`timescale 10ps / 10ps

`default_nettype none

module dds (
    input  wire logic [32-1:0] i_phase_inc,
    input  wire logic          i_phase_inc_valid,
    output      logic [36-1:0] o_cosine_data,
    output      logic [36-1:0] o_sine_data,
    input       logic          i_ready,
    input  wire logic          i_clock,
    input  wire logic          i_reset
);

// Phase increment
logic [32-1:0] phase_inc_reg;
logic [32-1:0] phase_accum;

always_ff @ (posedge i_clock) begin
    // Read input phase increment
    if (i_phase_inc_valid == 1'b1) begin
        phase_inc_reg <= i_phase_inc;
    end
    // Increment phase whenever an output is requested
    if (i_reset == 1'b1) begin
        phase_accum <= '0;
    end else if (i_ready == 1'b1) begin
        phase_accum <= phase_accum + phase_inc_reg;
    end
end

// Sine/Cosine Look Up Table
localparam integer WIDTH = 36;
localparam integer RESIDUAL_WIDTH = WIDTH-14;

logic signed [WIDTH-1:0]      cosine_reg0 /* synthesis syn_ramstyle="block_ram" */;
logic signed [WIDTH-1:0]      sine_reg0 /* synthesis syn_ramstyle="block_ram" */;
// logic [16+RESIDUAL_WIDTH-1:0] residual_reg0;

// Pipeline Stage 0
always_ff @ (posedge i_clock) begin
    if (i_ready == 1'b1) begin
        // Perform table look up
        case(phase_accum[32-1:32-14])
        0: begin
            cosine_reg0 <= 36'sb11111111111111111111111111111111111;
            sine_reg0   <= 36'sb0;
        end
        1: begin
            cosine_reg0 <= 36'sb11111111111111111111111011000100000;
            sine_reg0   <= 36'sb110010010000111111011010;
        end
        2: begin
            cosine_reg0 <= 36'sb11111111111111111111101100010000101;
            sine_reg0   <= 36'sb1100100100001111110110011;
        end
        3: begin
            cosine_reg0 <= 36'sb11111111111111111111010011100101011;
            sine_reg0   <= 36'sb10010110110010111110000111;
        end
        4: begin
            cosine_reg0 <= 36'sb11111111111111111110110001000010101;
            sine_reg0   <= 36'sb11001001000011111101010110;
        end
        5: begin
            cosine_reg0 <= 36'sb11111111111111111110000100101000010;
            sine_reg0   <= 36'sb11111011010100111100011101;
        end
        6: begin
            cosine_reg0 <= 36'sb11111111111111111101001110010110001;
            sine_reg0   <= 36'sb100101101100101111011011010;
        end
        7: begin
            cosine_reg0 <= 36'sb11111111111111111100001110001100011;
            sine_reg0   <= 36'sb101011111110110111010001100;
        end
        8: begin
            cosine_reg0 <= 36'sb11111111111111111011000100001011000;
            sine_reg0   <= 36'sb110010010000111111000110000;
        end
        9: begin
            cosine_reg0 <= 36'sb11111111111111111001110000010001111;
            sine_reg0   <= 36'sb111000100011000110111000100;
        end
        10: begin
            cosine_reg0 <= 36'sb11111111111111111000010010100001001;
            sine_reg0   <= 36'sb111110110101001110101000111;
        end
        11: begin
            cosine_reg0 <= 36'sb11111111111111110110101010111000111;
            sine_reg0   <= 36'sb1000101000111010110010110111;
        end
        12: begin
            cosine_reg0 <= 36'sb11111111111111110100111001011000111;
            sine_reg0   <= 36'sb1001011011001011110000010001;
        end
        13: begin
            cosine_reg0 <= 36'sb11111111111111110010111110000001001;
            sine_reg0   <= 36'sb1010001101011100101101010101;
        end
        14: begin
            cosine_reg0 <= 36'sb11111111111111110000111000110001111;
            sine_reg0   <= 36'sb1010111111101101101001111111;
        end
        15: begin
            cosine_reg0 <= 36'sb11111111111111101110101001101010111;
            sine_reg0   <= 36'sb1011110001111110100110001101;
        end
        16: begin
            cosine_reg0 <= 36'sb11111111111111101100010000101100011;
            sine_reg0   <= 36'sb1100100100001111100001111111;
        end
        17: begin
            cosine_reg0 <= 36'sb11111111111111101001101101110110001;
            sine_reg0   <= 36'sb1101010110100000011101010010;
        end
        18: begin
            cosine_reg0 <= 36'sb11111111111111100111000001001000010;
            sine_reg0   <= 36'sb1110001000110001011000000100;
        end
        19: begin
            cosine_reg0 <= 36'sb11111111111111100100001010100010110;
            sine_reg0   <= 36'sb1110111011000010010010010011;
        end
        20: begin
            cosine_reg0 <= 36'sb11111111111111100001001010000101100;
            sine_reg0   <= 36'sb1111101101010011001011111101;
        end
        21: begin
            cosine_reg0 <= 36'sb11111111111111011101111111110000110;
            sine_reg0   <= 36'sb10000011111100100000101000000;
        end
        22: begin
            cosine_reg0 <= 36'sb11111111111111011010101011100100011;
            sine_reg0   <= 36'sb10001010001110100111101011011;
        end
        23: begin
            cosine_reg0 <= 36'sb11111111111111010111001101100000010;
            sine_reg0   <= 36'sb10010000100000101110101001011;
        end
        24: begin
            cosine_reg0 <= 36'sb11111111111111010011100101100100101;
            sine_reg0   <= 36'sb10010110110010110101100001110;
        end
        25: begin
            cosine_reg0 <= 36'sb11111111111111001111110011110001010;
            sine_reg0   <= 36'sb10011101000100111100010100011;
        end
        26: begin
            cosine_reg0 <= 36'sb11111111111111001011111000000110011;
            sine_reg0   <= 36'sb10100011010111000011000001000;
        end
        27: begin
            cosine_reg0 <= 36'sb11111111111111000111110010100011110;
            sine_reg0   <= 36'sb10101001101001001001100111010;
        end
        28: begin
            cosine_reg0 <= 36'sb11111111111111000011100011001001101;
            sine_reg0   <= 36'sb10101111111011010000000111000;
        end
        29: begin
            cosine_reg0 <= 36'sb11111111111110111111001001110111111;
            sine_reg0   <= 36'sb10110110001101010110011111111;
        end
        30: begin
            cosine_reg0 <= 36'sb11111111111110111010100110101110011;
            sine_reg0   <= 36'sb10111100011111011100110001111;
        end
        31: begin
            cosine_reg0 <= 36'sb11111111111110110101111001101101011;
            sine_reg0   <= 36'sb11000010110001100010111100100;
        end
        32: begin
            cosine_reg0 <= 36'sb11111111111110110001000010110100110;
            sine_reg0   <= 36'sb11001001000011101000111111101;
        end
        33: begin
            cosine_reg0 <= 36'sb11111111111110101100000010000100100;
            sine_reg0   <= 36'sb11001111010101101110111011000;
        end
        34: begin
            cosine_reg0 <= 36'sb11111111111110100110110111011100101;
            sine_reg0   <= 36'sb11010101100111110100101110011;
        end
        35: begin
            cosine_reg0 <= 36'sb11111111111110100001100010111101010;
            sine_reg0   <= 36'sb11011011111001111010011001100;
        end
        36: begin
            cosine_reg0 <= 36'sb11111111111110011100000100100110001;
            sine_reg0   <= 36'sb11100010001011111111111100010;
        end
        37: begin
            cosine_reg0 <= 36'sb11111111111110010110011100010111100;
            sine_reg0   <= 36'sb11101000011110000101010110010;
        end
        38: begin
            cosine_reg0 <= 36'sb11111111111110010000101010010001010;
            sine_reg0   <= 36'sb11101110110000001010100111010;
        end
        39: begin
            cosine_reg0 <= 36'sb11111111111110001010101110010011100;
            sine_reg0   <= 36'sb11110101000010001111101111000;
        end
        40: begin
            cosine_reg0 <= 36'sb11111111111110000100101000011110000;
            sine_reg0   <= 36'sb11111011010100010100101101011;
        end
        41: begin
            cosine_reg0 <= 36'sb11111111111101111110011000110001000;
            sine_reg0   <= 36'sb100000001100110011001100010000;
        end
        42: begin
            cosine_reg0 <= 36'sb11111111111101110111111111001100100;
            sine_reg0   <= 36'sb100000111111000011110001100110;
        end
        43: begin
            cosine_reg0 <= 36'sb11111111111101110001011011110000011;
            sine_reg0   <= 36'sb100001110001010100010101101010;
        end
        44: begin
            cosine_reg0 <= 36'sb11111111111101101010101110011100101;
            sine_reg0   <= 36'sb100010100011100100111000011011;
        end
        45: begin
            cosine_reg0 <= 36'sb11111111111101100011110111010001011;
            sine_reg0   <= 36'sb100011010101110101011001110111;
        end
        46: begin
            cosine_reg0 <= 36'sb11111111111101011100110110001110100;
            sine_reg0   <= 36'sb100100001000000101111001111100;
        end
        47: begin
            cosine_reg0 <= 36'sb11111111111101010101101011010100001;
            sine_reg0   <= 36'sb100100111010010110011000100111;
        end
        48: begin
            cosine_reg0 <= 36'sb11111111111101001110010110100010010;
            sine_reg0   <= 36'sb100101101100100110110101111000;
        end
        49: begin
            cosine_reg0 <= 36'sb11111111111101000110110111111000110;
            sine_reg0   <= 36'sb100110011110110111010001101011;
        end
        50: begin
            cosine_reg0 <= 36'sb11111111111100111111001111010111110;
            sine_reg0   <= 36'sb100111010001000111101100000000;
        end
        51: begin
            cosine_reg0 <= 36'sb11111111111100110111011100111111001;
            sine_reg0   <= 36'sb101000000011011000000100110011;
        end
        52: begin
            cosine_reg0 <= 36'sb11111111111100101111100000101111000;
            sine_reg0   <= 36'sb101000110101101000011100000100;
        end
        53: begin
            cosine_reg0 <= 36'sb11111111111100100111011010100111011;
            sine_reg0   <= 36'sb101001100111111000110001110000;
        end
        54: begin
            cosine_reg0 <= 36'sb11111111111100011111001010101000010;
            sine_reg0   <= 36'sb101010011010001001000101110101;
        end
        55: begin
            cosine_reg0 <= 36'sb11111111111100010110110000110001101;
            sine_reg0   <= 36'sb101011001100011001011000010010;
        end
        56: begin
            cosine_reg0 <= 36'sb11111111111100001110001101000011011;
            sine_reg0   <= 36'sb101011111110101001101001000100;
        end
        57: begin
            cosine_reg0 <= 36'sb11111111111100000101011111011101110;
            sine_reg0   <= 36'sb101100110000111001111000001001;
        end
        58: begin
            cosine_reg0 <= 36'sb11111111111011111100101000000000100;
            sine_reg0   <= 36'sb101101100011001010000101100001;
        end
        59: begin
            cosine_reg0 <= 36'sb11111111111011110011100110101011110;
            sine_reg0   <= 36'sb101110010101011010010001000111;
        end
        60: begin
            cosine_reg0 <= 36'sb11111111111011101010011011011111101;
            sine_reg0   <= 36'sb101111000111101010011010111100;
        end
        61: begin
            cosine_reg0 <= 36'sb11111111111011100001000110011011111;
            sine_reg0   <= 36'sb101111111001111010100010111100;
        end
        62: begin
            cosine_reg0 <= 36'sb11111111111011010111100111100000110;
            sine_reg0   <= 36'sb110000101100001010101001000110;
        end
        63: begin
            cosine_reg0 <= 36'sb11111111111011001101111110101110001;
            sine_reg0   <= 36'sb110001011110011010101101011000;
        end
        64: begin
            cosine_reg0 <= 36'sb11111111111011000100001100000100000;
            sine_reg0   <= 36'sb110010010000101010101111101111;
        end
        65: begin
            cosine_reg0 <= 36'sb11111111111010111010001111100010100;
            sine_reg0   <= 36'sb110011000010111010110000001011;
        end
        66: begin
            cosine_reg0 <= 36'sb11111111111010110000001001001001011;
            sine_reg0   <= 36'sb110011110101001010101110101001;
        end
        67: begin
            cosine_reg0 <= 36'sb11111111111010100101111000111001000;
            sine_reg0   <= 36'sb110100100111011010101011000111;
        end
        68: begin
            cosine_reg0 <= 36'sb11111111111010011011011110110001000;
            sine_reg0   <= 36'sb110101011001101010100101100011;
        end
        69: begin
            cosine_reg0 <= 36'sb11111111111010010000111010110001101;
            sine_reg0   <= 36'sb110110001011111010011101111011;
        end
        70: begin
            cosine_reg0 <= 36'sb11111111111010000110001100111010111;
            sine_reg0   <= 36'sb110110111110001010010100001101;
        end
        71: begin
            cosine_reg0 <= 36'sb11111111111001111011010101001100101;
            sine_reg0   <= 36'sb110111110000011010001000011000;
        end
        72: begin
            cosine_reg0 <= 36'sb11111111111001110000010011100111000;
            sine_reg0   <= 36'sb111000100010101001111010011010;
        end
        73: begin
            cosine_reg0 <= 36'sb11111111111001100101001000001001111;
            sine_reg0   <= 36'sb111001010100111001101010010000;
        end
        74: begin
            cosine_reg0 <= 36'sb11111111111001011001110010110101011;
            sine_reg0   <= 36'sb111010000111001001010111111000;
        end
        75: begin
            cosine_reg0 <= 36'sb11111111111001001110010011101001100;
            sine_reg0   <= 36'sb111010111001011001000011010001;
        end
        76: begin
            cosine_reg0 <= 36'sb11111111111001000010101010100110010;
            sine_reg0   <= 36'sb111011101011101000101100011001;
        end
        77: begin
            cosine_reg0 <= 36'sb11111111111000110110110111101011101;
            sine_reg0   <= 36'sb111100011101111000010011001101;
        end
        78: begin
            cosine_reg0 <= 36'sb11111111111000101010111010111001101;
            sine_reg0   <= 36'sb111101010000000111110111101100;
        end
        79: begin
            cosine_reg0 <= 36'sb11111111111000011110110100010000010;
            sine_reg0   <= 36'sb111110000010010111011001110101;
        end
        80: begin
            cosine_reg0 <= 36'sb11111111111000010010100011101111011;
            sine_reg0   <= 36'sb111110110100100110111001100100;
        end
        81: begin
            cosine_reg0 <= 36'sb11111111111000000110001001010111010;
            sine_reg0   <= 36'sb111111100110110110010110111000;
        end
        82: begin
            cosine_reg0 <= 36'sb11111111110111111001100101000111111;
            sine_reg0   <= 36'sb1000000011001000101110001101111;
        end
        83: begin
            cosine_reg0 <= 36'sb11111111110111101100110111000001000;
            sine_reg0   <= 36'sb1000001001011010101001010000111;
        end
        84: begin
            cosine_reg0 <= 36'sb11111111110111011111111111000010111;
            sine_reg0   <= 36'sb1000001111101100100011111111110;
        end
        85: begin
            cosine_reg0 <= 36'sb11111111110111010010111101001101011;
            sine_reg0   <= 36'sb1000010101111110011110011010011;
        end
        86: begin
            cosine_reg0 <= 36'sb11111111110111000101110001100000101;
            sine_reg0   <= 36'sb1000011100010000011000100000011;
        end
        87: begin
            cosine_reg0 <= 36'sb11111111110110111000011011111100100;
            sine_reg0   <= 36'sb1000100010100010010010010001100;
        end
        88: begin
            cosine_reg0 <= 36'sb11111111110110101010111100100001000;
            sine_reg0   <= 36'sb1000101000110100001011101101101;
        end
        89: begin
            cosine_reg0 <= 36'sb11111111110110011101010011001110011;
            sine_reg0   <= 36'sb1000101111000110000100110100011;
        end
        90: begin
            cosine_reg0 <= 36'sb11111111110110001111100000000100011;
            sine_reg0   <= 36'sb1000110101010111111101100101101;
        end
        91: begin
            cosine_reg0 <= 36'sb11111111110110000001100011000011001;
            sine_reg0   <= 36'sb1000111011101001110110000001001;
        end
        92: begin
            cosine_reg0 <= 36'sb11111111110101110011011100001010100;
            sine_reg0   <= 36'sb1001000001111011101110000110100;
        end
        93: begin
            cosine_reg0 <= 36'sb11111111110101100101001011011010110;
            sine_reg0   <= 36'sb1001001000001101100101110101101;
        end
        94: begin
            cosine_reg0 <= 36'sb11111111110101010110110000110011101;
            sine_reg0   <= 36'sb1001001110011111011101001110001;
        end
        95: begin
            cosine_reg0 <= 36'sb11111111110101001000001100010101011;
            sine_reg0   <= 36'sb1001010100110001010100010000000;
        end
        96: begin
            cosine_reg0 <= 36'sb11111111110100111001011101111111111;
            sine_reg0   <= 36'sb1001011011000011001010111010110;
        end
        97: begin
            cosine_reg0 <= 36'sb11111111110100101010100101110011001;
            sine_reg0   <= 36'sb1001100001010101000001001110011;
        end
        98: begin
            cosine_reg0 <= 36'sb11111111110100011011100011101111001;
            sine_reg0   <= 36'sb1001100111100110110111001010011;
        end
        99: begin
            cosine_reg0 <= 36'sb11111111110100001100010111110011111;
            sine_reg0   <= 36'sb1001101101111000101100101110110;
        end
        100: begin
            cosine_reg0 <= 36'sb11111111110011111101000010000001100;
            sine_reg0   <= 36'sb1001110100001010100001111011001;
        end
        101: begin
            cosine_reg0 <= 36'sb11111111110011101101100010010111111;
            sine_reg0   <= 36'sb1001111010011100010110101111010;
        end
        102: begin
            cosine_reg0 <= 36'sb11111111110011011101111000110111001;
            sine_reg0   <= 36'sb1010000000101110001011001011000;
        end
        103: begin
            cosine_reg0 <= 36'sb11111111110011001110000101011111010;
            sine_reg0   <= 36'sb1010000110111111111111001110000;
        end
        104: begin
            cosine_reg0 <= 36'sb11111111110010111110001000010000001;
            sine_reg0   <= 36'sb1010001101010001110010111000000;
        end
        105: begin
            cosine_reg0 <= 36'sb11111111110010101110000001001001111;
            sine_reg0   <= 36'sb1010010011100011100110001000111;
        end
        106: begin
            cosine_reg0 <= 36'sb11111111110010011101110000001100100;
            sine_reg0   <= 36'sb1010011001110101011001000000010;
        end
        107: begin
            cosine_reg0 <= 36'sb11111111110010001101010101011000000;
            sine_reg0   <= 36'sb1010100000000111001011011110000;
        end
        108: begin
            cosine_reg0 <= 36'sb11111111110001111100110000101100011;
            sine_reg0   <= 36'sb1010100110011000111101100001111;
        end
        109: begin
            cosine_reg0 <= 36'sb11111111110001101100000010001001101;
            sine_reg0   <= 36'sb1010101100101010101111001011100;
        end
        110: begin
            cosine_reg0 <= 36'sb11111111110001011011001001101111110;
            sine_reg0   <= 36'sb1010110010111100100000011010111;
        end
        111: begin
            cosine_reg0 <= 36'sb11111111110001001010000111011110110;
            sine_reg0   <= 36'sb1010111001001110010001001111100;
        end
        112: begin
            cosine_reg0 <= 36'sb11111111110000111000111011010110110;
            sine_reg0   <= 36'sb1010111111100000000001101001010;
        end
        113: begin
            cosine_reg0 <= 36'sb11111111110000100111100101010111101;
            sine_reg0   <= 36'sb1011000101110001110001100111111;
        end
        114: begin
            cosine_reg0 <= 36'sb11111111110000010110000101100001100;
            sine_reg0   <= 36'sb1011001100000011100001001011010;
        end
        115: begin
            cosine_reg0 <= 36'sb11111111110000000100011011110100010;
            sine_reg0   <= 36'sb1011010010010101010000010010111;
        end
        116: begin
            cosine_reg0 <= 36'sb11111111101111110010101000010000000;
            sine_reg0   <= 36'sb1011011000100110111110111110110;
        end
        117: begin
            cosine_reg0 <= 36'sb11111111101111100000101010110100101;
            sine_reg0   <= 36'sb1011011110111000101101001110100;
        end
        118: begin
            cosine_reg0 <= 36'sb11111111101111001110100011100010011;
            sine_reg0   <= 36'sb1011100101001010011011000001111;
        end
        119: begin
            cosine_reg0 <= 36'sb11111111101110111100010010011001000;
            sine_reg0   <= 36'sb1011101011011100001000011000110;
        end
        120: begin
            cosine_reg0 <= 36'sb11111111101110101001110111011000110;
            sine_reg0   <= 36'sb1011110001101101110101010010110;
        end
        121: begin
            cosine_reg0 <= 36'sb11111111101110010111010010100001011;
            sine_reg0   <= 36'sb1011110111111111100001101111110;
        end
        122: begin
            cosine_reg0 <= 36'sb11111111101110000100100011110011001;
            sine_reg0   <= 36'sb1011111110010001001101101111011;
        end
        123: begin
            cosine_reg0 <= 36'sb11111111101101110001101011001101111;
            sine_reg0   <= 36'sb1100000100100010111001010001100;
        end
        124: begin
            cosine_reg0 <= 36'sb11111111101101011110101000110001110;
            sine_reg0   <= 36'sb1100001010110100100100010101111;
        end
        125: begin
            cosine_reg0 <= 36'sb11111111101101001011011100011110101;
            sine_reg0   <= 36'sb1100010001000110001110111100001;
        end
        126: begin
            cosine_reg0 <= 36'sb11111111101100111000000110010100100;
            sine_reg0   <= 36'sb1100010111010111111001000100010;
        end
        127: begin
            cosine_reg0 <= 36'sb11111111101100100100100110010011100;
            sine_reg0   <= 36'sb1100011101101001100010101101110;
        end
        128: begin
            cosine_reg0 <= 36'sb11111111101100010000111100011011101;
            sine_reg0   <= 36'sb1100100011111011001011111000100;
        end
        129: begin
            cosine_reg0 <= 36'sb11111111101011111101001000101100111;
            sine_reg0   <= 36'sb1100101010001100110100100100010;
        end
        130: begin
            cosine_reg0 <= 36'sb11111111101011101001001011000111010;
            sine_reg0   <= 36'sb1100110000011110011100110000111;
        end
        131: begin
            cosine_reg0 <= 36'sb11111111101011010101000011101010110;
            sine_reg0   <= 36'sb1100110110110000000100011101111;
        end
        132: begin
            cosine_reg0 <= 36'sb11111111101011000000110010010111011;
            sine_reg0   <= 36'sb1100111101000001101011101011010;
        end
        133: begin
            cosine_reg0 <= 36'sb11111111101010101100010111001101001;
            sine_reg0   <= 36'sb1101000011010011010010011000101;
        end
        134: begin
            cosine_reg0 <= 36'sb11111111101010010111110010001100000;
            sine_reg0   <= 36'sb1101001001100100111000100101111;
        end
        135: begin
            cosine_reg0 <= 36'sb11111111101010000011000011010100001;
            sine_reg0   <= 36'sb1101001111110110011110010010101;
        end
        136: begin
            cosine_reg0 <= 36'sb11111111101001101110001010100101011;
            sine_reg0   <= 36'sb1101010110001000000011011110101;
        end
        137: begin
            cosine_reg0 <= 36'sb11111111101001011001001000000000000;
            sine_reg0   <= 36'sb1101011100011001101000001001110;
        end
        138: begin
            cosine_reg0 <= 36'sb11111111101001000011111011100011101;
            sine_reg0   <= 36'sb1101100010101011001100010011110;
        end
        139: begin
            cosine_reg0 <= 36'sb11111111101000101110100101010000101;
            sine_reg0   <= 36'sb1101101000111100101111111100010;
        end
        140: begin
            cosine_reg0 <= 36'sb11111111101000011001000101000110111;
            sine_reg0   <= 36'sb1101101111001110010011000011010;
        end
        141: begin
            cosine_reg0 <= 36'sb11111111101000000011011011000110010;
            sine_reg0   <= 36'sb1101110101011111110101101000010;
        end
        142: begin
            cosine_reg0 <= 36'sb11111111100111101101100111001111000;
            sine_reg0   <= 36'sb1101111011110001010111101011000;
        end
        143: begin
            cosine_reg0 <= 36'sb11111111100111010111101001100001000;
            sine_reg0   <= 36'sb1110000010000010111001001011100;
        end
        144: begin
            cosine_reg0 <= 36'sb11111111100111000001100001111100010;
            sine_reg0   <= 36'sb1110001000010100011010001001011;
        end
        145: begin
            cosine_reg0 <= 36'sb11111111100110101011010000100000111;
            sine_reg0   <= 36'sb1110001110100101111010100100011;
        end
        146: begin
            cosine_reg0 <= 36'sb11111111100110010100110101001110111;
            sine_reg0   <= 36'sb1110010100110111011010011100010;
        end
        147: begin
            cosine_reg0 <= 36'sb11111111100101111110010000000110001;
            sine_reg0   <= 36'sb1110011011001000111001110000110;
        end
        148: begin
            cosine_reg0 <= 36'sb11111111100101100111100001000110110;
            sine_reg0   <= 36'sb1110100001011010011000100001110;
        end
        149: begin
            cosine_reg0 <= 36'sb11111111100101010000101000010000101;
            sine_reg0   <= 36'sb1110100111101011110110101110111;
        end
        150: begin
            cosine_reg0 <= 36'sb11111111100100111001100101100100000;
            sine_reg0   <= 36'sb1110101101111101010100010111111;
        end
        151: begin
            cosine_reg0 <= 36'sb11111111100100100010011001000000110;
            sine_reg0   <= 36'sb1110110100001110110001011100101;
        end
        152: begin
            cosine_reg0 <= 36'sb11111111100100001011000010100110111;
            sine_reg0   <= 36'sb1110111010100000001101111100110;
        end
        153: begin
            cosine_reg0 <= 36'sb11111111100011110011100010010110100;
            sine_reg0   <= 36'sb1111000000110001101001111000001;
        end
        154: begin
            cosine_reg0 <= 36'sb11111111100011011011111000001111100;
            sine_reg0   <= 36'sb1111000111000011000101001110011;
        end
        155: begin
            cosine_reg0 <= 36'sb11111111100011000100000100010001111;
            sine_reg0   <= 36'sb1111001101010100011111111111100;
        end
        156: begin
            cosine_reg0 <= 36'sb11111111100010101100000110011101111;
            sine_reg0   <= 36'sb1111010011100101111010001011000;
        end
        157: begin
            cosine_reg0 <= 36'sb11111111100010010011111110110011010;
            sine_reg0   <= 36'sb1111011001110111010011110000110;
        end
        158: begin
            cosine_reg0 <= 36'sb11111111100001111011101101010010000;
            sine_reg0   <= 36'sb1111100000001000101100110000100;
        end
        159: begin
            cosine_reg0 <= 36'sb11111111100001100011010001111010011;
            sine_reg0   <= 36'sb1111100110011010000101001010000;
        end
        160: begin
            cosine_reg0 <= 36'sb11111111100001001010101100101100011;
            sine_reg0   <= 36'sb1111101100101011011100111101000;
        end
        161: begin
            cosine_reg0 <= 36'sb11111111100000110001111101100111110;
            sine_reg0   <= 36'sb1111110010111100110100001001010;
        end
        162: begin
            cosine_reg0 <= 36'sb11111111100000011001000100101100110;
            sine_reg0   <= 36'sb1111111001001110001010101110100;
        end
        163: begin
            cosine_reg0 <= 36'sb11111111100000000000000001111011010;
            sine_reg0   <= 36'sb1111111111011111100000101100101;
        end
        164: begin
            cosine_reg0 <= 36'sb11111111011111100110110101010011011;
            sine_reg0   <= 36'sb10000000101110000110110000011010;
        end
        165: begin
            cosine_reg0 <= 36'sb11111111011111001101011110110101001;
            sine_reg0   <= 36'sb10000001100000010001010110010001;
        end
        166: begin
            cosine_reg0 <= 36'sb11111111011110110011111110100000011;
            sine_reg0   <= 36'sb10000010010010011011110111001001;
        end
        167: begin
            cosine_reg0 <= 36'sb11111111011110011010010100010101011;
            sine_reg0   <= 36'sb10000011000100100110010010111111;
        end
        168: begin
            cosine_reg0 <= 36'sb11111111011110000000100000010100000;
            sine_reg0   <= 36'sb10000011110110110000101001110010;
        end
        169: begin
            cosine_reg0 <= 36'sb11111111011101100110100010011100010;
            sine_reg0   <= 36'sb10000100101000111010111011100000;
        end
        170: begin
            cosine_reg0 <= 36'sb11111111011101001100011010101110001;
            sine_reg0   <= 36'sb10000101011011000101001000000110;
        end
        171: begin
            cosine_reg0 <= 36'sb11111111011100110010001001001001110;
            sine_reg0   <= 36'sb10000110001101001111001111100011;
        end
        172: begin
            cosine_reg0 <= 36'sb11111111011100010111101101101111000;
            sine_reg0   <= 36'sb10000110111111011001010001110101;
        end
        173: begin
            cosine_reg0 <= 36'sb11111111011011111101001000011110000;
            sine_reg0   <= 36'sb10000111110001100011001110111010;
        end
        174: begin
            cosine_reg0 <= 36'sb11111111011011100010011001010110110;
            sine_reg0   <= 36'sb10001000100011101101000110110000;
        end
        175: begin
            cosine_reg0 <= 36'sb11111111011011000111100000011001010;
            sine_reg0   <= 36'sb10001001010101110110111001010101;
        end
        176: begin
            cosine_reg0 <= 36'sb11111111011010101100011101100101101;
            sine_reg0   <= 36'sb10001010001000000000100110100111;
        end
        177: begin
            cosine_reg0 <= 36'sb11111111011010010001010000111011101;
            sine_reg0   <= 36'sb10001010111010001010001110100100;
        end
        178: begin
            cosine_reg0 <= 36'sb11111111011001110101111010011011100;
            sine_reg0   <= 36'sb10001011101100010011110001001010;
        end
        179: begin
            cosine_reg0 <= 36'sb11111111011001011010011010000101001;
            sine_reg0   <= 36'sb10001100011110011101001110011000;
        end
        180: begin
            cosine_reg0 <= 36'sb11111111011000111110101111111000101;
            sine_reg0   <= 36'sb10001101010000100110100110001011;
        end
        181: begin
            cosine_reg0 <= 36'sb11111111011000100010111011110110000;
            sine_reg0   <= 36'sb10001110000010101111111000100010;
        end
        182: begin
            cosine_reg0 <= 36'sb11111111011000000110111101111101010;
            sine_reg0   <= 36'sb10001110110100111001000101011010;
        end
        183: begin
            cosine_reg0 <= 36'sb11111111010111101010110110001110011;
            sine_reg0   <= 36'sb10001111100111000010001100110010;
        end
        184: begin
            cosine_reg0 <= 36'sb11111111010111001110100100101001011;
            sine_reg0   <= 36'sb10010000011001001011001110100111;
        end
        185: begin
            cosine_reg0 <= 36'sb11111111010110110010001001001110010;
            sine_reg0   <= 36'sb10010001001011010100001010111000;
        end
        186: begin
            cosine_reg0 <= 36'sb11111111010110010101100011111101001;
            sine_reg0   <= 36'sb10010001111101011101000001100011;
        end
        187: begin
            cosine_reg0 <= 36'sb11111111010101111000110100110110000;
            sine_reg0   <= 36'sb10010010101111100101110010100110;
        end
        188: begin
            cosine_reg0 <= 36'sb11111111010101011011111011111000110;
            sine_reg0   <= 36'sb10010011100001101110011101111111;
        end
        189: begin
            cosine_reg0 <= 36'sb11111111010100111110111001000101100;
            sine_reg0   <= 36'sb10010100010011110111000011101100;
        end
        190: begin
            cosine_reg0 <= 36'sb11111111010100100001101100011100010;
            sine_reg0   <= 36'sb10010101000101111111100011101010;
        end
        191: begin
            cosine_reg0 <= 36'sb11111111010100000100010101111101001;
            sine_reg0   <= 36'sb10010101111000000111111101111001;
        end
        192: begin
            cosine_reg0 <= 36'sb11111111010011100110110101100111111;
            sine_reg0   <= 36'sb10010110101010010000010010010110;
        end
        193: begin
            cosine_reg0 <= 36'sb11111111010011001001001011011100110;
            sine_reg0   <= 36'sb10010111011100011000100001000000;
        end
        194: begin
            cosine_reg0 <= 36'sb11111111010010101011010111011011110;
            sine_reg0   <= 36'sb10011000001110100000101001110011;
        end
        195: begin
            cosine_reg0 <= 36'sb11111111010010001101011001100100111;
            sine_reg0   <= 36'sb10011001000000101000101100101111;
        end
        196: begin
            cosine_reg0 <= 36'sb11111111010001101111010001111000000;
            sine_reg0   <= 36'sb10011001110010110000101001110010;
        end
        197: begin
            cosine_reg0 <= 36'sb11111111010001010001000000010101010;
            sine_reg0   <= 36'sb10011010100100111000100000111001;
        end
        198: begin
            cosine_reg0 <= 36'sb11111111010000110010100100111100110;
            sine_reg0   <= 36'sb10011011010111000000010010000011;
        end
        199: begin
            cosine_reg0 <= 36'sb11111111010000010011111111101110011;
            sine_reg0   <= 36'sb10011100001001000111111101001101;
        end
        200: begin
            cosine_reg0 <= 36'sb11111111001111110101010000101010001;
            sine_reg0   <= 36'sb10011100111011001111100010010110;
        end
        201: begin
            cosine_reg0 <= 36'sb11111111001111010110010111110000001;
            sine_reg0   <= 36'sb10011101101101010111000001011100;
        end
        202: begin
            cosine_reg0 <= 36'sb11111111001110110111010101000000011;
            sine_reg0   <= 36'sb10011110011111011110011010011101;
        end
        203: begin
            cosine_reg0 <= 36'sb11111111001110011000001000011010110;
            sine_reg0   <= 36'sb10011111010001100101101101010110;
        end
        204: begin
            cosine_reg0 <= 36'sb11111111001101111000110001111111100;
            sine_reg0   <= 36'sb10100000000011101100111010000111;
        end
        205: begin
            cosine_reg0 <= 36'sb11111111001101011001010001101110100;
            sine_reg0   <= 36'sb10100000110101110100000000101101;
        end
        206: begin
            cosine_reg0 <= 36'sb11111111001100111001100111100111110;
            sine_reg0   <= 36'sb10100001100111111011000001000110;
        end
        207: begin
            cosine_reg0 <= 36'sb11111111001100011001110011101011011;
            sine_reg0   <= 36'sb10100010011010000001111011010000;
        end
        208: begin
            cosine_reg0 <= 36'sb11111111001011111001110101111001011;
            sine_reg0   <= 36'sb10100011001100001000101111001001;
        end
        209: begin
            cosine_reg0 <= 36'sb11111111001011011001101110010001101;
            sine_reg0   <= 36'sb10100011111110001111011100110000;
        end
        210: begin
            cosine_reg0 <= 36'sb11111111001010111001011100110100010;
            sine_reg0   <= 36'sb10100100110000010110000100000010;
        end
        211: begin
            cosine_reg0 <= 36'sb11111111001010011001000001100001011;
            sine_reg0   <= 36'sb10100101100010011100100100111110;
        end
        212: begin
            cosine_reg0 <= 36'sb11111111001001111000011100011000110;
            sine_reg0   <= 36'sb10100110010100100010111111100001;
        end
        213: begin
            cosine_reg0 <= 36'sb11111111001001010111101101011010110;
            sine_reg0   <= 36'sb10100111000110101001010011101010;
        end
        214: begin
            cosine_reg0 <= 36'sb11111111001000110110110100100111000;
            sine_reg0   <= 36'sb10100111111000101111100001010110;
        end
        215: begin
            cosine_reg0 <= 36'sb11111111001000010101110001111101111;
            sine_reg0   <= 36'sb10101000101010110101101000100100;
        end
        216: begin
            cosine_reg0 <= 36'sb11111111000111110100100101011111001;
            sine_reg0   <= 36'sb10101001011100111011101001010010;
        end
        217: begin
            cosine_reg0 <= 36'sb11111111000111010011001111001011000;
            sine_reg0   <= 36'sb10101010001111000001100011011110;
        end
        218: begin
            cosine_reg0 <= 36'sb11111111000110110001101111000001011;
            sine_reg0   <= 36'sb10101011000001000111010111000110;
        end
        219: begin
            cosine_reg0 <= 36'sb11111111000110010000000101000010010;
            sine_reg0   <= 36'sb10101011110011001101000100001000;
        end
        220: begin
            cosine_reg0 <= 36'sb11111111000101101110010001001101110;
            sine_reg0   <= 36'sb10101100100101010010101010100010;
        end
        221: begin
            cosine_reg0 <= 36'sb11111111000101001100010011100011111;
            sine_reg0   <= 36'sb10101101010111011000001010010010;
        end
        222: begin
            cosine_reg0 <= 36'sb11111111000100101010001100000100100;
            sine_reg0   <= 36'sb10101110001001011101100011010111;
        end
        223: begin
            cosine_reg0 <= 36'sb11111111000100000111111010101111111;
            sine_reg0   <= 36'sb10101110111011100010110101101110;
        end
        224: begin
            cosine_reg0 <= 36'sb11111111000011100101011111100101110;
            sine_reg0   <= 36'sb10101111101101101000000001010101;
        end
        225: begin
            cosine_reg0 <= 36'sb11111111000011000010111010100110100;
            sine_reg0   <= 36'sb10110000011111101101000110001010;
        end
        226: begin
            cosine_reg0 <= 36'sb11111111000010100000001011110001110;
            sine_reg0   <= 36'sb10110001010001110010000100001100;
        end
        227: begin
            cosine_reg0 <= 36'sb11111111000001111101010011000111111;
            sine_reg0   <= 36'sb10110010000011110110111011011001;
        end
        228: begin
            cosine_reg0 <= 36'sb11111111000001011010010000101000101;
            sine_reg0   <= 36'sb10110010110101111011101011101110;
        end
        229: begin
            cosine_reg0 <= 36'sb11111111000000110111000100010100001;
            sine_reg0   <= 36'sb10110011101000000000010101001011;
        end
        230: begin
            cosine_reg0 <= 36'sb11111111000000010011101110001010100;
            sine_reg0   <= 36'sb10110100011010000100110111101011;
        end
        231: begin
            cosine_reg0 <= 36'sb11111110111111110000001110001011101;
            sine_reg0   <= 36'sb10110101001100001001010011001111;
        end
        232: begin
            cosine_reg0 <= 36'sb11111110111111001100100100010111101;
            sine_reg0   <= 36'sb10110101111110001101100111110100;
        end
        233: begin
            cosine_reg0 <= 36'sb11111110111110101000110000101110011;
            sine_reg0   <= 36'sb10110110110000010001110101010111;
        end
        234: begin
            cosine_reg0 <= 36'sb11111110111110000100110011010000001;
            sine_reg0   <= 36'sb10110111100010010101111011111000;
        end
        235: begin
            cosine_reg0 <= 36'sb11111110111101100000101011111100101;
            sine_reg0   <= 36'sb10111000010100011001111011010100;
        end
        236: begin
            cosine_reg0 <= 36'sb11111110111100111100011010110100001;
            sine_reg0   <= 36'sb10111001000110011101110011101001;
        end
        237: begin
            cosine_reg0 <= 36'sb11111110111100010111111111110110100;
            sine_reg0   <= 36'sb10111001111000100001100100110101;
        end
        238: begin
            cosine_reg0 <= 36'sb11111110111011110011011011000011110;
            sine_reg0   <= 36'sb10111010101010100101001110110111;
        end
        239: begin
            cosine_reg0 <= 36'sb11111110111011001110101100011100001;
            sine_reg0   <= 36'sb10111011011100101000110001101100;
        end
        240: begin
            cosine_reg0 <= 36'sb11111110111010101001110011111111011;
            sine_reg0   <= 36'sb10111100001110101100001101010011;
        end
        241: begin
            cosine_reg0 <= 36'sb11111110111010000100110001101101110;
            sine_reg0   <= 36'sb10111101000000101111100001101001;
        end
        242: begin
            cosine_reg0 <= 36'sb11111110111001011111100101100111001;
            sine_reg0   <= 36'sb10111101110010110010101110101101;
        end
        243: begin
            cosine_reg0 <= 36'sb11111110111000111010001111101011101;
            sine_reg0   <= 36'sb10111110100100110101110100011100;
        end
        244: begin
            cosine_reg0 <= 36'sb11111110111000010100101111111011001;
            sine_reg0   <= 36'sb10111111010110111000110010110110;
        end
        245: begin
            cosine_reg0 <= 36'sb11111110110111101111000110010101110;
            sine_reg0   <= 36'sb11000000001000111011101001110111;
        end
        246: begin
            cosine_reg0 <= 36'sb11111110110111001001010010111011100;
            sine_reg0   <= 36'sb11000000111010111110011001011110;
        end
        247: begin
            cosine_reg0 <= 36'sb11111110110110100011010101101100011;
            sine_reg0   <= 36'sb11000001101101000001000001101001;
        end
        248: begin
            cosine_reg0 <= 36'sb11111110110101111101001110101000100;
            sine_reg0   <= 36'sb11000010011111000011100010010110;
        end
        249: begin
            cosine_reg0 <= 36'sb11111110110101010110111101101111110;
            sine_reg0   <= 36'sb11000011010001000101111011100011;
        end
        250: begin
            cosine_reg0 <= 36'sb11111110110100110000100011000010011;
            sine_reg0   <= 36'sb11000100000011001000001101001111;
        end
        251: begin
            cosine_reg0 <= 36'sb11111110110100001001111110100000001;
            sine_reg0   <= 36'sb11000100110101001010010111010110;
        end
        252: begin
            cosine_reg0 <= 36'sb11111110110011100011010000001001001;
            sine_reg0   <= 36'sb11000101100111001100011001111000;
        end
        253: begin
            cosine_reg0 <= 36'sb11111110110010111100010111111101100;
            sine_reg0   <= 36'sb11000110011001001110010100110011;
        end
        254: begin
            cosine_reg0 <= 36'sb11111110110010010101010101111101001;
            sine_reg0   <= 36'sb11000111001011010000001000000100;
        end
        255: begin
            cosine_reg0 <= 36'sb11111110110001101110001010001000001;
            sine_reg0   <= 36'sb11000111111101010001110011101001;
        end
        256: begin
            cosine_reg0 <= 36'sb11111110110001000110110100011110011;
            sine_reg0   <= 36'sb11001000101111010011010111100001;
        end
        257: begin
            cosine_reg0 <= 36'sb11111110110000011111010101000000001;
            sine_reg0   <= 36'sb11001001100001010100110011101010;
        end
        258: begin
            cosine_reg0 <= 36'sb11111110101111110111101011101101010;
            sine_reg0   <= 36'sb11001010010011010110001000000010;
        end
        259: begin
            cosine_reg0 <= 36'sb11111110101111001111111000100101111;
            sine_reg0   <= 36'sb11001011000101010111010100100110;
        end
        260: begin
            cosine_reg0 <= 36'sb11111110101110100111111011101001111;
            sine_reg0   <= 36'sb11001011110111011000011001010101;
        end
        261: begin
            cosine_reg0 <= 36'sb11111110101101111111110100111001011;
            sine_reg0   <= 36'sb11001100101001011001010110001110;
        end
        262: begin
            cosine_reg0 <= 36'sb11111110101101010111100100010100100;
            sine_reg0   <= 36'sb11001101011011011010001011001101;
        end
        263: begin
            cosine_reg0 <= 36'sb11111110101100101111001001111011000;
            sine_reg0   <= 36'sb11001110001101011010111000010001;
        end
        264: begin
            cosine_reg0 <= 36'sb11111110101100000110100101101101001;
            sine_reg0   <= 36'sb11001110111111011011011101011001;
        end
        265: begin
            cosine_reg0 <= 36'sb11111110101011011101110111101010110;
            sine_reg0   <= 36'sb11001111110001011011111010100010;
        end
        266: begin
            cosine_reg0 <= 36'sb11111110101010110100111111110100001;
            sine_reg0   <= 36'sb11010000100011011100001111101010;
        end
        267: begin
            cosine_reg0 <= 36'sb11111110101010001011111110001001000;
            sine_reg0   <= 36'sb11010001010101011100011100110000;
        end
        268: begin
            cosine_reg0 <= 36'sb11111110101001100010110010101001101;
            sine_reg0   <= 36'sb11010010000111011100100001110001;
        end
        269: begin
            cosine_reg0 <= 36'sb11111110101000111001011101010101111;
            sine_reg0   <= 36'sb11010010111001011100011110101100;
        end
        270: begin
            cosine_reg0 <= 36'sb11111110101000001111111110001101110;
            sine_reg0   <= 36'sb11010011101011011100010011011110;
        end
        271: begin
            cosine_reg0 <= 36'sb11111110100111100110010101010001100;
            sine_reg0   <= 36'sb11010100011101011100000000000110;
        end
        272: begin
            cosine_reg0 <= 36'sb11111110100110111100100010100001000;
            sine_reg0   <= 36'sb11010101001111011011100100100010;
        end
        273: begin
            cosine_reg0 <= 36'sb11111110100110010010100101111100001;
            sine_reg0   <= 36'sb11010110000001011011000000110000;
        end
        274: begin
            cosine_reg0 <= 36'sb11111110100101101000011111100011001;
            sine_reg0   <= 36'sb11010110110011011010010100101110;
        end
        275: begin
            cosine_reg0 <= 36'sb11111110100100111110001111010110000;
            sine_reg0   <= 36'sb11010111100101011001100000011001;
        end
        276: begin
            cosine_reg0 <= 36'sb11111110100100010011110101010100110;
            sine_reg0   <= 36'sb11011000010111011000100011110001;
        end
        277: begin
            cosine_reg0 <= 36'sb11111110100011101001010001011111011;
            sine_reg0   <= 36'sb11011001001001010111011110110011;
        end
        278: begin
            cosine_reg0 <= 36'sb11111110100010111110100011110101111;
            sine_reg0   <= 36'sb11011001111011010110010001011101;
        end
        279: begin
            cosine_reg0 <= 36'sb11111110100010010011101100011000010;
            sine_reg0   <= 36'sb11011010101101010100111011101101;
        end
        280: begin
            cosine_reg0 <= 36'sb11111110100001101000101011000110101;
            sine_reg0   <= 36'sb11011011011111010011011101100010;
        end
        281: begin
            cosine_reg0 <= 36'sb11111110100000111101100000000001000;
            sine_reg0   <= 36'sb11011100010001010001110110111001;
        end
        282: begin
            cosine_reg0 <= 36'sb11111110100000010010001011000111011;
            sine_reg0   <= 36'sb11011101000011010000000111110000;
        end
        283: begin
            cosine_reg0 <= 36'sb11111110011111100110101100011001110;
            sine_reg0   <= 36'sb11011101110101001110010000000111;
        end
        284: begin
            cosine_reg0 <= 36'sb11111110011110111011000011111000010;
            sine_reg0   <= 36'sb11011110100111001100001111111001;
        end
        285: begin
            cosine_reg0 <= 36'sb11111110011110001111010001100010111;
            sine_reg0   <= 36'sb11011111011001001010000111000111;
        end
        286: begin
            cosine_reg0 <= 36'sb11111110011101100011010101011001100;
            sine_reg0   <= 36'sb11100000001011000111110101101101;
        end
        287: begin
            cosine_reg0 <= 36'sb11111110011100110111001111011100011;
            sine_reg0   <= 36'sb11100000111101000101011011101011;
        end
        288: begin
            cosine_reg0 <= 36'sb11111110011100001010111111101011010;
            sine_reg0   <= 36'sb11100001101111000010111000111101;
        end
        289: begin
            cosine_reg0 <= 36'sb11111110011011011110100110000110100;
            sine_reg0   <= 36'sb11100010100001000000001101100010;
        end
        290: begin
            cosine_reg0 <= 36'sb11111110011010110010000010101101111;
            sine_reg0   <= 36'sb11100011010010111101011001011000;
        end
        291: begin
            cosine_reg0 <= 36'sb11111110011010000101010101100001100;
            sine_reg0   <= 36'sb11100100000100111010011100011110;
        end
        292: begin
            cosine_reg0 <= 36'sb11111110011001011000011110100001100;
            sine_reg0   <= 36'sb11100100110110110111010110110001;
        end
        293: begin
            cosine_reg0 <= 36'sb11111110011000101011011101101101101;
            sine_reg0   <= 36'sb11100101101000110100001000001111;
        end
        294: begin
            cosine_reg0 <= 36'sb11111110010111111110010011000110010;
            sine_reg0   <= 36'sb11100110011010110000110000110110;
        end
        295: begin
            cosine_reg0 <= 36'sb11111110010111010000111110101011001;
            sine_reg0   <= 36'sb11100111001100101101010000100101;
        end
        296: begin
            cosine_reg0 <= 36'sb11111110010110100011100000011100011;
            sine_reg0   <= 36'sb11100111111110101001100111011001;
        end
        297: begin
            cosine_reg0 <= 36'sb11111110010101110101111000011010001;
            sine_reg0   <= 36'sb11101000110000100101110101010001;
        end
        298: begin
            cosine_reg0 <= 36'sb11111110010101001000000110100100010;
            sine_reg0   <= 36'sb11101001100010100001111010001011;
        end
        299: begin
            cosine_reg0 <= 36'sb11111110010100011010001010111010111;
            sine_reg0   <= 36'sb11101010010100011101110110000101;
        end
        300: begin
            cosine_reg0 <= 36'sb11111110010011101100000101011110000;
            sine_reg0   <= 36'sb11101011000110011001101000111100;
        end
        301: begin
            cosine_reg0 <= 36'sb11111110010010111101110110001101101;
            sine_reg0   <= 36'sb11101011111000010101010010101111;
        end
        302: begin
            cosine_reg0 <= 36'sb11111110010010001111011101001001110;
            sine_reg0   <= 36'sb11101100101010010000110011011101;
        end
        303: begin
            cosine_reg0 <= 36'sb11111110010001100000111010010010100;
            sine_reg0   <= 36'sb11101101011100001100001011000010;
        end
        304: begin
            cosine_reg0 <= 36'sb11111110010000110010001101100111111;
            sine_reg0   <= 36'sb11101110001110000111011001011101;
        end
        305: begin
            cosine_reg0 <= 36'sb11111110010000000011010111001001111;
            sine_reg0   <= 36'sb11101111000000000010011110101101;
        end
        306: begin
            cosine_reg0 <= 36'sb11111110001111010100010110111000100;
            sine_reg0   <= 36'sb11101111110001111101011010101111;
        end
        307: begin
            cosine_reg0 <= 36'sb11111110001110100101001100110011110;
            sine_reg0   <= 36'sb11110000100011111000001101100001;
        end
        308: begin
            cosine_reg0 <= 36'sb11111110001101110101111000111011111;
            sine_reg0   <= 36'sb11110001010101110010110111000010;
        end
        309: begin
            cosine_reg0 <= 36'sb11111110001101000110011011010000101;
            sine_reg0   <= 36'sb11110010000111101101010111001111;
        end
        310: begin
            cosine_reg0 <= 36'sb11111110001100010110110011110010010;
            sine_reg0   <= 36'sb11110010111001100111101110000111;
        end
        311: begin
            cosine_reg0 <= 36'sb11111110001011100111000010100000101;
            sine_reg0   <= 36'sb11110011101011100001111011101000;
        end
        312: begin
            cosine_reg0 <= 36'sb11111110001010110111000111011011110;
            sine_reg0   <= 36'sb11110100011101011011111111101111;
        end
        313: begin
            cosine_reg0 <= 36'sb11111110001010000111000010100011111;
            sine_reg0   <= 36'sb11110101001111010101111010011011;
        end
        314: begin
            cosine_reg0 <= 36'sb11111110001001010110110011111000111;
            sine_reg0   <= 36'sb11110110000001001111101011101010;
        end
        315: begin
            cosine_reg0 <= 36'sb11111110001000100110011011011010110;
            sine_reg0   <= 36'sb11110110110011001001010011011010;
        end
        316: begin
            cosine_reg0 <= 36'sb11111110000111110101111001001001100;
            sine_reg0   <= 36'sb11110111100101000010110001101001;
        end
        317: begin
            cosine_reg0 <= 36'sb11111110000111000101001101000101011;
            sine_reg0   <= 36'sb11111000010110111100000110010101;
        end
        318: begin
            cosine_reg0 <= 36'sb11111110000110010100010111001110001;
            sine_reg0   <= 36'sb11111001001000110101010001011101;
        end
        319: begin
            cosine_reg0 <= 36'sb11111110000101100011010111100100000;
            sine_reg0   <= 36'sb11111001111010101110010010111101;
        end
        320: begin
            cosine_reg0 <= 36'sb11111110000100110010001110000110111;
            sine_reg0   <= 36'sb11111010101100100111001010110101;
        end
        321: begin
            cosine_reg0 <= 36'sb11111110000100000000111010110111000;
            sine_reg0   <= 36'sb11111011011110011111111001000011;
        end
        322: begin
            cosine_reg0 <= 36'sb11111110000011001111011101110100001;
            sine_reg0   <= 36'sb11111100010000011000011101100011;
        end
        323: begin
            cosine_reg0 <= 36'sb11111110000010011101110110111110011;
            sine_reg0   <= 36'sb11111101000010010000111000010110;
        end
        324: begin
            cosine_reg0 <= 36'sb11111110000001101100000110010101111;
            sine_reg0   <= 36'sb11111101110100001001001001011000;
        end
        325: begin
            cosine_reg0 <= 36'sb11111110000000111010001011111010100;
            sine_reg0   <= 36'sb11111110100110000001010000101000;
        end
        326: begin
            cosine_reg0 <= 36'sb11111110000000001000000111101100100;
            sine_reg0   <= 36'sb11111111010111111001001110000100;
        end
        327: begin
            cosine_reg0 <= 36'sb11111101111111010101111001101011110;
            sine_reg0   <= 36'sb100000000001001110001000001101001;
        end
        328: begin
            cosine_reg0 <= 36'sb11111101111110100011100001111000010;
            sine_reg0   <= 36'sb100000000111011101000101011010111;
        end
        329: begin
            cosine_reg0 <= 36'sb11111101111101110001000000010010000;
            sine_reg0   <= 36'sb100000001101101100000001011001010;
        end
        330: begin
            cosine_reg0 <= 36'sb11111101111100111110010100111001010;
            sine_reg0   <= 36'sb100000010011111010111100001000010;
        end
        331: begin
            cosine_reg0 <= 36'sb11111101111100001011011111101101111;
            sine_reg0   <= 36'sb100000011010001001110101100111100;
        end
        332: begin
            cosine_reg0 <= 36'sb11111101111011011000100000110000000;
            sine_reg0   <= 36'sb100000100000011000101101110110110;
        end
        333: begin
            cosine_reg0 <= 36'sb11111101111010100101010111111111100;
            sine_reg0   <= 36'sb100000100110100111100100110101111;
        end
        334: begin
            cosine_reg0 <= 36'sb11111101111001110010000101011100011;
            sine_reg0   <= 36'sb100000101100110110011010100100100;
        end
        335: begin
            cosine_reg0 <= 36'sb11111101111000111110101001000111000;
            sine_reg0   <= 36'sb100000110011000101001111000010011;
        end
        336: begin
            cosine_reg0 <= 36'sb11111101111000001011000010111111000;
            sine_reg0   <= 36'sb100000111001010100000010001111100;
        end
        337: begin
            cosine_reg0 <= 36'sb11111101110111010111010011000100101;
            sine_reg0   <= 36'sb100000111111100010110100001011010;
        end
        338: begin
            cosine_reg0 <= 36'sb11111101110110100011011001010111111;
            sine_reg0   <= 36'sb100001000101110001100100110101110;
        end
        339: begin
            cosine_reg0 <= 36'sb11111101110101101111010101111000110;
            sine_reg0   <= 36'sb100001001100000000010100001110100;
        end
        340: begin
            cosine_reg0 <= 36'sb11111101110100111011001000100111011;
            sine_reg0   <= 36'sb100001010010001111000010010101011;
        end
        341: begin
            cosine_reg0 <= 36'sb11111101110100000110110001100011101;
            sine_reg0   <= 36'sb100001011000011101101111001010010;
        end
        342: begin
            cosine_reg0 <= 36'sb11111101110011010010010000101101110;
            sine_reg0   <= 36'sb100001011110101100011010101100101;
        end
        343: begin
            cosine_reg0 <= 36'sb11111101110010011101100110000101100;
            sine_reg0   <= 36'sb100001100100111011000100111100011;
        end
        344: begin
            cosine_reg0 <= 36'sb11111101110001101000110001101011001;
            sine_reg0   <= 36'sb100001101011001001101101111001011;
        end
        345: begin
            cosine_reg0 <= 36'sb11111101110000110011110011011110100;
            sine_reg0   <= 36'sb100001110001011000010101100011010;
        end
        346: begin
            cosine_reg0 <= 36'sb11111101101111111110101011011111110;
            sine_reg0   <= 36'sb100001110111100110111011111001110;
        end
        347: begin
            cosine_reg0 <= 36'sb11111101101111001001011001101111000;
            sine_reg0   <= 36'sb100001111101110101100000111100110;
        end
        348: begin
            cosine_reg0 <= 36'sb11111101101110010011111110001100001;
            sine_reg0   <= 36'sb100010000100000100000100101011111;
        end
        349: begin
            cosine_reg0 <= 36'sb11111101101101011110011000110111010;
            sine_reg0   <= 36'sb100010001010010010100111000111000;
        end
        350: begin
            cosine_reg0 <= 36'sb11111101101100101000101001110000010;
            sine_reg0   <= 36'sb100010010000100001001000001101111;
        end
        351: begin
            cosine_reg0 <= 36'sb11111101101011110010110000110111011;
            sine_reg0   <= 36'sb100010010110101111101000000000001;
        end
        352: begin
            cosine_reg0 <= 36'sb11111101101010111100101110001100100;
            sine_reg0   <= 36'sb100010011100111110000110011101110;
        end
        353: begin
            cosine_reg0 <= 36'sb11111101101010000110100001101111111;
            sine_reg0   <= 36'sb100010100011001100100011100110010;
        end
        354: begin
            cosine_reg0 <= 36'sb11111101101001010000001011100001010;
            sine_reg0   <= 36'sb100010101001011010111111011001100;
        end
        355: begin
            cosine_reg0 <= 36'sb11111101101000011001101011100000110;
            sine_reg0   <= 36'sb100010101111101001011001110111010;
        end
        356: begin
            cosine_reg0 <= 36'sb11111101100111100011000001101110100;
            sine_reg0   <= 36'sb100010110101110111110010111111011;
        end
        357: begin
            cosine_reg0 <= 36'sb11111101100110101100001110001010011;
            sine_reg0   <= 36'sb100010111100000110001010110001011;
        end
        358: begin
            cosine_reg0 <= 36'sb11111101100101110101010000110100101;
            sine_reg0   <= 36'sb100011000010010100100001001101010;
        end
        359: begin
            cosine_reg0 <= 36'sb11111101100100111110001001101101001;
            sine_reg0   <= 36'sb100011001000100010110110010010110;
        end
        360: begin
            cosine_reg0 <= 36'sb11111101100100000110111000110011111;
            sine_reg0   <= 36'sb100011001110110001001010000001100;
        end
        361: begin
            cosine_reg0 <= 36'sb11111101100011001111011110001001001;
            sine_reg0   <= 36'sb100011010100111111011100011001010;
        end
        362: begin
            cosine_reg0 <= 36'sb11111101100010010111111001101100101;
            sine_reg0   <= 36'sb100011011011001101101101011001111;
        end
        363: begin
            cosine_reg0 <= 36'sb11111101100001100000001011011110101;
            sine_reg0   <= 36'sb100011100001011011111101000011001;
        end
        364: begin
            cosine_reg0 <= 36'sb11111101100000101000010011011111001;
            sine_reg0   <= 36'sb100011100111101010001011010100110;
        end
        365: begin
            cosine_reg0 <= 36'sb11111101011111110000010001101110000;
            sine_reg0   <= 36'sb100011101101111000011000001110100;
        end
        366: begin
            cosine_reg0 <= 36'sb11111101011110111000000110001011100;
            sine_reg0   <= 36'sb100011110100000110100011110000000;
        end
        367: begin
            cosine_reg0 <= 36'sb11111101011101111111110000110111100;
            sine_reg0   <= 36'sb100011111010010100101101111001010;
        end
        368: begin
            cosine_reg0 <= 36'sb11111101011101000111010001110010001;
            sine_reg0   <= 36'sb100100000000100010110110101001111;
        end
        369: begin
            cosine_reg0 <= 36'sb11111101011100001110101000111011011;
            sine_reg0   <= 36'sb100100000110110000111110000001101;
        end
        370: begin
            cosine_reg0 <= 36'sb11111101011011010101110110010011010;
            sine_reg0   <= 36'sb100100001100111111000100000000010;
        end
        371: begin
            cosine_reg0 <= 36'sb11111101011010011100111001111001110;
            sine_reg0   <= 36'sb100100010011001101001000100101101;
        end
        372: begin
            cosine_reg0 <= 36'sb11111101011001100011110011101111001;
            sine_reg0   <= 36'sb100100011001011011001011110001011;
        end
        373: begin
            cosine_reg0 <= 36'sb11111101011000101010100011110011001;
            sine_reg0   <= 36'sb100100011111101001001101100011010;
        end
        374: begin
            cosine_reg0 <= 36'sb11111101010111110001001010000110000;
            sine_reg0   <= 36'sb100100100101110111001101111011010;
        end
        375: begin
            cosine_reg0 <= 36'sb11111101010110110111100110100111110;
            sine_reg0   <= 36'sb100100101100000101001100111000111;
        end
        376: begin
            cosine_reg0 <= 36'sb11111101010101111101111001011000010;
            sine_reg0   <= 36'sb100100110010010011001010011100000;
        end
        377: begin
            cosine_reg0 <= 36'sb11111101010101000100000010010111110;
            sine_reg0   <= 36'sb100100111000100001000110100100010;
        end
        378: begin
            cosine_reg0 <= 36'sb11111101010100001010000001100110001;
            sine_reg0   <= 36'sb100100111110101111000001010001101;
        end
        379: begin
            cosine_reg0 <= 36'sb11111101010011001111110111000011100;
            sine_reg0   <= 36'sb100101000100111100111010100011110;
        end
        380: begin
            cosine_reg0 <= 36'sb11111101010010010101100010101111111;
            sine_reg0   <= 36'sb100101001011001010110010011010011;
        end
        381: begin
            cosine_reg0 <= 36'sb11111101010001011011000100101011010;
            sine_reg0   <= 36'sb100101010001011000101000110101010;
        end
        382: begin
            cosine_reg0 <= 36'sb11111101010000100000011100110101110;
            sine_reg0   <= 36'sb100101010111100110011101110100001;
        end
        383: begin
            cosine_reg0 <= 36'sb11111101001111100101101011001111011;
            sine_reg0   <= 36'sb100101011101110100010001010110111;
        end
        384: begin
            cosine_reg0 <= 36'sb11111101001110101010101111111000001;
            sine_reg0   <= 36'sb100101100100000010000011011101001;
        end
        385: begin
            cosine_reg0 <= 36'sb11111101001101101111101010110000001;
            sine_reg0   <= 36'sb100101101010001111110100000110101;
        end
        386: begin
            cosine_reg0 <= 36'sb11111101001100110100011011110111010;
            sine_reg0   <= 36'sb100101110000011101100011010011011;
        end
        387: begin
            cosine_reg0 <= 36'sb11111101001011111001000011001101101;
            sine_reg0   <= 36'sb100101110110101011010001000010111;
        end
        388: begin
            cosine_reg0 <= 36'sb11111101001010111101100000110011011;
            sine_reg0   <= 36'sb100101111100111000111101010101000;
        end
        389: begin
            cosine_reg0 <= 36'sb11111101001010000001110100101000011;
            sine_reg0   <= 36'sb100110000011000110101000001001011;
        end
        390: begin
            cosine_reg0 <= 36'sb11111101001001000101111110101100110;
            sine_reg0   <= 36'sb100110001001010100010001100000000;
        end
        391: begin
            cosine_reg0 <= 36'sb11111101001000001001111111000000100;
            sine_reg0   <= 36'sb100110001111100001111001011000011;
        end
        392: begin
            cosine_reg0 <= 36'sb11111101000111001101110101100011110;
            sine_reg0   <= 36'sb100110010101101111011111110010100;
        end
        393: begin
            cosine_reg0 <= 36'sb11111101000110010001100010010110011;
            sine_reg0   <= 36'sb100110011011111101000100101110000;
        end
        394: begin
            cosine_reg0 <= 36'sb11111101000101010101000101011000100;
            sine_reg0   <= 36'sb100110100010001010101000001010101;
        end
        395: begin
            cosine_reg0 <= 36'sb11111101000100011000011110101010010;
            sine_reg0   <= 36'sb100110101000011000001010001000010;
        end
        396: begin
            cosine_reg0 <= 36'sb11111101000011011011101110001011101;
            sine_reg0   <= 36'sb100110101110100101101010100110100;
        end
        397: begin
            cosine_reg0 <= 36'sb11111101000010011110110011111100100;
            sine_reg0   <= 36'sb100110110100110011001001100101010;
        end
        398: begin
            cosine_reg0 <= 36'sb11111101000001100001101111111101001;
            sine_reg0   <= 36'sb100110111011000000100111000100001;
        end
        399: begin
            cosine_reg0 <= 36'sb11111101000000100100100010001101011;
            sine_reg0   <= 36'sb100111000001001110000011000011000;
        end
        400: begin
            cosine_reg0 <= 36'sb11111100111111100111001010101101010;
            sine_reg0   <= 36'sb100111000111011011011101100001101;
        end
        401: begin
            cosine_reg0 <= 36'sb11111100111110101001101001011101000;
            sine_reg0   <= 36'sb100111001101101000110110011111101;
        end
        402: begin
            cosine_reg0 <= 36'sb11111100111101101011111110011100101;
            sine_reg0   <= 36'sb100111010011110110001101111101000;
        end
        403: begin
            cosine_reg0 <= 36'sb11111100111100101110001001101100000;
            sine_reg0   <= 36'sb100111011010000011100011111001011;
        end
        404: begin
            cosine_reg0 <= 36'sb11111100111011110000001011001011010;
            sine_reg0   <= 36'sb100111100000010000111000010100011;
        end
        405: begin
            cosine_reg0 <= 36'sb11111100111010110010000010111010011;
            sine_reg0   <= 36'sb100111100110011110001011001110000;
        end
        406: begin
            cosine_reg0 <= 36'sb11111100111001110011110000111001100;
            sine_reg0   <= 36'sb100111101100101011011100100110000;
        end
        407: begin
            cosine_reg0 <= 36'sb11111100111000110101010101001000101;
            sine_reg0   <= 36'sb100111110010111000101100011011111;
        end
        408: begin
            cosine_reg0 <= 36'sb11111100110111110110101111100111110;
            sine_reg0   <= 36'sb100111111001000101111010101111110;
        end
        409: begin
            cosine_reg0 <= 36'sb11111100110110111000000000010110111;
            sine_reg0   <= 36'sb100111111111010011000111100001000;
        end
        410: begin
            cosine_reg0 <= 36'sb11111100110101111001000111010110010;
            sine_reg0   <= 36'sb101000000101100000010010101111110;
        end
        411: begin
            cosine_reg0 <= 36'sb11111100110100111010000100100101101;
            sine_reg0   <= 36'sb101000001011101101011100011011100;
        end
        412: begin
            cosine_reg0 <= 36'sb11111100110011111010111000000101010;
            sine_reg0   <= 36'sb101000010001111010100100100100001;
        end
        413: begin
            cosine_reg0 <= 36'sb11111100110010111011100001110101000;
            sine_reg0   <= 36'sb101000011000000111101011001001011;
        end
        414: begin
            cosine_reg0 <= 36'sb11111100110001111100000001110101001;
            sine_reg0   <= 36'sb101000011110010100110000001010111;
        end
        415: begin
            cosine_reg0 <= 36'sb11111100110000111100011000000101100;
            sine_reg0   <= 36'sb101000100100100001110011101000101;
        end
        416: begin
            cosine_reg0 <= 36'sb11111100101111111100100100100110001;
            sine_reg0   <= 36'sb101000101010101110110101100010010;
        end
        417: begin
            cosine_reg0 <= 36'sb11111100101110111100100111010111010;
            sine_reg0   <= 36'sb101000110000111011110101110111101;
        end
        418: begin
            cosine_reg0 <= 36'sb11111100101101111100100000011000101;
            sine_reg0   <= 36'sb101000110111001000110100101000010;
        end
        419: begin
            cosine_reg0 <= 36'sb11111100101100111100001111101010100;
            sine_reg0   <= 36'sb101000111101010101110001110100010;
        end
        420: begin
            cosine_reg0 <= 36'sb11111100101011111011110101001100111;
            sine_reg0   <= 36'sb101001000011100010101101011011000;
        end
        421: begin
            cosine_reg0 <= 36'sb11111100101010111011010000111111111;
            sine_reg0   <= 36'sb101001001001101111100111011100100;
        end
        422: begin
            cosine_reg0 <= 36'sb11111100101001111010100011000011010;
            sine_reg0   <= 36'sb101001001111111100011111111000100;
        end
        423: begin
            cosine_reg0 <= 36'sb11111100101000111001101011010111011;
            sine_reg0   <= 36'sb101001010110001001010110101110110;
        end
        424: begin
            cosine_reg0 <= 36'sb11111100100111111000101001111100000;
            sine_reg0   <= 36'sb101001011100010110001011111110111;
        end
        425: begin
            cosine_reg0 <= 36'sb11111100100110110111011110110001011;
            sine_reg0   <= 36'sb101001100010100010111111101000111;
        end
        426: begin
            cosine_reg0 <= 36'sb11111100100101110110001001110111100;
            sine_reg0   <= 36'sb101001101000101111110001101100010;
        end
        427: begin
            cosine_reg0 <= 36'sb11111100100100110100101011001110011;
            sine_reg0   <= 36'sb101001101110111100100010001001000;
        end
        428: begin
            cosine_reg0 <= 36'sb11111100100011110011000010110110000;
            sine_reg0   <= 36'sb101001110101001001010000111110110;
        end
        429: begin
            cosine_reg0 <= 36'sb11111100100010110001010000101110100;
            sine_reg0   <= 36'sb101001111011010101111110001101010;
        end
        430: begin
            cosine_reg0 <= 36'sb11111100100001101111010100110111111;
            sine_reg0   <= 36'sb101010000001100010101001110100011;
        end
        431: begin
            cosine_reg0 <= 36'sb11111100100000101101001111010010001;
            sine_reg0   <= 36'sb101010000111101111010011110011110;
        end
        432: begin
            cosine_reg0 <= 36'sb11111100011111101010111111111101011;
            sine_reg0   <= 36'sb101010001101111011111100001011001;
        end
        433: begin
            cosine_reg0 <= 36'sb11111100011110101000100110111001100;
            sine_reg0   <= 36'sb101010010100001000100010111010100;
        end
        434: begin
            cosine_reg0 <= 36'sb11111100011101100110000100000110110;
            sine_reg0   <= 36'sb101010011010010101001000000001011;
        end
        435: begin
            cosine_reg0 <= 36'sb11111100011100100011010111100101001;
            sine_reg0   <= 36'sb101010100000100001101011011111100;
        end
        436: begin
            cosine_reg0 <= 36'sb11111100011011100000100001010100100;
            sine_reg0   <= 36'sb101010100110101110001101010100111;
        end
        437: begin
            cosine_reg0 <= 36'sb11111100011010011101100001010101001;
            sine_reg0   <= 36'sb101010101100111010101101100001001;
        end
        438: begin
            cosine_reg0 <= 36'sb11111100011001011010010111100110111;
            sine_reg0   <= 36'sb101010110011000111001100000100000;
        end
        439: begin
            cosine_reg0 <= 36'sb11111100011000010111000100001001111;
            sine_reg0   <= 36'sb101010111001010011101000111101010;
        end
        440: begin
            cosine_reg0 <= 36'sb11111100010111010011100110111110010;
            sine_reg0   <= 36'sb101010111111100000000100001100101;
        end
        441: begin
            cosine_reg0 <= 36'sb11111100010110010000000000000011111;
            sine_reg0   <= 36'sb101011000101101100011101110010000;
        end
        442: begin
            cosine_reg0 <= 36'sb11111100010101001100001111011010110;
            sine_reg0   <= 36'sb101011001011111000110101101101000;
        end
        443: begin
            cosine_reg0 <= 36'sb11111100010100001000010101000011001;
            sine_reg0   <= 36'sb101011010010000101001011111101100;
        end
        444: begin
            cosine_reg0 <= 36'sb11111100010011000100010000111101000;
            sine_reg0   <= 36'sb101011011000010001100000100011001;
        end
        445: begin
            cosine_reg0 <= 36'sb11111100010010000000000011001000010;
            sine_reg0   <= 36'sb101011011110011101110011011101110;
        end
        446: begin
            cosine_reg0 <= 36'sb11111100010000111011101011100101001;
            sine_reg0   <= 36'sb101011100100101010000100101101001;
        end
        447: begin
            cosine_reg0 <= 36'sb11111100001111110111001010010011100;
            sine_reg0   <= 36'sb101011101010110110010100010001000;
        end
        448: begin
            cosine_reg0 <= 36'sb11111100001110110010011111010011011;
            sine_reg0   <= 36'sb101011110001000010100010001001001;
        end
        449: begin
            cosine_reg0 <= 36'sb11111100001101101101101010100101000;
            sine_reg0   <= 36'sb101011110111001110101110010101001;
        end
        450: begin
            cosine_reg0 <= 36'sb11111100001100101000101100001000011;
            sine_reg0   <= 36'sb101011111101011010111000110101000;
        end
        451: begin
            cosine_reg0 <= 36'sb11111100001011100011100011111101011;
            sine_reg0   <= 36'sb101100000011100111000001101000100;
        end
        452: begin
            cosine_reg0 <= 36'sb11111100001010011110010010000100001;
            sine_reg0   <= 36'sb101100001001110011001000101111001;
        end
        453: begin
            cosine_reg0 <= 36'sb11111100001001011000110110011100110;
            sine_reg0   <= 36'sb101100001111111111001110001001000;
        end
        454: begin
            cosine_reg0 <= 36'sb11111100001000010011010001000111010;
            sine_reg0   <= 36'sb101100010110001011010001110101100;
        end
        455: begin
            cosine_reg0 <= 36'sb11111100000111001101100010000011101;
            sine_reg0   <= 36'sb101100011100010111010011110100110;
        end
        456: begin
            cosine_reg0 <= 36'sb11111100000110000111101001010001111;
            sine_reg0   <= 36'sb101100100010100011010100000110010;
        end
        457: begin
            cosine_reg0 <= 36'sb11111100000101000001100110110010001;
            sine_reg0   <= 36'sb101100101000101111010010101001111;
        end
        458: begin
            cosine_reg0 <= 36'sb11111100000011111011011010100100100;
            sine_reg0   <= 36'sb101100101110111011001111011111010;
        end
        459: begin
            cosine_reg0 <= 36'sb11111100000010110101000100101000111;
            sine_reg0   <= 36'sb101100110101000111001010100110011;
        end
        460: begin
            cosine_reg0 <= 36'sb11111100000001101110100100111111010;
            sine_reg0   <= 36'sb101100111011010011000011111110111;
        end
        461: begin
            cosine_reg0 <= 36'sb11111100000000100111111011100111111;
            sine_reg0   <= 36'sb101101000001011110111011101000100;
        end
        462: begin
            cosine_reg0 <= 36'sb11111011111111100001001000100010110;
            sine_reg0   <= 36'sb101101000111101010110001100011000;
        end
        463: begin
            cosine_reg0 <= 36'sb11111011111110011010001011101111110;
            sine_reg0   <= 36'sb101101001101110110100101101110010;
        end
        464: begin
            cosine_reg0 <= 36'sb11111011111101010011000101001111001;
            sine_reg0   <= 36'sb101101010100000010011000001001111;
        end
        465: begin
            cosine_reg0 <= 36'sb11111011111100001011110101000000110;
            sine_reg0   <= 36'sb101101011010001110001000110101110;
        end
        466: begin
            cosine_reg0 <= 36'sb11111011111011000100011011000100110;
            sine_reg0   <= 36'sb101101100000011001110111110001100;
        end
        467: begin
            cosine_reg0 <= 36'sb11111011111001111100110111011011001;
            sine_reg0   <= 36'sb101101100110100101100100111101000;
        end
        468: begin
            cosine_reg0 <= 36'sb11111011111000110101001010000100000;
            sine_reg0   <= 36'sb101101101100110001010000011000000;
        end
        469: begin
            cosine_reg0 <= 36'sb11111011110111101101010010111111010;
            sine_reg0   <= 36'sb101101110010111100111010000010010;
        end
        470: begin
            cosine_reg0 <= 36'sb11111011110110100101010010001101001;
            sine_reg0   <= 36'sb101101111001001000100001111011100;
        end
        471: begin
            cosine_reg0 <= 36'sb11111011110101011101000111101101101;
            sine_reg0   <= 36'sb101101111111010100001000000011100;
        end
        472: begin
            cosine_reg0 <= 36'sb11111011110100010100110011100000110;
            sine_reg0   <= 36'sb101110000101011111101100011010000;
        end
        473: begin
            cosine_reg0 <= 36'sb11111011110011001100010101100110011;
            sine_reg0   <= 36'sb101110001011101011001110111110111;
        end
        474: begin
            cosine_reg0 <= 36'sb11111011110010000011101101111110111;
            sine_reg0   <= 36'sb101110010001110110101111110001110;
        end
        475: begin
            cosine_reg0 <= 36'sb11111011110000111010111100101010001;
            sine_reg0   <= 36'sb101110011000000010001110110010011;
        end
        476: begin
            cosine_reg0 <= 36'sb11111011101111110010000001101000001;
            sine_reg0   <= 36'sb101110011110001101101100000000101;
        end
        477: begin
            cosine_reg0 <= 36'sb11111011101110101000111100111000111;
            sine_reg0   <= 36'sb101110100100011001000111011100010;
        end
        478: begin
            cosine_reg0 <= 36'sb11111011101101011111101110011100101;
            sine_reg0   <= 36'sb101110101010100100100001000100111;
        end
        479: begin
            cosine_reg0 <= 36'sb11111011101100010110010110010011010;
            sine_reg0   <= 36'sb101110110000101111111000111010100;
        end
        480: begin
            cosine_reg0 <= 36'sb11111011101011001100110100011100111;
            sine_reg0   <= 36'sb101110110110111011001110111100101;
        end
        481: begin
            cosine_reg0 <= 36'sb11111011101010000011001000111001100;
            sine_reg0   <= 36'sb101110111101000110100011001011001;
        end
        482: begin
            cosine_reg0 <= 36'sb11111011101000111001010011101001010;
            sine_reg0   <= 36'sb101111000011010001110101100101111;
        end
        483: begin
            cosine_reg0 <= 36'sb11111011100111101111010100101100000;
            sine_reg0   <= 36'sb101111001001011101000110001100011;
        end
        484: begin
            cosine_reg0 <= 36'sb11111011100110100101001100000010000;
            sine_reg0   <= 36'sb101111001111101000010100111110101;
        end
        485: begin
            cosine_reg0 <= 36'sb11111011100101011010111001101011001;
            sine_reg0   <= 36'sb101111010101110011100001111100011;
        end
        486: begin
            cosine_reg0 <= 36'sb11111011100100010000011101100111100;
            sine_reg0   <= 36'sb101111011011111110101101000101010;
        end
        487: begin
            cosine_reg0 <= 36'sb11111011100011000101110111110111010;
            sine_reg0   <= 36'sb101111100010001001110110011001001;
        end
        488: begin
            cosine_reg0 <= 36'sb11111011100001111011001000011010010;
            sine_reg0   <= 36'sb101111101000010100111101110111101;
        end
        489: begin
            cosine_reg0 <= 36'sb11111011100000110000001111010000101;
            sine_reg0   <= 36'sb101111101110100000000011100000101;
        end
        490: begin
            cosine_reg0 <= 36'sb11111011011111100101001100011010011;
            sine_reg0   <= 36'sb101111110100101011000111010011111;
        end
        491: begin
            cosine_reg0 <= 36'sb11111011011110011001111111110111101;
            sine_reg0   <= 36'sb101111111010110110001001010001001;
        end
        492: begin
            cosine_reg0 <= 36'sb11111011011101001110101001101000100;
            sine_reg0   <= 36'sb110000000001000001001001011000010;
        end
        493: begin
            cosine_reg0 <= 36'sb11111011011100000011001001101100110;
            sine_reg0   <= 36'sb110000000111001100000111101000110;
        end
        494: begin
            cosine_reg0 <= 36'sb11111011011010110111100000000100110;
            sine_reg0   <= 36'sb110000001101010111000100000010101;
        end
        495: begin
            cosine_reg0 <= 36'sb11111011011001101011101100110000010;
            sine_reg0   <= 36'sb110000010011100001111110100101100;
        end
        496: begin
            cosine_reg0 <= 36'sb11111011011000011111101111101111100;
            sine_reg0   <= 36'sb110000011001101100110111010001010;
        end
        497: begin
            cosine_reg0 <= 36'sb11111011010111010011101001000010101;
            sine_reg0   <= 36'sb110000011111110111101110000101100;
        end
        498: begin
            cosine_reg0 <= 36'sb11111011010110000111011000101001011;
            sine_reg0   <= 36'sb110000100110000010100011000010001;
        end
        499: begin
            cosine_reg0 <= 36'sb11111011010100111010111110100100000;
            sine_reg0   <= 36'sb110000101100001101010110000110110;
        end
        500: begin
            cosine_reg0 <= 36'sb11111011010011101110011010110010100;
            sine_reg0   <= 36'sb110000110010011000000111010011011;
        end
        501: begin
            cosine_reg0 <= 36'sb11111011010010100001101101010100111;
            sine_reg0   <= 36'sb110000111000100010110110100111101;
        end
        502: begin
            cosine_reg0 <= 36'sb11111011010001010100110110001011010;
            sine_reg0   <= 36'sb110000111110101101100100000011001;
        end
        503: begin
            cosine_reg0 <= 36'sb11111011010000000111110101010101101;
            sine_reg0   <= 36'sb110001000100111000001111100101111;
        end
        504: begin
            cosine_reg0 <= 36'sb11111011001110111010101010110100001;
            sine_reg0   <= 36'sb110001001011000010111001001111100;
        end
        505: begin
            cosine_reg0 <= 36'sb11111011001101101101010110100110110;
            sine_reg0   <= 36'sb110001010001001101100000111111111;
        end
        506: begin
            cosine_reg0 <= 36'sb11111011001100011111111000101101011;
            sine_reg0   <= 36'sb110001010111011000000110110110100;
        end
        507: begin
            cosine_reg0 <= 36'sb11111011001011010010010001001000011;
            sine_reg0   <= 36'sb110001011101100010101010110011100;
        end
        508: begin
            cosine_reg0 <= 36'sb11111011001010000100011111110111100;
            sine_reg0   <= 36'sb110001100011101101001100110110011;
        end
        509: begin
            cosine_reg0 <= 36'sb11111011001000110110100100111011000;
            sine_reg0   <= 36'sb110001101001110111101100111111000;
        end
        510: begin
            cosine_reg0 <= 36'sb11111011000111101000100000010010110;
            sine_reg0   <= 36'sb110001110000000010001011001101001;
        end
        511: begin
            cosine_reg0 <= 36'sb11111011000110011010010001111111000;
            sine_reg0   <= 36'sb110001110110001100100111100000100;
        end
        512: begin
            cosine_reg0 <= 36'sb11111011000101001011111001111111101;
            sine_reg0   <= 36'sb110001111100010111000001111000110;
        end
        513: begin
            cosine_reg0 <= 36'sb11111011000011111101011000010100110;
            sine_reg0   <= 36'sb110010000010100001011010010101111;
        end
        514: begin
            cosine_reg0 <= 36'sb11111011000010101110101100111110011;
            sine_reg0   <= 36'sb110010001000101011110000110111101;
        end
        515: begin
            cosine_reg0 <= 36'sb11111011000001011111110111111100101;
            sine_reg0   <= 36'sb110010001110110110000101011101100;
        end
        516: begin
            cosine_reg0 <= 36'sb11111011000000010000111001001111011;
            sine_reg0   <= 36'sb110010010101000000011000000111100;
        end
        517: begin
            cosine_reg0 <= 36'sb11111010111111000001110000110110111;
            sine_reg0   <= 36'sb110010011011001010101000110101011;
        end
        518: begin
            cosine_reg0 <= 36'sb11111010111101110010011110110011001;
            sine_reg0   <= 36'sb110010100001010100110111100110110;
        end
        519: begin
            cosine_reg0 <= 36'sb11111010111100100011000011000100001;
            sine_reg0   <= 36'sb110010100111011111000100011011100;
        end
        520: begin
            cosine_reg0 <= 36'sb11111010111011010011011101101010000;
            sine_reg0   <= 36'sb110010101101101001001111010011011;
        end
        521: begin
            cosine_reg0 <= 36'sb11111010111010000011101110100100101;
            sine_reg0   <= 36'sb110010110011110011011000001110001;
        end
        522: begin
            cosine_reg0 <= 36'sb11111010111000110011110101110100010;
            sine_reg0   <= 36'sb110010111001111101011111001011100;
        end
        523: begin
            cosine_reg0 <= 36'sb11111010110111100011110011011000110;
            sine_reg0   <= 36'sb110011000000000111100100001011010;
        end
        524: begin
            cosine_reg0 <= 36'sb11111010110110010011100111010010011;
            sine_reg0   <= 36'sb110011000110010001100111001101001;
        end
        525: begin
            cosine_reg0 <= 36'sb11111010110101000011010001100001000;
            sine_reg0   <= 36'sb110011001100011011101000010001000;
        end
        526: begin
            cosine_reg0 <= 36'sb11111010110011110010110010000100110;
            sine_reg0   <= 36'sb110011010010100101100111010110100;
        end
        527: begin
            cosine_reg0 <= 36'sb11111010110010100010001000111101101;
            sine_reg0   <= 36'sb110011011000101111100100011101100;
        end
        528: begin
            cosine_reg0 <= 36'sb11111010110001010001010110001011101;
            sine_reg0   <= 36'sb110011011110111001011111100101110;
        end
        529: begin
            cosine_reg0 <= 36'sb11111010110000000000011001101111000;
            sine_reg0   <= 36'sb110011100101000011011000101110111;
        end
        530: begin
            cosine_reg0 <= 36'sb11111010101110101111010011100111101;
            sine_reg0   <= 36'sb110011101011001101001111111000110;
        end
        531: begin
            cosine_reg0 <= 36'sb11111010101101011110000011110101101;
            sine_reg0   <= 36'sb110011110001010111000101000011001;
        end
        532: begin
            cosine_reg0 <= 36'sb11111010101100001100101010011000111;
            sine_reg0   <= 36'sb110011110111100000111000001101110;
        end
        533: begin
            cosine_reg0 <= 36'sb11111010101010111011000111010001110;
            sine_reg0   <= 36'sb110011111101101010101001011000011;
        end
        534: begin
            cosine_reg0 <= 36'sb11111010101001101001011010100000000;
            sine_reg0   <= 36'sb110100000011110100011000100010111;
        end
        535: begin
            cosine_reg0 <= 36'sb11111010101000010111100100000011111;
            sine_reg0   <= 36'sb110100001001111110000101101100111;
        end
        536: begin
            cosine_reg0 <= 36'sb11111010100111000101100011111101011;
            sine_reg0   <= 36'sb110100010000000111110000110110001;
        end
        537: begin
            cosine_reg0 <= 36'sb11111010100101110011011010001100100;
            sine_reg0   <= 36'sb110100010110010001011001111110100;
        end
        538: begin
            cosine_reg0 <= 36'sb11111010100100100001000110110001010;
            sine_reg0   <= 36'sb110100011100011011000001000101110;
        end
        539: begin
            cosine_reg0 <= 36'sb11111010100011001110101001101011110;
            sine_reg0   <= 36'sb110100100010100100100110001011101;
        end
        540: begin
            cosine_reg0 <= 36'sb11111010100001111100000010111100000;
            sine_reg0   <= 36'sb110100101000101110001001001111110;
        end
        541: begin
            cosine_reg0 <= 36'sb11111010100000101001010010100010010;
            sine_reg0   <= 36'sb110100101110110111101010010010000;
        end
        542: begin
            cosine_reg0 <= 36'sb11111010011111010110011000011110010;
            sine_reg0   <= 36'sb110100110101000001001001010010010;
        end
        543: begin
            cosine_reg0 <= 36'sb11111010011110000011010100110000010;
            sine_reg0   <= 36'sb110100111011001010100110010000001;
        end
        544: begin
            cosine_reg0 <= 36'sb11111010011100110000000111011000010;
            sine_reg0   <= 36'sb110101000001010100000001001011011;
        end
        545: begin
            cosine_reg0 <= 36'sb11111010011011011100110000010110010;
            sine_reg0   <= 36'sb110101000111011101011010000011110;
        end
        546: begin
            cosine_reg0 <= 36'sb11111010011010001001001111101010011;
            sine_reg0   <= 36'sb110101001101100110110000111001001;
        end
        547: begin
            cosine_reg0 <= 36'sb11111010011000110101100101010100101;
            sine_reg0   <= 36'sb110101010011110000000101101011010;
        end
        548: begin
            cosine_reg0 <= 36'sb11111010010111100001110001010101000;
            sine_reg0   <= 36'sb110101011001111001011000011001110;
        end
        549: begin
            cosine_reg0 <= 36'sb11111010010110001101110011101011110;
            sine_reg0   <= 36'sb110101100000000010101001000100100;
        end
        550: begin
            cosine_reg0 <= 36'sb11111010010100111001101100011000110;
            sine_reg0   <= 36'sb110101100110001011110111101011011;
        end
        551: begin
            cosine_reg0 <= 36'sb11111010010011100101011011011100000;
            sine_reg0   <= 36'sb110101101100010101000100001101111;
        end
        552: begin
            cosine_reg0 <= 36'sb11111010010010010001000000110101110;
            sine_reg0   <= 36'sb110101110010011110001110101011111;
        end
        553: begin
            cosine_reg0 <= 36'sb11111010010000111100011100100110000;
            sine_reg0   <= 36'sb110101111000100111010111000101010;
        end
        554: begin
            cosine_reg0 <= 36'sb11111010001111100111101110101100101;
            sine_reg0   <= 36'sb110101111110110000011101011001101;
        end
        555: begin
            cosine_reg0 <= 36'sb11111010001110010010110111001001110;
            sine_reg0   <= 36'sb110110000100111001100001101000110;
        end
        556: begin
            cosine_reg0 <= 36'sb11111010001100111101110101111101101;
            sine_reg0   <= 36'sb110110001011000010100011110010100;
        end
        557: begin
            cosine_reg0 <= 36'sb11111010001011101000101011001000001;
            sine_reg0   <= 36'sb110110010001001011100011110110101;
        end
        558: begin
            cosine_reg0 <= 36'sb11111010001010010011010110101001010;
            sine_reg0   <= 36'sb110110010111010100100001110100110;
        end
        559: begin
            cosine_reg0 <= 36'sb11111010001000111101111000100001001;
            sine_reg0   <= 36'sb110110011101011101011101101100110;
        end
        560: begin
            cosine_reg0 <= 36'sb11111010000111101000010000101111111;
            sine_reg0   <= 36'sb110110100011100110010111011110100;
        end
        561: begin
            cosine_reg0 <= 36'sb11111010000110010010011111010101011;
            sine_reg0   <= 36'sb110110101001101111001111001001100;
        end
        562: begin
            cosine_reg0 <= 36'sb11111010000100111100100100010001111;
            sine_reg0   <= 36'sb110110101111111000000100101101110;
        end
        563: begin
            cosine_reg0 <= 36'sb11111010000011100110011111100101011;
            sine_reg0   <= 36'sb110110110110000000111000001010111;
        end
        564: begin
            cosine_reg0 <= 36'sb11111010000010010000010001001111110;
            sine_reg0   <= 36'sb110110111100001001101001100000101;
        end
        565: begin
            cosine_reg0 <= 36'sb11111010000000111001111001010001011;
            sine_reg0   <= 36'sb110111000010010010011000101110111;
        end
        566: begin
            cosine_reg0 <= 36'sb11111001111111100011010111101010000;
            sine_reg0   <= 36'sb110111001000011011000101110101010;
        end
        567: begin
            cosine_reg0 <= 36'sb11111001111110001100101100011001110;
            sine_reg0   <= 36'sb110111001110100011110000110011110;
        end
        568: begin
            cosine_reg0 <= 36'sb11111001111100110101110111100000110;
            sine_reg0   <= 36'sb110111010100101100011001101001111;
        end
        569: begin
            cosine_reg0 <= 36'sb11111001111011011110111000111111000;
            sine_reg0   <= 36'sb110111011010110101000000010111100;
        end
        570: begin
            cosine_reg0 <= 36'sb11111001111010000111110000110100101;
            sine_reg0   <= 36'sb110111100000111101100100111100011;
        end
        571: begin
            cosine_reg0 <= 36'sb11111001111000110000011111000001101;
            sine_reg0   <= 36'sb110111100111000110000111011000010;
        end
        572: begin
            cosine_reg0 <= 36'sb11111001110111011001000011100110000;
            sine_reg0   <= 36'sb110111101101001110100111101011000;
        end
        573: begin
            cosine_reg0 <= 36'sb11111001110110000001011110100001111;
            sine_reg0   <= 36'sb110111110011010111000101110100010;
        end
        574: begin
            cosine_reg0 <= 36'sb11111001110100101001101111110101011;
            sine_reg0   <= 36'sb110111111001011111100001110011111;
        end
        575: begin
            cosine_reg0 <= 36'sb11111001110011010001110111100000011;
            sine_reg0   <= 36'sb110111111111100111111011101001100;
        end
        576: begin
            cosine_reg0 <= 36'sb11111001110001111001110101100011000;
            sine_reg0   <= 36'sb111000000101110000010011010101000;
        end
        577: begin
            cosine_reg0 <= 36'sb11111001110000100001101001111101011;
            sine_reg0   <= 36'sb111000001011111000101000110110000;
        end
        578: begin
            cosine_reg0 <= 36'sb11111001101111001001010100101111100;
            sine_reg0   <= 36'sb111000010010000000111100001100100;
        end
        579: begin
            cosine_reg0 <= 36'sb11111001101101110000110101111001011;
            sine_reg0   <= 36'sb111000011000001001001101011000001;
        end
        580: begin
            cosine_reg0 <= 36'sb11111001101100011000001101011011001;
            sine_reg0   <= 36'sb111000011110010001011100011000101;
        end
        581: begin
            cosine_reg0 <= 36'sb11111001101010111111011011010100110;
            sine_reg0   <= 36'sb111000100100011001101001001101110;
        end
        582: begin
            cosine_reg0 <= 36'sb11111001101001100110011111100110011;
            sine_reg0   <= 36'sb111000101010100001110011110111010;
        end
        583: begin
            cosine_reg0 <= 36'sb11111001101000001101011010010000000;
            sine_reg0   <= 36'sb111000110000101001111100010101000;
        end
        584: begin
            cosine_reg0 <= 36'sb11111001100110110100001011010001110;
            sine_reg0   <= 36'sb111000110110110010000010100110110;
        end
        585: begin
            cosine_reg0 <= 36'sb11111001100101011010110010101011100;
            sine_reg0   <= 36'sb111000111100111010000110101100001;
        end
        586: begin
            cosine_reg0 <= 36'sb11111001100100000001010000011101100;
            sine_reg0   <= 36'sb111001000011000010001000100101000;
        end
        587: begin
            cosine_reg0 <= 36'sb11111001100010100111100100100111110;
            sine_reg0   <= 36'sb111001001001001010001000010001001;
        end
        588: begin
            cosine_reg0 <= 36'sb11111001100001001101101111001010010;
            sine_reg0   <= 36'sb111001001111010010000101110000010;
        end
        589: begin
            cosine_reg0 <= 36'sb11111001011111110011110000000101001;
            sine_reg0   <= 36'sb111001010101011010000001000010001;
        end
        590: begin
            cosine_reg0 <= 36'sb11111001011110011001100111011000010;
            sine_reg0   <= 36'sb111001011011100001111010000110101;
        end
        591: begin
            cosine_reg0 <= 36'sb11111001011100111111010101000100000;
            sine_reg0   <= 36'sb111001100001101001110000111101011;
        end
        592: begin
            cosine_reg0 <= 36'sb11111001011011100100111001001000001;
            sine_reg0   <= 36'sb111001100111110001100101100110001;
        end
        593: begin
            cosine_reg0 <= 36'sb11111001011010001010010011100100111;
            sine_reg0   <= 36'sb111001101101111001011000000000110;
        end
        594: begin
            cosine_reg0 <= 36'sb11111001011000101111100100011010010;
            sine_reg0   <= 36'sb111001110100000001001000001101000;
        end
        595: begin
            cosine_reg0 <= 36'sb11111001010111010100101011101000010;
            sine_reg0   <= 36'sb111001111010001000110110001010100;
        end
        596: begin
            cosine_reg0 <= 36'sb11111001010101111001101001001110111;
            sine_reg0   <= 36'sb111010000000010000100001111001001;
        end
        597: begin
            cosine_reg0 <= 36'sb11111001010100011110011101001110011;
            sine_reg0   <= 36'sb111010000110011000001011011000110;
        end
        598: begin
            cosine_reg0 <= 36'sb11111001010011000011000111100110110;
            sine_reg0   <= 36'sb111010001100011111110010101000111;
        end
        599: begin
            cosine_reg0 <= 36'sb11111001010001100111101000010111111;
            sine_reg0   <= 36'sb111010010010100111010111101001100;
        end
        600: begin
            cosine_reg0 <= 36'sb11111001010000001011111111100010001;
            sine_reg0   <= 36'sb111010011000101110111010011010011;
        end
        601: begin
            cosine_reg0 <= 36'sb11111001001110110000001101000101010;
            sine_reg0   <= 36'sb111010011110110110011010111011000;
        end
        602: begin
            cosine_reg0 <= 36'sb11111001001101010100010001000001011;
            sine_reg0   <= 36'sb111010100100111101111001001011100;
        end
        603: begin
            cosine_reg0 <= 36'sb11111001001011111000001011010110101;
            sine_reg0   <= 36'sb111010101011000101010101001011011;
        end
        604: begin
            cosine_reg0 <= 36'sb11111001001010011011111100000101001;
            sine_reg0   <= 36'sb111010110001001100101110111010100;
        end
        605: begin
            cosine_reg0 <= 36'sb11111001001000111111100011001100110;
            sine_reg0   <= 36'sb111010110111010100000110011000101;
        end
        606: begin
            cosine_reg0 <= 36'sb11111001000111100011000000101101101;
            sine_reg0   <= 36'sb111010111101011011011011100101100;
        end
        607: begin
            cosine_reg0 <= 36'sb11111001000110000110010100101000000;
            sine_reg0   <= 36'sb111011000011100010101110100000111;
        end
        608: begin
            cosine_reg0 <= 36'sb11111001000100101001011110111011101;
            sine_reg0   <= 36'sb111011001001101001111111001010100;
        end
        609: begin
            cosine_reg0 <= 36'sb11111001000011001100011111101000101;
            sine_reg0   <= 36'sb111011001111110001001101100010010;
        end
        610: begin
            cosine_reg0 <= 36'sb11111001000001101111010110101111010;
            sine_reg0   <= 36'sb111011010101111000011001100111110;
        end
        611: begin
            cosine_reg0 <= 36'sb11111001000000010010000100001111011;
            sine_reg0   <= 36'sb111011011011111111100011011010111;
        end
        612: begin
            cosine_reg0 <= 36'sb11111000111110110100101000001001000;
            sine_reg0   <= 36'sb111011100010000110101010111011011;
        end
        613: begin
            cosine_reg0 <= 36'sb11111000111101010111000010011100100;
            sine_reg0   <= 36'sb111011101000001101110000001001000;
        end
        614: begin
            cosine_reg0 <= 36'sb11111000111011111001010011001001100;
            sine_reg0   <= 36'sb111011101110010100110011000011011;
        end
        615: begin
            cosine_reg0 <= 36'sb11111000111010011011011010010000011;
            sine_reg0   <= 36'sb111011110100011011110011101010100;
        end
        616: begin
            cosine_reg0 <= 36'sb11111000111000111101010111110001001;
            sine_reg0   <= 36'sb111011111010100010110001111110000;
        end
        617: begin
            cosine_reg0 <= 36'sb11111000110111011111001011101011110;
            sine_reg0   <= 36'sb111100000000101001101101111101101;
        end
        618: begin
            cosine_reg0 <= 36'sb11111000110110000000110110000000010;
            sine_reg0   <= 36'sb111100000110110000100111101001010;
        end
        619: begin
            cosine_reg0 <= 36'sb11111000110100100010010110101110111;
            sine_reg0   <= 36'sb111100001100110111011111000000100;
        end
        620: begin
            cosine_reg0 <= 36'sb11111000110011000011101101110111100;
            sine_reg0   <= 36'sb111100010010111110010100000011010;
        end
        621: begin
            cosine_reg0 <= 36'sb11111000110001100100111011011010001;
            sine_reg0   <= 36'sb111100011001000101000110110001010;
        end
        622: begin
            cosine_reg0 <= 36'sb11111000110000000101111111010111000;
            sine_reg0   <= 36'sb111100011111001011110111001010001;
        end
        623: begin
            cosine_reg0 <= 36'sb11111000101110100110111001101110001;
            sine_reg0   <= 36'sb111100100101010010100101001101111;
        end
        624: begin
            cosine_reg0 <= 36'sb11111000101101000111101010011111101;
            sine_reg0   <= 36'sb111100101011011001010000111100001;
        end
        625: begin
            cosine_reg0 <= 36'sb11111000101011101000010001101011011;
            sine_reg0   <= 36'sb111100110001011111111010010100101;
        end
        626: begin
            cosine_reg0 <= 36'sb11111000101010001000101111010001100;
            sine_reg0   <= 36'sb111100110111100110100001010111001;
        end
        627: begin
            cosine_reg0 <= 36'sb11111000101000101001000011010010001;
            sine_reg0   <= 36'sb111100111101101101000110000011100;
        end
        628: begin
            cosine_reg0 <= 36'sb11111000100111001001001101101101010;
            sine_reg0   <= 36'sb111101000011110011101000011001100;
        end
        629: begin
            cosine_reg0 <= 36'sb11111000100101101001001110100011000;
            sine_reg0   <= 36'sb111101001001111010001000011000110;
        end
        630: begin
            cosine_reg0 <= 36'sb11111000100100001001000101110011011;
            sine_reg0   <= 36'sb111101010000000000100110000001001;
        end
        631: begin
            cosine_reg0 <= 36'sb11111000100010101000110011011110011;
            sine_reg0   <= 36'sb111101010110000111000001010010011;
        end
        632: begin
            cosine_reg0 <= 36'sb11111000100001001000010111100100001;
            sine_reg0   <= 36'sb111101011100001101011010001100011;
        end
        633: begin
            cosine_reg0 <= 36'sb11111000011111100111110010000100110;
            sine_reg0   <= 36'sb111101100010010011110000101110101;
        end
        634: begin
            cosine_reg0 <= 36'sb11111000011110000111000011000000010;
            sine_reg0   <= 36'sb111101101000011010000100111001001;
        end
        635: begin
            cosine_reg0 <= 36'sb11111000011100100110001010010110101;
            sine_reg0   <= 36'sb111101101110100000010110101011100;
        end
        636: begin
            cosine_reg0 <= 36'sb11111000011011000101001000001000000;
            sine_reg0   <= 36'sb111101110100100110100110000101101;
        end
        637: begin
            cosine_reg0 <= 36'sb11111000011001100011111100010100011;
            sine_reg0   <= 36'sb111101111010101100110011000111001;
        end
        638: begin
            cosine_reg0 <= 36'sb11111000011000000010100110111011111;
            sine_reg0   <= 36'sb111110000000110010111101101111111;
        end
        639: begin
            cosine_reg0 <= 36'sb11111000010110100001000111111110101;
            sine_reg0   <= 36'sb111110000110111001000101111111110;
        end
        640: begin
            cosine_reg0 <= 36'sb11111000010100111111011111011100100;
            sine_reg0   <= 36'sb111110001100111111001011110110010;
        end
        641: begin
            cosine_reg0 <= 36'sb11111000010011011101101101010101101;
            sine_reg0   <= 36'sb111110010011000101001111010011010;
        end
        642: begin
            cosine_reg0 <= 36'sb11111000010001111011110001101010001;
            sine_reg0   <= 36'sb111110011001001011010000010110101;
        end
        643: begin
            cosine_reg0 <= 36'sb11111000010000011001101100011010000;
            sine_reg0   <= 36'sb111110011111010001001111000000000;
        end
        644: begin
            cosine_reg0 <= 36'sb11111000001110110111011101100101011;
            sine_reg0   <= 36'sb111110100101010111001011001111010;
        end
        645: begin
            cosine_reg0 <= 36'sb11111000001101010101000101001100001;
            sine_reg0   <= 36'sb111110101011011101000101000100000;
        end
        646: begin
            cosine_reg0 <= 36'sb11111000001011110010100011001110101;
            sine_reg0   <= 36'sb111110110001100010111100011110001;
        end
        647: begin
            cosine_reg0 <= 36'sb11111000001010001111110111101100101;
            sine_reg0   <= 36'sb111110110111101000110001011101011;
        end
        648: begin
            cosine_reg0 <= 36'sb11111000001000101101000010100110011;
            sine_reg0   <= 36'sb111110111101101110100100000001100;
        end
        649: begin
            cosine_reg0 <= 36'sb11111000000111001010000011111011111;
            sine_reg0   <= 36'sb111111000011110100010100001010010;
        end
        650: begin
            cosine_reg0 <= 36'sb11111000000101100110111011101101001;
            sine_reg0   <= 36'sb111111001001111010000001110111011;
        end
        651: begin
            cosine_reg0 <= 36'sb11111000000100000011101001111010010;
            sine_reg0   <= 36'sb111111001111111111101101001000110;
        end
        652: begin
            cosine_reg0 <= 36'sb11111000000010100000001110100011011;
            sine_reg0   <= 36'sb111111010110000101010101111110000;
        end
        653: begin
            cosine_reg0 <= 36'sb11111000000000111100101001101000100;
            sine_reg0   <= 36'sb111111011100001010111100010110111;
        end
        654: begin
            cosine_reg0 <= 36'sb11110111111111011000111011001001101;
            sine_reg0   <= 36'sb111111100010010000100000010011011;
        end
        655: begin
            cosine_reg0 <= 36'sb11110111111101110101000011000110111;
            sine_reg0   <= 36'sb111111101000010110000001110011000;
        end
        656: begin
            cosine_reg0 <= 36'sb11110111111100010001000001100000010;
            sine_reg0   <= 36'sb111111101110011011100000110101110;
        end
        657: begin
            cosine_reg0 <= 36'sb11110111111010101100110110010101111;
            sine_reg0   <= 36'sb111111110100100000111101011011001;
        end
        658: begin
            cosine_reg0 <= 36'sb11110111111001001000100001100111110;
            sine_reg0   <= 36'sb111111111010100110010111100011001;
        end
        659: begin
            cosine_reg0 <= 36'sb11110111110111100100000011010110001;
            sine_reg0   <= 36'sb1000000000000101011101111001101011;
        end
        660: begin
            cosine_reg0 <= 36'sb11110111110101111111011011100000110;
            sine_reg0   <= 36'sb1000000000110110001000100011001110;
        end
        661: begin
            cosine_reg0 <= 36'sb11110111110100011010101010000111111;
            sine_reg0   <= 36'sb1000000001100110110010111000111111;
        end
        662: begin
            cosine_reg0 <= 36'sb11110111110010110101101111001011101;
            sine_reg0   <= 36'sb1000000010010111011100111010111101;
        end
        663: begin
            cosine_reg0 <= 36'sb11110111110001010000101010101011111;
            sine_reg0   <= 36'sb1000000011001000000110101001000101;
        end
        664: begin
            cosine_reg0 <= 36'sb11110111101111101011011100101000110;
            sine_reg0   <= 36'sb1000000011111000110000000011010111;
        end
        665: begin
            cosine_reg0 <= 36'sb11110111101110000110000101000010011;
            sine_reg0   <= 36'sb1000000100101001011001001001110000;
        end
        666: begin
            cosine_reg0 <= 36'sb11110111101100100000100011111000111;
            sine_reg0   <= 36'sb1000000101011010000001111100001110;
        end
        667: begin
            cosine_reg0 <= 36'sb11110111101010111010111001001100001;
            sine_reg0   <= 36'sb1000000110001010101010011010101111;
        end
        668: begin
            cosine_reg0 <= 36'sb11110111101001010101000100111100010;
            sine_reg0   <= 36'sb1000000110111011010010100101010010;
        end
        669: begin
            cosine_reg0 <= 36'sb11110111100111101111000111001001011;
            sine_reg0   <= 36'sb1000000111101011111010011011110101;
        end
        670: begin
            cosine_reg0 <= 36'sb11110111100110001000111111110011100;
            sine_reg0   <= 36'sb1000001000011100100001111110010101;
        end
        671: begin
            cosine_reg0 <= 36'sb11110111100100100010101110111010101;
            sine_reg0   <= 36'sb1000001001001101001001001100110001;
        end
        672: begin
            cosine_reg0 <= 36'sb11110111100010111100010100011111000;
            sine_reg0   <= 36'sb1000001001111101110000000111000111;
        end
        673: begin
            cosine_reg0 <= 36'sb11110111100001010101110000100000101;
            sine_reg0   <= 36'sb1000001010101110010110101101010101;
        end
        674: begin
            cosine_reg0 <= 36'sb11110111011111101111000010111111011;
            sine_reg0   <= 36'sb1000001011011110111100111111011001;
        end
        675: begin
            cosine_reg0 <= 36'sb11110111011110001000001011111011100;
            sine_reg0   <= 36'sb1000001100001111100010111101010010;
        end
        676: begin
            cosine_reg0 <= 36'sb11110111011100100001001011010101001;
            sine_reg0   <= 36'sb1000001101000000001000100110111101;
        end
        677: begin
            cosine_reg0 <= 36'sb11110111011010111010000001001100001;
            sine_reg0   <= 36'sb1000001101110000101101111100011001;
        end
        678: begin
            cosine_reg0 <= 36'sb11110111011001010010101101100000101;
            sine_reg0   <= 36'sb1000001110100001010010111101100011;
        end
        679: begin
            cosine_reg0 <= 36'sb11110111010111101011010000010010101;
            sine_reg0   <= 36'sb1000001111010001110111101010011011;
        end
        680: begin
            cosine_reg0 <= 36'sb11110111010110000011101001100010011;
            sine_reg0   <= 36'sb1000010000000010011100000010111101;
        end
        681: begin
            cosine_reg0 <= 36'sb11110111010100011011111001001111111;
            sine_reg0   <= 36'sb1000010000110011000000000111001001;
        end
        682: begin
            cosine_reg0 <= 36'sb11110111010010110011111111011011000;
            sine_reg0   <= 36'sb1000010001100011100011110110111011;
        end
        683: begin
            cosine_reg0 <= 36'sb11110111010001001011111100000100000;
            sine_reg0   <= 36'sb1000010010010100000111010010010100;
        end
        684: begin
            cosine_reg0 <= 36'sb11110111001111100011101111001010111;
            sine_reg0   <= 36'sb1000010011000100101010011001001111;
        end
        685: begin
            cosine_reg0 <= 36'sb11110111001101111011011000101111110;
            sine_reg0   <= 36'sb1000010011110101001101001011101100;
        end
        686: begin
            cosine_reg0 <= 36'sb11110111001100010010111000110010101;
            sine_reg0   <= 36'sb1000010100100101101111101001101001;
        end
        687: begin
            cosine_reg0 <= 36'sb11110111001010101010001111010011101;
            sine_reg0   <= 36'sb1000010101010110010001110011000100;
        end
        688: begin
            cosine_reg0 <= 36'sb11110111001001000001011100010010110;
            sine_reg0   <= 36'sb1000010110000110110011100111111011;
        end
        689: begin
            cosine_reg0 <= 36'sb11110111000111011000011111110000000;
            sine_reg0   <= 36'sb1000010110110111010101001000001100;
        end
        690: begin
            cosine_reg0 <= 36'sb11110111000101101111011001101011101;
            sine_reg0   <= 36'sb1000010111100111110110010011110110;
        end
        691: begin
            cosine_reg0 <= 36'sb11110111000100000110001010000101100;
            sine_reg0   <= 36'sb1000011000011000010111001010110101;
        end
        692: begin
            cosine_reg0 <= 36'sb11110111000010011100110000111101110;
            sine_reg0   <= 36'sb1000011001001000110111101101001010;
        end
        693: begin
            cosine_reg0 <= 36'sb11110111000000110011001110010100100;
            sine_reg0   <= 36'sb1000011001111001010111111010110001;
        end
        694: begin
            cosine_reg0 <= 36'sb11110110111111001001100010001001110;
            sine_reg0   <= 36'sb1000011010101001110111110011101000;
        end
        695: begin
            cosine_reg0 <= 36'sb11110110111101011111101100011101101;
            sine_reg0   <= 36'sb1000011011011010010111010111101111;
        end
        696: begin
            cosine_reg0 <= 36'sb11110110111011110101101101010000001;
            sine_reg0   <= 36'sb1000011100001010110110100111000011;
        end
        697: begin
            cosine_reg0 <= 36'sb11110110111010001011100100100001011;
            sine_reg0   <= 36'sb1000011100111011010101100001100010;
        end
        698: begin
            cosine_reg0 <= 36'sb11110110111000100001010010010001011;
            sine_reg0   <= 36'sb1000011101101011110100000111001010;
        end
        699: begin
            cosine_reg0 <= 36'sb11110110110110110110110110100000001;
            sine_reg0   <= 36'sb1000011110011100010010010111111001;
        end
        700: begin
            cosine_reg0 <= 36'sb11110110110101001100010001001101111;
            sine_reg0   <= 36'sb1000011111001100110000010011101111;
        end
        701: begin
            cosine_reg0 <= 36'sb11110110110011100001100010011010101;
            sine_reg0   <= 36'sb1000011111111101001101111010101000;
        end
        702: begin
            cosine_reg0 <= 36'sb11110110110001110110101010000110011;
            sine_reg0   <= 36'sb1000100000101101101011001100100010;
        end
        703: begin
            cosine_reg0 <= 36'sb11110110110000001011101000010001001;
            sine_reg0   <= 36'sb1000100001011110001000001001011101;
        end
        704: begin
            cosine_reg0 <= 36'sb11110110101110100000011100111011001;
            sine_reg0   <= 36'sb1000100010001110100100110001010110;
        end
        705: begin
            cosine_reg0 <= 36'sb11110110101100110101001000000100011;
            sine_reg0   <= 36'sb1000100010111111000001000100001011;
        end
        706: begin
            cosine_reg0 <= 36'sb11110110101011001001101001101100111;
            sine_reg0   <= 36'sb1000100011101111011101000001111011;
        end
        707: begin
            cosine_reg0 <= 36'sb11110110101001011110000001110100110;
            sine_reg0   <= 36'sb1000100100011111111000101010100011;
        end
        708: begin
            cosine_reg0 <= 36'sb11110110100111110010010000011100000;
            sine_reg0   <= 36'sb1000100101010000010011111110000001;
        end
        709: begin
            cosine_reg0 <= 36'sb11110110100110000110010101100010110;
            sine_reg0   <= 36'sb1000100110000000101110111100010100;
        end
        710: begin
            cosine_reg0 <= 36'sb11110110100100011010010001001001001;
            sine_reg0   <= 36'sb1000100110110001001001100101011011;
        end
        711: begin
            cosine_reg0 <= 36'sb11110110100010101110000011001111000;
            sine_reg0   <= 36'sb1000100111100001100011111001010010;
        end
        712: begin
            cosine_reg0 <= 36'sb11110110100001000001101011110100101;
            sine_reg0   <= 36'sb1000101000010001111101110111111001;
        end
        713: begin
            cosine_reg0 <= 36'sb11110110011111010101001010111010000;
            sine_reg0   <= 36'sb1000101001000010010111100001001100;
        end
        714: begin
            cosine_reg0 <= 36'sb11110110011101101000100000011111010;
            sine_reg0   <= 36'sb1000101001110010110000110101001100;
        end
        715: begin
            cosine_reg0 <= 36'sb11110110011011111011101100100100010;
            sine_reg0   <= 36'sb1000101010100011001001110011110100;
        end
        716: begin
            cosine_reg0 <= 36'sb11110110011010001110101111001001010;
            sine_reg0   <= 36'sb1000101011010011100010011101000101;
        end
        717: begin
            cosine_reg0 <= 36'sb11110110011000100001101000001110010;
            sine_reg0   <= 36'sb1000101100000011111010110000111011;
        end
        718: begin
            cosine_reg0 <= 36'sb11110110010110110100010111110011011;
            sine_reg0   <= 36'sb1000101100110100010010101111010101;
        end
        719: begin
            cosine_reg0 <= 36'sb11110110010101000110111101111000101;
            sine_reg0   <= 36'sb1000101101100100101010011000010010;
        end
        720: begin
            cosine_reg0 <= 36'sb11110110010011011001011010011110000;
            sine_reg0   <= 36'sb1000101110010101000001101011101111;
        end
        721: begin
            cosine_reg0 <= 36'sb11110110010001101011101101100011110;
            sine_reg0   <= 36'sb1000101111000101011000101001101010;
        end
        722: begin
            cosine_reg0 <= 36'sb11110110001111111101110111001001110;
            sine_reg0   <= 36'sb1000101111110101101111010010000001;
        end
        723: begin
            cosine_reg0 <= 36'sb11110110001110001111110111010000001;
            sine_reg0   <= 36'sb1000110000100110000101100100110011;
        end
        724: begin
            cosine_reg0 <= 36'sb11110110001100100001101101110111001;
            sine_reg0   <= 36'sb1000110001010110011011100001111110;
        end
        725: begin
            cosine_reg0 <= 36'sb11110110001010110011011010111110100;
            sine_reg0   <= 36'sb1000110010000110110001001001100000;
        end
        726: begin
            cosine_reg0 <= 36'sb11110110001001000100111110100110100;
            sine_reg0   <= 36'sb1000110010110111000110011011010111;
        end
        727: begin
            cosine_reg0 <= 36'sb11110110000111010110011000101111010;
            sine_reg0   <= 36'sb1000110011100111011011010111100001;
        end
        728: begin
            cosine_reg0 <= 36'sb11110110000101100111101001011000110;
            sine_reg0   <= 36'sb1000110100010111101111111101111101;
        end
        729: begin
            cosine_reg0 <= 36'sb11110110000011111000110000100011000;
            sine_reg0   <= 36'sb1000110101001000000100001110101000;
        end
        730: begin
            cosine_reg0 <= 36'sb11110110000010001001101110001110001;
            sine_reg0   <= 36'sb1000110101111000011000001001100000;
        end
        731: begin
            cosine_reg0 <= 36'sb11110110000000011010100010011010001;
            sine_reg0   <= 36'sb1000110110101000101011101110100101;
        end
        732: begin
            cosine_reg0 <= 36'sb11110101111110101011001101000111010;
            sine_reg0   <= 36'sb1000110111011000111110111101110011;
        end
        733: begin
            cosine_reg0 <= 36'sb11110101111100111011101110010101011;
            sine_reg0   <= 36'sb1000111000001001010001110111001001;
        end
        734: begin
            cosine_reg0 <= 36'sb11110101111011001100000110000100101;
            sine_reg0   <= 36'sb1000111000111001100100011010100110;
        end
        735: begin
            cosine_reg0 <= 36'sb11110101111001011100010100010101001;
            sine_reg0   <= 36'sb1000111001101001110110101000000110;
        end
        736: begin
            cosine_reg0 <= 36'sb11110101110111101100011001000110111;
            sine_reg0   <= 36'sb1000111010011010001000011111101001;
        end
        737: begin
            cosine_reg0 <= 36'sb11110101110101111100010100011010000;
            sine_reg0   <= 36'sb1000111011001010011010000001001101;
        end
        738: begin
            cosine_reg0 <= 36'sb11110101110100001100000110001110011;
            sine_reg0   <= 36'sb1000111011111010101011001100101111;
        end
        739: begin
            cosine_reg0 <= 36'sb11110101110010011011101110100100011;
            sine_reg0   <= 36'sb1000111100101010111100000010001111;
        end
        740: begin
            cosine_reg0 <= 36'sb11110101110000101011001101011011111;
            sine_reg0   <= 36'sb1000111101011011001100100001101001;
        end
        741: begin
            cosine_reg0 <= 36'sb11110101101110111010100010110101000;
            sine_reg0   <= 36'sb1000111110001011011100101010111100;
        end
        742: begin
            cosine_reg0 <= 36'sb11110101101101001001101110101111111;
            sine_reg0   <= 36'sb1000111110111011101100011110000111;
        end
        743: begin
            cosine_reg0 <= 36'sb11110101101011011000110001001100011;
            sine_reg0   <= 36'sb1000111111101011111011111011000111;
        end
        744: begin
            cosine_reg0 <= 36'sb11110101101001100111101010001010110;
            sine_reg0   <= 36'sb1001000000011100001011000001111011;
        end
        745: begin
            cosine_reg0 <= 36'sb11110101100111110110011001101011000;
            sine_reg0   <= 36'sb1001000001001100011001110010100000;
        end
        746: begin
            cosine_reg0 <= 36'sb11110101100110000100111111101101001;
            sine_reg0   <= 36'sb1001000001111100101000001100110101;
        end
        747: begin
            cosine_reg0 <= 36'sb11110101100100010011011100010001011;
            sine_reg0   <= 36'sb1001000010101100110110010000111000;
        end
        748: begin
            cosine_reg0 <= 36'sb11110101100010100001101111010111101;
            sine_reg0   <= 36'sb1001000011011101000011111110100111;
        end
        749: begin
            cosine_reg0 <= 36'sb11110101100000101111111001000000001;
            sine_reg0   <= 36'sb1001000100001101010001010110000001;
        end
        750: begin
            cosine_reg0 <= 36'sb11110101011110111101111001001010111;
            sine_reg0   <= 36'sb1001000100111101011110010111000011;
        end
        751: begin
            cosine_reg0 <= 36'sb11110101011101001011101111110111110;
            sine_reg0   <= 36'sb1001000101101101101011000001101011;
        end
        752: begin
            cosine_reg0 <= 36'sb11110101011011011001011101000111001;
            sine_reg0   <= 36'sb1001000110011101110111010101111000;
        end
        753: begin
            cosine_reg0 <= 36'sb11110101011001100111000000111000111;
            sine_reg0   <= 36'sb1001000111001110000011010011101000;
        end
        754: begin
            cosine_reg0 <= 36'sb11110101010111110100011011001101001;
            sine_reg0   <= 36'sb1001000111111110001110111010111001;
        end
        755: begin
            cosine_reg0 <= 36'sb11110101010110000001101100000100000;
            sine_reg0   <= 36'sb1001001000101110011010001011101001;
        end
        756: begin
            cosine_reg0 <= 36'sb11110101010100001110110011011101100;
            sine_reg0   <= 36'sb1001001001011110100101000101110110;
        end
        757: begin
            cosine_reg0 <= 36'sb11110101010010011011110001011001101;
            sine_reg0   <= 36'sb1001001010001110101111101001011111;
        end
        758: begin
            cosine_reg0 <= 36'sb11110101010000101000100101111000101;
            sine_reg0   <= 36'sb1001001010111110111001110110100001;
        end
        759: begin
            cosine_reg0 <= 36'sb11110101001110110101010000111010011;
            sine_reg0   <= 36'sb1001001011101111000011101100111011;
        end
        760: begin
            cosine_reg0 <= 36'sb11110101001101000001110010011111001;
            sine_reg0   <= 36'sb1001001100011111001101001100101010;
        end
        761: begin
            cosine_reg0 <= 36'sb11110101001011001110001010100110110;
            sine_reg0   <= 36'sb1001001101001111010110010101101110;
        end
        762: begin
            cosine_reg0 <= 36'sb11110101001001011010011001010001100;
            sine_reg0   <= 36'sb1001001101111111011111001000000100;
        end
        763: begin
            cosine_reg0 <= 36'sb11110101000111100110011110011111011;
            sine_reg0   <= 36'sb1001001110101111100111100011101010;
        end
        764: begin
            cosine_reg0 <= 36'sb11110101000101110010011010010000100;
            sine_reg0   <= 36'sb1001001111011111101111101000011110;
        end
        765: begin
            cosine_reg0 <= 36'sb11110101000011111110001100100100110;
            sine_reg0   <= 36'sb1001010000001111110111010110011111;
        end
        766: begin
            cosine_reg0 <= 36'sb11110101000010001001110101011100100;
            sine_reg0   <= 36'sb1001010000111111111110101101101011;
        end
        767: begin
            cosine_reg0 <= 36'sb11110101000000010101010100110111100;
            sine_reg0   <= 36'sb1001010001110000000101101101111111;
        end
        768: begin
            cosine_reg0 <= 36'sb11110100111110100000101010110110001;
            sine_reg0   <= 36'sb1001010010100000001100010111011010;
        end
        769: begin
            cosine_reg0 <= 36'sb11110100111100101011110111011000001;
            sine_reg0   <= 36'sb1001010011010000010010101001111011;
        end
        770: begin
            cosine_reg0 <= 36'sb11110100111010110110111010011101111;
            sine_reg0   <= 36'sb1001010100000000011000100101011111;
        end
        771: begin
            cosine_reg0 <= 36'sb11110100111001000001110100000111010;
            sine_reg0   <= 36'sb1001010100110000011110001010000100;
        end
        772: begin
            cosine_reg0 <= 36'sb11110100110111001100100100010100011;
            sine_reg0   <= 36'sb1001010101100000100011010111101001;
        end
        773: begin
            cosine_reg0 <= 36'sb11110100110101010111001011000101011;
            sine_reg0   <= 36'sb1001010110010000101000001110001011;
        end
        774: begin
            cosine_reg0 <= 36'sb11110100110011100001101000011010010;
            sine_reg0   <= 36'sb1001010111000000101100101101101010;
        end
        775: begin
            cosine_reg0 <= 36'sb11110100110001101011111100010011000;
            sine_reg0   <= 36'sb1001010111110000110000110110000010;
        end
        776: begin
            cosine_reg0 <= 36'sb11110100101111110110000110101111111;
            sine_reg0   <= 36'sb1001011000100000110100100111010010;
        end
        777: begin
            cosine_reg0 <= 36'sb11110100101110000000000111110000111;
            sine_reg0   <= 36'sb1001011001010000111000000001011001;
        end
        778: begin
            cosine_reg0 <= 36'sb11110100101100001001111111010110001;
            sine_reg0   <= 36'sb1001011010000000111011000100010100;
        end
        779: begin
            cosine_reg0 <= 36'sb11110100101010010011101101011111100;
            sine_reg0   <= 36'sb1001011010110000111101110000000010;
        end
        780: begin
            cosine_reg0 <= 36'sb11110100101000011101010010001101010;
            sine_reg0   <= 36'sb1001011011100001000000000100100001;
        end
        781: begin
            cosine_reg0 <= 36'sb11110100100110100110101101011111011;
            sine_reg0   <= 36'sb1001011100010001000010000001101110;
        end
        782: begin
            cosine_reg0 <= 36'sb11110100100100101111111111010110000;
            sine_reg0   <= 36'sb1001011101000001000011100111101001;
        end
        783: begin
            cosine_reg0 <= 36'sb11110100100010111001000111110001001;
            sine_reg0   <= 36'sb1001011101110001000100110110001110;
        end
        784: begin
            cosine_reg0 <= 36'sb11110100100001000010000110110000111;
            sine_reg0   <= 36'sb1001011110100001000101101101011101;
        end
        785: begin
            cosine_reg0 <= 36'sb11110100011111001010111100010101010;
            sine_reg0   <= 36'sb1001011111010001000110001101010100;
        end
        786: begin
            cosine_reg0 <= 36'sb11110100011101010011101000011110011;
            sine_reg0   <= 36'sb1001100000000001000110010101110000;
        end
        787: begin
            cosine_reg0 <= 36'sb11110100011011011100001011001100011;
            sine_reg0   <= 36'sb1001100000110001000110000110110000;
        end
        788: begin
            cosine_reg0 <= 36'sb11110100011001100100100100011111010;
            sine_reg0   <= 36'sb1001100001100001000101100000010001;
        end
        789: begin
            cosine_reg0 <= 36'sb11110100010111101100110100010111001;
            sine_reg0   <= 36'sb1001100010010001000100100010010011;
        end
        790: begin
            cosine_reg0 <= 36'sb11110100010101110100111010110100001;
            sine_reg0   <= 36'sb1001100011000001000011001100110011;
        end
        791: begin
            cosine_reg0 <= 36'sb11110100010011111100110111110110001;
            sine_reg0   <= 36'sb1001100011110001000001011111110000;
        end
        792: begin
            cosine_reg0 <= 36'sb11110100010010000100101011011101010;
            sine_reg0   <= 36'sb1001100100100000111111011011000111;
        end
        793: begin
            cosine_reg0 <= 36'sb11110100010000001100010101101001110;
            sine_reg0   <= 36'sb1001100101010000111100111110110110;
        end
        794: begin
            cosine_reg0 <= 36'sb11110100001110010011110110011011100;
            sine_reg0   <= 36'sb1001100110000000111010001010111101;
        end
        795: begin
            cosine_reg0 <= 36'sb11110100001100011011001101110010110;
            sine_reg0   <= 36'sb1001100110110000110110111111011000;
        end
        796: begin
            cosine_reg0 <= 36'sb11110100001010100010011011101111011;
            sine_reg0   <= 36'sb1001100111100000110011011100000111;
        end
        797: begin
            cosine_reg0 <= 36'sb11110100001000101001100000010001101;
            sine_reg0   <= 36'sb1001101000010000101111100001000111;
        end
        798: begin
            cosine_reg0 <= 36'sb11110100000110110000011011011001100;
            sine_reg0   <= 36'sb1001101001000000101011001110010110;
        end
        799: begin
            cosine_reg0 <= 36'sb11110100000100110111001101000111000;
            sine_reg0   <= 36'sb1001101001110000100110100011110011;
        end
        800: begin
            cosine_reg0 <= 36'sb11110100000010111101110101011010010;
            sine_reg0   <= 36'sb1001101010100000100001100001011100;
        end
        801: begin
            cosine_reg0 <= 36'sb11110100000001000100010100010011011;
            sine_reg0   <= 36'sb1001101011010000011100000111001110;
        end
        802: begin
            cosine_reg0 <= 36'sb11110011111111001010101001110010100;
            sine_reg0   <= 36'sb1001101100000000010110010101001001;
        end
        803: begin
            cosine_reg0 <= 36'sb11110011111101010000110101110111100;
            sine_reg0   <= 36'sb1001101100110000010000001011001010;
        end
        804: begin
            cosine_reg0 <= 36'sb11110011111011010110111000100010101;
            sine_reg0   <= 36'sb1001101101100000001001101001001111;
        end
        805: begin
            cosine_reg0 <= 36'sb11110011111001011100110001110011111;
            sine_reg0   <= 36'sb1001101110010000000010101111010111;
        end
        806: begin
            cosine_reg0 <= 36'sb11110011110111100010100001101011010;
            sine_reg0   <= 36'sb1001101110111111111011011101011111;
        end
        807: begin
            cosine_reg0 <= 36'sb11110011110101101000001000001001000;
            sine_reg0   <= 36'sb1001101111101111110011110011100110;
        end
        808: begin
            cosine_reg0 <= 36'sb11110011110011101101100101001101000;
            sine_reg0   <= 36'sb1001110000011111101011110001101010;
        end
        809: begin
            cosine_reg0 <= 36'sb11110011110001110010111000110111100;
            sine_reg0   <= 36'sb1001110001001111100011010111101001;
        end
        810: begin
            cosine_reg0 <= 36'sb11110011101111111000000011001000100;
            sine_reg0   <= 36'sb1001110001111111011010100101100010;
        end
        811: begin
            cosine_reg0 <= 36'sb11110011101101111101000100000000001;
            sine_reg0   <= 36'sb1001110010101111010001011011010010;
        end
        812: begin
            cosine_reg0 <= 36'sb11110011101100000001111011011110011;
            sine_reg0   <= 36'sb1001110011011111000111111000110111;
        end
        813: begin
            cosine_reg0 <= 36'sb11110011101010000110101001100011010;
            sine_reg0   <= 36'sb1001110100001110111101111110010000;
        end
        814: begin
            cosine_reg0 <= 36'sb11110011101000001011001110001111000;
            sine_reg0   <= 36'sb1001110100111110110011101011011100;
        end
        815: begin
            cosine_reg0 <= 36'sb11110011100110001111101001100001101;
            sine_reg0   <= 36'sb1001110101101110101001000000010111;
        end
        816: begin
            cosine_reg0 <= 36'sb11110011100100010011111011011011010;
            sine_reg0   <= 36'sb1001110110011110011101111101000000;
        end
        817: begin
            cosine_reg0 <= 36'sb11110011100010011000000011111011110;
            sine_reg0   <= 36'sb1001110111001110010010100001010110;
        end
        818: begin
            cosine_reg0 <= 36'sb11110011100000011100000011000011100;
            sine_reg0   <= 36'sb1001110111111110000110101101010110;
        end
        819: begin
            cosine_reg0 <= 36'sb11110011011110011111111000110010011;
            sine_reg0   <= 36'sb1001111000101101111010100000111111;
        end
        820: begin
            cosine_reg0 <= 36'sb11110011011100100011100101001000100;
            sine_reg0   <= 36'sb1001111001011101101101111100001111;
        end
        821: begin
            cosine_reg0 <= 36'sb11110011011010100111001000000101111;
            sine_reg0   <= 36'sb1001111010001101100000111111000100;
        end
        822: begin
            cosine_reg0 <= 36'sb11110011011000101010100001101010101;
            sine_reg0   <= 36'sb1001111010111101010011101001011100;
        end
        823: begin
            cosine_reg0 <= 36'sb11110011010110101101110001110111000;
            sine_reg0   <= 36'sb1001111011101101000101111011010101;
        end
        824: begin
            cosine_reg0 <= 36'sb11110011010100110000111000101010110;
            sine_reg0   <= 36'sb1001111100011100110111110100101110;
        end
        825: begin
            cosine_reg0 <= 36'sb11110011010010110011110110000110010;
            sine_reg0   <= 36'sb1001111101001100101001010101100100;
        end
        826: begin
            cosine_reg0 <= 36'sb11110011010000110110101010001001011;
            sine_reg0   <= 36'sb1001111101111100011010011101110110;
        end
        827: begin
            cosine_reg0 <= 36'sb11110011001110111001010100110100011;
            sine_reg0   <= 36'sb1001111110101100001011001101100010;
        end
        828: begin
            cosine_reg0 <= 36'sb11110011001100111011110110000111001;
            sine_reg0   <= 36'sb1001111111011011111011100100100110;
        end
        829: begin
            cosine_reg0 <= 36'sb11110011001010111110001110000001110;
            sine_reg0   <= 36'sb1010000000001011101011100011000000;
        end
        830: begin
            cosine_reg0 <= 36'sb11110011001001000000011100100100100;
            sine_reg0   <= 36'sb1010000000111011011011001000101111;
        end
        831: begin
            cosine_reg0 <= 36'sb11110011000111000010100001101111010;
            sine_reg0   <= 36'sb1010000001101011001010010101110001;
        end
        832: begin
            cosine_reg0 <= 36'sb11110011000101000100011101100010001;
            sine_reg0   <= 36'sb1010000010011010111001001010000011;
        end
        833: begin
            cosine_reg0 <= 36'sb11110011000011000110001111111101010;
            sine_reg0   <= 36'sb1010000011001010100111100101100100;
        end
        834: begin
            cosine_reg0 <= 36'sb11110011000001000111111001000000110;
            sine_reg0   <= 36'sb1010000011111010010101101000010010;
        end
        835: begin
            cosine_reg0 <= 36'sb11110010111111001001011000101100101;
            sine_reg0   <= 36'sb1010000100101010000011010010001011;
        end
        836: begin
            cosine_reg0 <= 36'sb11110010111101001010101111000000111;
            sine_reg0   <= 36'sb1010000101011001110000100011001101;
        end
        837: begin
            cosine_reg0 <= 36'sb11110010111011001011111011111101101;
            sine_reg0   <= 36'sb1010000110001001011101011011011000;
        end
        838: begin
            cosine_reg0 <= 36'sb11110010111001001100111111100011001;
            sine_reg0   <= 36'sb1010000110111001001001111010100111;
        end
        839: begin
            cosine_reg0 <= 36'sb11110010110111001101111001110001001;
            sine_reg0   <= 36'sb1010000111101000110110000000111011;
        end
        840: begin
            cosine_reg0 <= 36'sb11110010110101001110101010101000000;
            sine_reg0   <= 36'sb1010001000011000100001101110010001;
        end
        841: begin
            cosine_reg0 <= 36'sb11110010110011001111010010000111110;
            sine_reg0   <= 36'sb1010001001001000001101000010100111;
        end
        842: begin
            cosine_reg0 <= 36'sb11110010110001001111110000010000011;
            sine_reg0   <= 36'sb1010001001110111110111111101111011;
        end
        843: begin
            cosine_reg0 <= 36'sb11110010101111010000000101000001111;
            sine_reg0   <= 36'sb1010001010100111100010100000001100;
        end
        844: begin
            cosine_reg0 <= 36'sb11110010101101010000010000011100101;
            sine_reg0   <= 36'sb1010001011010111001100101001010111;
        end
        845: begin
            cosine_reg0 <= 36'sb11110010101011010000010010100000011;
            sine_reg0   <= 36'sb1010001100000110110110011001011011;
        end
        846: begin
            cosine_reg0 <= 36'sb11110010101001010000001011001101011;
            sine_reg0   <= 36'sb1010001100110110011111110000010111;
        end
        847: begin
            cosine_reg0 <= 36'sb11110010100111001111111010100011110;
            sine_reg0   <= 36'sb1010001101100110001000101110000111;
        end
        848: begin
            cosine_reg0 <= 36'sb11110010100101001111100000100011100;
            sine_reg0   <= 36'sb1010001110010101110001010010101011;
        end
        849: begin
            cosine_reg0 <= 36'sb11110010100011001110111101001100101;
            sine_reg0   <= 36'sb1010001111000101011001011110000000;
        end
        850: begin
            cosine_reg0 <= 36'sb11110010100001001110010000011111010;
            sine_reg0   <= 36'sb1010001111110101000001010000000101;
        end
        851: begin
            cosine_reg0 <= 36'sb11110010011111001101011010011011101;
            sine_reg0   <= 36'sb1010010000100100101000101000110111;
        end
        852: begin
            cosine_reg0 <= 36'sb11110010011101001100011011000001101;
            sine_reg0   <= 36'sb1010010001010100001111101000010110;
        end
        853: begin
            cosine_reg0 <= 36'sb11110010011011001011010010010001011;
            sine_reg0   <= 36'sb1010010010000011110110001110011110;
        end
        854: begin
            cosine_reg0 <= 36'sb11110010011001001010000000001010111;
            sine_reg0   <= 36'sb1010010010110011011100011011001111;
        end
        855: begin
            cosine_reg0 <= 36'sb11110010010111001000100100101110011;
            sine_reg0   <= 36'sb1010010011100011000010001110100111;
        end
        856: begin
            cosine_reg0 <= 36'sb11110010010101000110111111111100000;
            sine_reg0   <= 36'sb1010010100010010100111101000100011;
        end
        857: begin
            cosine_reg0 <= 36'sb11110010010011000101010001110011100;
            sine_reg0   <= 36'sb1010010101000010001100101001000010;
        end
        858: begin
            cosine_reg0 <= 36'sb11110010010001000011011010010101010;
            sine_reg0   <= 36'sb1010010101110001110001010000000010;
        end
        859: begin
            cosine_reg0 <= 36'sb11110010001111000001011001100001010;
            sine_reg0   <= 36'sb1010010110100001010101011101100001;
        end
        860: begin
            cosine_reg0 <= 36'sb11110010001100111111001111010111100;
            sine_reg0   <= 36'sb1010010111010000111001010001011101;
        end
        861: begin
            cosine_reg0 <= 36'sb11110010001010111100111011111000001;
            sine_reg0   <= 36'sb1010011000000000011100101011110101;
        end
        862: begin
            cosine_reg0 <= 36'sb11110010001000111010011111000011010;
            sine_reg0   <= 36'sb1010011000101111111111101100100110;
        end
        863: begin
            cosine_reg0 <= 36'sb11110010000110110111111000111001000;
            sine_reg0   <= 36'sb1010011001011111100010010011110000;
        end
        864: begin
            cosine_reg0 <= 36'sb11110010000100110101001001011001010;
            sine_reg0   <= 36'sb1010011010001111000100100001001111;
        end
        865: begin
            cosine_reg0 <= 36'sb11110010000010110010010000100100010;
            sine_reg0   <= 36'sb1010011010111110100110010101000010;
        end
        866: begin
            cosine_reg0 <= 36'sb11110010000000101111001110011010000;
            sine_reg0   <= 36'sb1010011011101110000111101111001000;
        end
        867: begin
            cosine_reg0 <= 36'sb11110001111110101100000010111010101;
            sine_reg0   <= 36'sb1010011100011101101000101111011110;
        end
        868: begin
            cosine_reg0 <= 36'sb11110001111100101000101110000110010;
            sine_reg0   <= 36'sb1010011101001101001001010110000010;
        end
        869: begin
            cosine_reg0 <= 36'sb11110001111010100101001111111100111;
            sine_reg0   <= 36'sb1010011101111100101001100010110100;
        end
        870: begin
            cosine_reg0 <= 36'sb11110001111000100001101000011110100;
            sine_reg0   <= 36'sb1010011110101100001001010101110000;
        end
        871: begin
            cosine_reg0 <= 36'sb11110001110110011101110111101011011;
            sine_reg0   <= 36'sb1010011111011011101000101110110110;
        end
        872: begin
            cosine_reg0 <= 36'sb11110001110100011001111101100011101;
            sine_reg0   <= 36'sb1010100000001011000111101110000011;
        end
        873: begin
            cosine_reg0 <= 36'sb11110001110010010101111010000111000;
            sine_reg0   <= 36'sb1010100000111010100110010011010101;
        end
        874: begin
            cosine_reg0 <= 36'sb11110001110000010001101101010101111;
            sine_reg0   <= 36'sb1010100001101010000100011110101011;
        end
        875: begin
            cosine_reg0 <= 36'sb11110001101110001101010111010000010;
            sine_reg0   <= 36'sb1010100010011001100010010000000011;
        end
        876: begin
            cosine_reg0 <= 36'sb11110001101100001000110111110110010;
            sine_reg0   <= 36'sb1010100011001000111111100111011011;
        end
        877: begin
            cosine_reg0 <= 36'sb11110001101010000100001111000111111;
            sine_reg0   <= 36'sb1010100011111000011100100100110001;
        end
        878: begin
            cosine_reg0 <= 36'sb11110001100111111111011101000101010;
            sine_reg0   <= 36'sb1010100100100111111001001000000011;
        end
        879: begin
            cosine_reg0 <= 36'sb11110001100101111010100001101110011;
            sine_reg0   <= 36'sb1010100101010111010101010001010000;
        end
        880: begin
            cosine_reg0 <= 36'sb11110001100011110101011101000011011;
            sine_reg0   <= 36'sb1010100110000110110001000000010110;
        end
        881: begin
            cosine_reg0 <= 36'sb11110001100001110000001111000100011;
            sine_reg0   <= 36'sb1010100110110110001100010101010010;
        end
        882: begin
            cosine_reg0 <= 36'sb11110001011111101010110111110001100;
            sine_reg0   <= 36'sb1010100111100101100111010000000011;
        end
        883: begin
            cosine_reg0 <= 36'sb11110001011101100101010111001010110;
            sine_reg0   <= 36'sb1010101000010101000001110000101000;
        end
        884: begin
            cosine_reg0 <= 36'sb11110001011011011111101101010000001;
            sine_reg0   <= 36'sb1010101001000100011011110110111110;
        end
        885: begin
            cosine_reg0 <= 36'sb11110001011001011001111010000001111;
            sine_reg0   <= 36'sb1010101001110011110101100011000011;
        end
        886: begin
            cosine_reg0 <= 36'sb11110001010111010011111101100000000;
            sine_reg0   <= 36'sb1010101010100011001110110100110110;
        end
        887: begin
            cosine_reg0 <= 36'sb11110001010101001101110111101010101;
            sine_reg0   <= 36'sb1010101011010010100111101100010101;
        end
        888: begin
            cosine_reg0 <= 36'sb11110001010011000111101000100001101;
            sine_reg0   <= 36'sb1010101100000010000000001001011110;
        end
        889: begin
            cosine_reg0 <= 36'sb11110001010001000001010000000101011;
            sine_reg0   <= 36'sb1010101100110001011000001100001111;
        end
        890: begin
            cosine_reg0 <= 36'sb11110001001110111010101110010101110;
            sine_reg0   <= 36'sb1010101101100000101111110100100111;
        end
        891: begin
            cosine_reg0 <= 36'sb11110001001100110100000011010011000;
            sine_reg0   <= 36'sb1010101110010000000111000010100011;
        end
        892: begin
            cosine_reg0 <= 36'sb11110001001010101101001110111101001;
            sine_reg0   <= 36'sb1010101110111111011101110110000010;
        end
        893: begin
            cosine_reg0 <= 36'sb11110001001000100110010001010100001;
            sine_reg0   <= 36'sb1010101111101110110100001111000010;
        end
        894: begin
            cosine_reg0 <= 36'sb11110001000110011111001010011000001;
            sine_reg0   <= 36'sb1010110000011110001010001101100001;
        end
        895: begin
            cosine_reg0 <= 36'sb11110001000100010111111010001001010;
            sine_reg0   <= 36'sb1010110001001101011111110001011101;
        end
        896: begin
            cosine_reg0 <= 36'sb11110001000010010000100000100111101;
            sine_reg0   <= 36'sb1010110001111100110100111010110101;
        end
        897: begin
            cosine_reg0 <= 36'sb11110001000000001000111101110011001;
            sine_reg0   <= 36'sb1010110010101100001001101001100110;
        end
        898: begin
            cosine_reg0 <= 36'sb11110000111110000001010001101100001;
            sine_reg0   <= 36'sb1010110011011011011101111101101111;
        end
        899: begin
            cosine_reg0 <= 36'sb11110000111011111001011100010010100;
            sine_reg0   <= 36'sb1010110100001010110001110111001110;
        end
        900: begin
            cosine_reg0 <= 36'sb11110000111001110001011101100110011;
            sine_reg0   <= 36'sb1010110100111010000101010110000010;
        end
        901: begin
            cosine_reg0 <= 36'sb11110000110111101001010101100111111;
            sine_reg0   <= 36'sb1010110101101001011000011010000111;
        end
        902: begin
            cosine_reg0 <= 36'sb11110000110101100001000100010111001;
            sine_reg0   <= 36'sb1010110110011000101011000011011101;
        end
        903: begin
            cosine_reg0 <= 36'sb11110000110011011000101001110100000;
            sine_reg0   <= 36'sb1010110111000111111101010010000010;
        end
        904: begin
            cosine_reg0 <= 36'sb11110000110001010000000101111110110;
            sine_reg0   <= 36'sb1010110111110111001111000101110011;
        end
        905: begin
            cosine_reg0 <= 36'sb11110000101111000111011000110111100;
            sine_reg0   <= 36'sb1010111000100110100000011110110000;
        end
        906: begin
            cosine_reg0 <= 36'sb11110000101100111110100010011110001;
            sine_reg0   <= 36'sb1010111001010101110001011100110110;
        end
        907: begin
            cosine_reg0 <= 36'sb11110000101010110101100010110011000;
            sine_reg0   <= 36'sb1010111010000101000010000000000011;
        end
        908: begin
            cosine_reg0 <= 36'sb11110000101000101100011001110101111;
            sine_reg0   <= 36'sb1010111010110100010010001000010110;
        end
        909: begin
            cosine_reg0 <= 36'sb11110000100110100011000111100111001;
            sine_reg0   <= 36'sb1010111011100011100001110101101100;
        end
        910: begin
            cosine_reg0 <= 36'sb11110000100100011001101100000110110;
            sine_reg0   <= 36'sb1010111100010010110001001000000100;
        end
        911: begin
            cosine_reg0 <= 36'sb11110000100010010000000111010100110;
            sine_reg0   <= 36'sb1010111101000001111111111111011101;
        end
        912: begin
            cosine_reg0 <= 36'sb11110000100000000110011001010001001;
            sine_reg0   <= 36'sb1010111101110001001110011011110011;
        end
        913: begin
            cosine_reg0 <= 36'sb11110000011101111100100001111100010;
            sine_reg0   <= 36'sb1010111110100000011100011101000111;
        end
        914: begin
            cosine_reg0 <= 36'sb11110000011011110010100001010110000;
            sine_reg0   <= 36'sb1010111111001111101010000011010100;
        end
        915: begin
            cosine_reg0 <= 36'sb11110000011001101000010111011110100;
            sine_reg0   <= 36'sb1010111111111110110111001110011011;
        end
        916: begin
            cosine_reg0 <= 36'sb11110000010111011110000100010101110;
            sine_reg0   <= 36'sb1011000000101110000011111110011001;
        end
        917: begin
            cosine_reg0 <= 36'sb11110000010101010011100111111100000;
            sine_reg0   <= 36'sb1011000001011101010000010011001100;
        end
        918: begin
            cosine_reg0 <= 36'sb11110000010011001001000010010001010;
            sine_reg0   <= 36'sb1011000010001100011100001100110010;
        end
        919: begin
            cosine_reg0 <= 36'sb11110000010000111110010011010101101;
            sine_reg0   <= 36'sb1011000010111011100111101011001001;
        end
        920: begin
            cosine_reg0 <= 36'sb11110000001110110011011011001001001;
            sine_reg0   <= 36'sb1011000011101010110010101110010001;
        end
        921: begin
            cosine_reg0 <= 36'sb11110000001100101000011001101011111;
            sine_reg0   <= 36'sb1011000100011001111101010110000110;
        end
        922: begin
            cosine_reg0 <= 36'sb11110000001010011101001110111110000;
            sine_reg0   <= 36'sb1011000101001001000111100010100111;
        end
        923: begin
            cosine_reg0 <= 36'sb11110000001000010001111010111111100;
            sine_reg0   <= 36'sb1011000101111000010001010011110011;
        end
        924: begin
            cosine_reg0 <= 36'sb11110000000110000110011101110000100;
            sine_reg0   <= 36'sb1011000110100111011010101001100111;
        end
        925: begin
            cosine_reg0 <= 36'sb11110000000011111010110111010001001;
            sine_reg0   <= 36'sb1011000111010110100011100100000010;
        end
        926: begin
            cosine_reg0 <= 36'sb11110000000001101111000111100001011;
            sine_reg0   <= 36'sb1011001000000101101100000011000001;
        end
        927: begin
            cosine_reg0 <= 36'sb11101111111111100011001110100001011;
            sine_reg0   <= 36'sb1011001000110100110100000110100100;
        end
        928: begin
            cosine_reg0 <= 36'sb11101111111101010111001100010001010;
            sine_reg0   <= 36'sb1011001001100011111011101110101000;
        end
        929: begin
            cosine_reg0 <= 36'sb11101111111011001011000000110001001;
            sine_reg0   <= 36'sb1011001010010011000010111011001011;
        end
        930: begin
            cosine_reg0 <= 36'sb11101111111000111110101100000000111;
            sine_reg0   <= 36'sb1011001011000010001001101100001011;
        end
        931: begin
            cosine_reg0 <= 36'sb11101111110110110010001110000000111;
            sine_reg0   <= 36'sb1011001011110001010000000001100111;
        end
        932: begin
            cosine_reg0 <= 36'sb11101111110100100101100110110000111;
            sine_reg0   <= 36'sb1011001100100000010101111011011110;
        end
        933: begin
            cosine_reg0 <= 36'sb11101111110010011000110110010001010;
            sine_reg0   <= 36'sb1011001101001111011011011001101100;
        end
        934: begin
            cosine_reg0 <= 36'sb11101111110000001011111100100010000;
            sine_reg0   <= 36'sb1011001101111110100000011100010001;
        end
        935: begin
            cosine_reg0 <= 36'sb11101111101101111110111001100011001;
            sine_reg0   <= 36'sb1011001110101101100101000011001010;
        end
        936: begin
            cosine_reg0 <= 36'sb11101111101011110001101101010100110;
            sine_reg0   <= 36'sb1011001111011100101001001110010101;
        end
        937: begin
            cosine_reg0 <= 36'sb11101111101001100100010111110111000;
            sine_reg0   <= 36'sb1011010000001011101100111101110010;
        end
        938: begin
            cosine_reg0 <= 36'sb11101111100111010110111001001010000;
            sine_reg0   <= 36'sb1011010000111010110000010001011101;
        end
        939: begin
            cosine_reg0 <= 36'sb11101111100101001001010001001101101;
            sine_reg0   <= 36'sb1011010001101001110011001001010110;
        end
        940: begin
            cosine_reg0 <= 36'sb11101111100010111011100000000010010;
            sine_reg0   <= 36'sb1011010010011000110101100101011010;
        end
        941: begin
            cosine_reg0 <= 36'sb11101111100000101101100101100111110;
            sine_reg0   <= 36'sb1011010011000111110111100101101000;
        end
        942: begin
            cosine_reg0 <= 36'sb11101111011110011111100001111110010;
            sine_reg0   <= 36'sb1011010011110110111001001001111110;
        end
        943: begin
            cosine_reg0 <= 36'sb11101111011100010001010101000110000;
            sine_reg0   <= 36'sb1011010100100101111010010010011001;
        end
        944: begin
            cosine_reg0 <= 36'sb11101111011010000010111110111110111;
            sine_reg0   <= 36'sb1011010101010100111010111110111001;
        end
        945: begin
            cosine_reg0 <= 36'sb11101111010111110100011111101001000;
            sine_reg0   <= 36'sb1011010110000011111011001111011010;
        end
        946: begin
            cosine_reg0 <= 36'sb11101111010101100101110111000100100;
            sine_reg0   <= 36'sb1011010110110010111011000011111101;
        end
        947: begin
            cosine_reg0 <= 36'sb11101111010011010111000101010001100;
            sine_reg0   <= 36'sb1011010111100001111010011100011110;
        end
        948: begin
            cosine_reg0 <= 36'sb11101111010001001000001010010000000;
            sine_reg0   <= 36'sb1011011000010000111001011000111100;
        end
        949: begin
            cosine_reg0 <= 36'sb11101111001110111001000110000000001;
            sine_reg0   <= 36'sb1011011000111111110111111001010101;
        end
        950: begin
            cosine_reg0 <= 36'sb11101111001100101001111000100010000;
            sine_reg0   <= 36'sb1011011001101110110101111101101000;
        end
        951: begin
            cosine_reg0 <= 36'sb11101111001010011010100001110101110;
            sine_reg0   <= 36'sb1011011010011101110011100101110001;
        end
        952: begin
            cosine_reg0 <= 36'sb11101111001000001011000001111011010;
            sine_reg0   <= 36'sb1011011011001100110000110001110001;
        end
        953: begin
            cosine_reg0 <= 36'sb11101111000101111011011000110010111;
            sine_reg0   <= 36'sb1011011011111011101101100001100100;
        end
        954: begin
            cosine_reg0 <= 36'sb11101111000011101011100110011100100;
            sine_reg0   <= 36'sb1011011100101010101001110101001010;
        end
        955: begin
            cosine_reg0 <= 36'sb11101111000001011011101010111000010;
            sine_reg0   <= 36'sb1011011101011001100101101100011111;
        end
        956: begin
            cosine_reg0 <= 36'sb11101110111111001011100110000110010;
            sine_reg0   <= 36'sb1011011110001000100001000111100011;
        end
        957: begin
            cosine_reg0 <= 36'sb11101110111100111011011000000110100;
            sine_reg0   <= 36'sb1011011110110111011100000110010100;
        end
        958: begin
            cosine_reg0 <= 36'sb11101110111010101011000000111001010;
            sine_reg0   <= 36'sb1011011111100110010110101000101111;
        end
        959: begin
            cosine_reg0 <= 36'sb11101110111000011010100000011110100;
            sine_reg0   <= 36'sb1011100000010101010000101110110011;
        end
        960: begin
            cosine_reg0 <= 36'sb11101110110110001001110110110110010;
            sine_reg0   <= 36'sb1011100001000100001010011000011111;
        end
        961: begin
            cosine_reg0 <= 36'sb11101110110011111001000100000000110;
            sine_reg0   <= 36'sb1011100001110011000011100101110000;
        end
        962: begin
            cosine_reg0 <= 36'sb11101110110001101000000111111110000;
            sine_reg0   <= 36'sb1011100010100001111100010110100100;
        end
        963: begin
            cosine_reg0 <= 36'sb11101110101111010111000010101110001;
            sine_reg0   <= 36'sb1011100011010000110100101010111010;
        end
        964: begin
            cosine_reg0 <= 36'sb11101110101101000101110100010001001;
            sine_reg0   <= 36'sb1011100011111111101100100010110001;
        end
        965: begin
            cosine_reg0 <= 36'sb11101110101010110100011100100111001;
            sine_reg0   <= 36'sb1011100100101110100011111110000101;
        end
        966: begin
            cosine_reg0 <= 36'sb11101110101000100010111011110000010;
            sine_reg0   <= 36'sb1011100101011101011010111100110101;
        end
        967: begin
            cosine_reg0 <= 36'sb11101110100110010001010001101100101;
            sine_reg0   <= 36'sb1011100110001100010001011111000001;
        end
        968: begin
            cosine_reg0 <= 36'sb11101110100011111111011110011100010;
            sine_reg0   <= 36'sb1011100110111011000111100100100100;
        end
        969: begin
            cosine_reg0 <= 36'sb11101110100001101101100001111111010;
            sine_reg0   <= 36'sb1011100111101001111101001101011111;
        end
        970: begin
            cosine_reg0 <= 36'sb11101110011111011011011100010101101;
            sine_reg0   <= 36'sb1011101000011000110010011001101111;
        end
        971: begin
            cosine_reg0 <= 36'sb11101110011101001001001101011111101;
            sine_reg0   <= 36'sb1011101001000111100111001001010010;
        end
        972: begin
            cosine_reg0 <= 36'sb11101110011010110110110101011101010;
            sine_reg0   <= 36'sb1011101001110110011011011100000111;
        end
        973: begin
            cosine_reg0 <= 36'sb11101110011000100100010100001110101;
            sine_reg0   <= 36'sb1011101010100101001111010010001011;
        end
        974: begin
            cosine_reg0 <= 36'sb11101110010110010001101001110011110;
            sine_reg0   <= 36'sb1011101011010100000010101011011101;
        end
        975: begin
            cosine_reg0 <= 36'sb11101110010011111110110110001100111;
            sine_reg0   <= 36'sb1011101100000010110101100111111100;
        end
        976: begin
            cosine_reg0 <= 36'sb11101110010001101011111001011001111;
            sine_reg0   <= 36'sb1011101100110001101000000111100100;
        end
        977: begin
            cosine_reg0 <= 36'sb11101110001111011000110011011011000;
            sine_reg0   <= 36'sb1011101101100000011010001010010101;
        end
        978: begin
            cosine_reg0 <= 36'sb11101110001101000101100100010000011;
            sine_reg0   <= 36'sb1011101110001111001011110000001101;
        end
        979: begin
            cosine_reg0 <= 36'sb11101110001010110010001011111001111;
            sine_reg0   <= 36'sb1011101110111101111100111001001001;
        end
        980: begin
            cosine_reg0 <= 36'sb11101110001000011110101010010111110;
            sine_reg0   <= 36'sb1011101111101100101101100101001001;
        end
        981: begin
            cosine_reg0 <= 36'sb11101110000110001010111111101010001;
            sine_reg0   <= 36'sb1011110000011011011101110100001010;
        end
        982: begin
            cosine_reg0 <= 36'sb11101110000011110111001011110001000;
            sine_reg0   <= 36'sb1011110001001010001101100110001010;
        end
        983: begin
            cosine_reg0 <= 36'sb11101110000001100011001110101100011;
            sine_reg0   <= 36'sb1011110001111000111100111011001000;
        end
        984: begin
            cosine_reg0 <= 36'sb11101101111111001111001000011100100;
            sine_reg0   <= 36'sb1011110010100111101011110011000010;
        end
        985: begin
            cosine_reg0 <= 36'sb11101101111100111010111001000001100;
            sine_reg0   <= 36'sb1011110011010110011010001101110110;
        end
        986: begin
            cosine_reg0 <= 36'sb11101101111010100110100000011011011;
            sine_reg0   <= 36'sb1011110100000101001000001011100010;
        end
        987: begin
            cosine_reg0 <= 36'sb11101101111000010001111110101010001;
            sine_reg0   <= 36'sb1011110100110011110101101100000101;
        end
        988: begin
            cosine_reg0 <= 36'sb11101101110101111101010011101110000;
            sine_reg0   <= 36'sb1011110101100010100010101111011100;
        end
        989: begin
            cosine_reg0 <= 36'sb11101101110011101000011111100110111;
            sine_reg0   <= 36'sb1011110110010001001111010101100110;
        end
        990: begin
            cosine_reg0 <= 36'sb11101101110001010011100010010101001;
            sine_reg0   <= 36'sb1011110110111111111011011110100001;
        end
        991: begin
            cosine_reg0 <= 36'sb11101101101110111110011011111000110;
            sine_reg0   <= 36'sb1011110111101110100111001010001100;
        end
        992: begin
            cosine_reg0 <= 36'sb11101101101100101001001100010001101;
            sine_reg0   <= 36'sb1011111000011101010010011000100011;
        end
        993: begin
            cosine_reg0 <= 36'sb11101101101010010011110011100000001;
            sine_reg0   <= 36'sb1011111001001011111101001001100111;
        end
        994: begin
            cosine_reg0 <= 36'sb11101101100111111110010001100100001;
            sine_reg0   <= 36'sb1011111001111010100111011101010100;
        end
        995: begin
            cosine_reg0 <= 36'sb11101101100101101000100110011101111;
            sine_reg0   <= 36'sb1011111010101001010001010011101001;
        end
        996: begin
            cosine_reg0 <= 36'sb11101101100011010010110010001101100;
            sine_reg0   <= 36'sb1011111011010111111010101100100101;
        end
        997: begin
            cosine_reg0 <= 36'sb11101101100000111100110100110010111;
            sine_reg0   <= 36'sb1011111100000110100011101000000101;
        end
        998: begin
            cosine_reg0 <= 36'sb11101101011110100110101110001110001;
            sine_reg0   <= 36'sb1011111100110101001100000110001000;
        end
        999: begin
            cosine_reg0 <= 36'sb11101101011100010000011110011111101;
            sine_reg0   <= 36'sb1011111101100011110100000110101011;
        end
        1000: begin
            cosine_reg0 <= 36'sb11101101011001111010000101100111001;
            sine_reg0   <= 36'sb1011111110010010011011101001101110;
        end
        1001: begin
            cosine_reg0 <= 36'sb11101101010111100011100011100100111;
            sine_reg0   <= 36'sb1011111111000001000010101111001110;
        end
        1002: begin
            cosine_reg0 <= 36'sb11101101010101001100111000011000111;
            sine_reg0   <= 36'sb1011111111101111101001010111001001;
        end
        1003: begin
            cosine_reg0 <= 36'sb11101101010010110110000100000011011;
            sine_reg0   <= 36'sb1100000000011110001111100001011110;
        end
        1004: begin
            cosine_reg0 <= 36'sb11101101010000011111000110100100011;
            sine_reg0   <= 36'sb1100000001001100110101001110001011;
        end
        1005: begin
            cosine_reg0 <= 36'sb11101101001110000111111111111011111;
            sine_reg0   <= 36'sb1100000001111011011010011101001110;
        end
        1006: begin
            cosine_reg0 <= 36'sb11101101001011110000110000001010001;
            sine_reg0   <= 36'sb1100000010101001111111001110100101;
        end
        1007: begin
            cosine_reg0 <= 36'sb11101101001001011001010111001111010;
            sine_reg0   <= 36'sb1100000011011000100011100010001111;
        end
        1008: begin
            cosine_reg0 <= 36'sb11101101000111000001110101001011001;
            sine_reg0   <= 36'sb1100000100000111000111011000001001;
        end
        1009: begin
            cosine_reg0 <= 36'sb11101101000100101010001001111101111;
            sine_reg0   <= 36'sb1100000100110101101010110000010011;
        end
        1010: begin
            cosine_reg0 <= 36'sb11101101000010010010010101100111111;
            sine_reg0   <= 36'sb1100000101100100001101101010101001;
        end
        1011: begin
            cosine_reg0 <= 36'sb11101100111111111010011000001000111;
            sine_reg0   <= 36'sb1100000110010010110000000111001011;
        end
        1012: begin
            cosine_reg0 <= 36'sb11101100111101100010010001100001001;
            sine_reg0   <= 36'sb1100000111000001010010000101110110;
        end
        1013: begin
            cosine_reg0 <= 36'sb11101100111011001010000001110000101;
            sine_reg0   <= 36'sb1100000111101111110011100110101001;
        end
        1014: begin
            cosine_reg0 <= 36'sb11101100111000110001101000110111101;
            sine_reg0   <= 36'sb1100001000011110010100101001100010;
        end
        1015: begin
            cosine_reg0 <= 36'sb11101100110110011001000110110110001;
            sine_reg0   <= 36'sb1100001001001100110101001110011111;
        end
        1016: begin
            cosine_reg0 <= 36'sb11101100110100000000011011101100010;
            sine_reg0   <= 36'sb1100001001111011010101010101011110;
        end
        1017: begin
            cosine_reg0 <= 36'sb11101100110001100111100111011010000;
            sine_reg0   <= 36'sb1100001010101001110100111110011110;
        end
        1018: begin
            cosine_reg0 <= 36'sb11101100101111001110101001111111101;
            sine_reg0   <= 36'sb1100001011011000010100001001011101;
        end
        1019: begin
            cosine_reg0 <= 36'sb11101100101100110101100011011101000;
            sine_reg0   <= 36'sb1100001100000110110010110110011000;
        end
        1020: begin
            cosine_reg0 <= 36'sb11101100101010011100010011110010011;
            sine_reg0   <= 36'sb1100001100110101010001000101001111;
        end
        1021: begin
            cosine_reg0 <= 36'sb11101100101000000010111010111111111;
            sine_reg0   <= 36'sb1100001101100011101110110101111111;
        end
        1022: begin
            cosine_reg0 <= 36'sb11101100100101101001011001000101100;
            sine_reg0   <= 36'sb1100001110010010001100001000100111;
        end
        1023: begin
            cosine_reg0 <= 36'sb11101100100011001111101110000011010;
            sine_reg0   <= 36'sb1100001111000000101000111101000100;
        end
        1024: begin
            cosine_reg0 <= 36'sb11101100100000110101111001111001100;
            sine_reg0   <= 36'sb1100001111101111000101010011010101;
        end
        1025: begin
            cosine_reg0 <= 36'sb11101100011110011011111100101000001;
            sine_reg0   <= 36'sb1100010000011101100001001011011001;
        end
        1026: begin
            cosine_reg0 <= 36'sb11101100011100000001110110001111010;
            sine_reg0   <= 36'sb1100010001001011111100100101001101;
        end
        1027: begin
            cosine_reg0 <= 36'sb11101100011001100111100110101110111;
            sine_reg0   <= 36'sb1100010001111010010111100000110000;
        end
        1028: begin
            cosine_reg0 <= 36'sb11101100010111001101001110000111011;
            sine_reg0   <= 36'sb1100010010101000110001111101111111;
        end
        1029: begin
            cosine_reg0 <= 36'sb11101100010100110010101100011000101;
            sine_reg0   <= 36'sb1100010011010111001011111100111010;
        end
        1030: begin
            cosine_reg0 <= 36'sb11101100010010011000000001100010110;
            sine_reg0   <= 36'sb1100010100000101100101011101011110;
        end
        1031: begin
            cosine_reg0 <= 36'sb11101100001111111101001101100101111;
            sine_reg0   <= 36'sb1100010100110011111110011111101001;
        end
        1032: begin
            cosine_reg0 <= 36'sb11101100001101100010010000100010000;
            sine_reg0   <= 36'sb1100010101100010010111000011011010;
        end
        1033: begin
            cosine_reg0 <= 36'sb11101100001011000111001010010111011;
            sine_reg0   <= 36'sb1100010110010000101111001000101111;
        end
        1034: begin
            cosine_reg0 <= 36'sb11101100001000101011111011000110000;
            sine_reg0   <= 36'sb1100010110111111000110101111100110;
        end
        1035: begin
            cosine_reg0 <= 36'sb11101100000110010000100010101110000;
            sine_reg0   <= 36'sb1100010111101101011101110111111110;
        end
        1036: begin
            cosine_reg0 <= 36'sb11101100000011110101000001001111100;
            sine_reg0   <= 36'sb1100011000011011110100100001110100;
        end
        1037: begin
            cosine_reg0 <= 36'sb11101100000001011001010110101010100;
            sine_reg0   <= 36'sb1100011001001010001010101101000110;
        end
        1038: begin
            cosine_reg0 <= 36'sb11101011111110111101100010111111001;
            sine_reg0   <= 36'sb1100011001111000100000011001110100;
        end
        1039: begin
            cosine_reg0 <= 36'sb11101011111100100001100110001101100;
            sine_reg0   <= 36'sb1100011010100110110101100111111011;
        end
        1040: begin
            cosine_reg0 <= 36'sb11101011111010000101100000010101101;
            sine_reg0   <= 36'sb1100011011010101001010010111011001;
        end
        1041: begin
            cosine_reg0 <= 36'sb11101011110111101001010001010111110;
            sine_reg0   <= 36'sb1100011100000011011110101000001100;
        end
        1042: begin
            cosine_reg0 <= 36'sb11101011110101001100111001010011111;
            sine_reg0   <= 36'sb1100011100110001110010011010010100;
        end
        1043: begin
            cosine_reg0 <= 36'sb11101011110010110000011000001010001;
            sine_reg0   <= 36'sb1100011101100000000101101101101110;
        end
        1044: begin
            cosine_reg0 <= 36'sb11101011110000010011101101111010101;
            sine_reg0   <= 36'sb1100011110001110011000100010010111;
        end
        1045: begin
            cosine_reg0 <= 36'sb11101011101101110110111010100101011;
            sine_reg0   <= 36'sb1100011110111100101010111000010000;
        end
        1046: begin
            cosine_reg0 <= 36'sb11101011101011011001111110001010100;
            sine_reg0   <= 36'sb1100011111101010111100101111010101;
        end
        1047: begin
            cosine_reg0 <= 36'sb11101011101000111100111000101010000;
            sine_reg0   <= 36'sb1100100000011001001110000111100101;
        end
        1048: begin
            cosine_reg0 <= 36'sb11101011100110011111101010000100010;
            sine_reg0   <= 36'sb1100100001000111011111000000111110;
        end
        1049: begin
            cosine_reg0 <= 36'sb11101011100100000010010010011001001;
            sine_reg0   <= 36'sb1100100001110101101111011011011110;
        end
        1050: begin
            cosine_reg0 <= 36'sb11101011100001100100110001101000110;
            sine_reg0   <= 36'sb1100100010100011111111010111000100;
        end
        1051: begin
            cosine_reg0 <= 36'sb11101011011111000111000111110011010;
            sine_reg0   <= 36'sb1100100011010010001110110011101101;
        end
        1052: begin
            cosine_reg0 <= 36'sb11101011011100101001010100111000110;
            sine_reg0   <= 36'sb1100100100000000011101110001011001;
        end
        1053: begin
            cosine_reg0 <= 36'sb11101011011010001011011000111001010;
            sine_reg0   <= 36'sb1100100100101110101100010000000101;
        end
        1054: begin
            cosine_reg0 <= 36'sb11101011010111101101010011110101000;
            sine_reg0   <= 36'sb1100100101011100111010001111101111;
        end
        1055: begin
            cosine_reg0 <= 36'sb11101011010101001111000101101011111;
            sine_reg0   <= 36'sb1100100110001011000111110000010110;
        end
        1056: begin
            cosine_reg0 <= 36'sb11101011010010110000101110011110010;
            sine_reg0   <= 36'sb1100100110111001010100110001110111;
        end
        1057: begin
            cosine_reg0 <= 36'sb11101011010000010010001110001011111;
            sine_reg0   <= 36'sb1100100111100111100001010100010010;
        end
        1058: begin
            cosine_reg0 <= 36'sb11101011001101110011100100110101001;
            sine_reg0   <= 36'sb1100101000010101101101010111100100;
        end
        1059: begin
            cosine_reg0 <= 36'sb11101011001011010100110010011010000;
            sine_reg0   <= 36'sb1100101001000011111000111011101011;
        end
        1060: begin
            cosine_reg0 <= 36'sb11101011001000110101110110111010101;
            sine_reg0   <= 36'sb1100101001110010000100000000100111;
        end
        1061: begin
            cosine_reg0 <= 36'sb11101011000110010110110010010111000;
            sine_reg0   <= 36'sb1100101010100000001110100110010100;
        end
        1062: begin
            cosine_reg0 <= 36'sb11101011000011110111100100101111011;
            sine_reg0   <= 36'sb1100101011001110011000101100110001;
        end
        1063: begin
            cosine_reg0 <= 36'sb11101011000001011000001110000011110;
            sine_reg0   <= 36'sb1100101011111100100010010011111101;
        end
        1064: begin
            cosine_reg0 <= 36'sb11101010111110111000101110010100001;
            sine_reg0   <= 36'sb1100101100101010101011011011110101;
        end
        1065: begin
            cosine_reg0 <= 36'sb11101010111100011001000101100000110;
            sine_reg0   <= 36'sb1100101101011000110100000100011000;
        end
        1066: begin
            cosine_reg0 <= 36'sb11101010111001111001010011101001110;
            sine_reg0   <= 36'sb1100101110000110111100001101100100;
        end
        1067: begin
            cosine_reg0 <= 36'sb11101010110111011001011000101111001;
            sine_reg0   <= 36'sb1100101110110101000011110111011000;
        end
        1068: begin
            cosine_reg0 <= 36'sb11101010110100111001010100110001000;
            sine_reg0   <= 36'sb1100101111100011001011000001110001;
        end
        1069: begin
            cosine_reg0 <= 36'sb11101010110010011001000111101111011;
            sine_reg0   <= 36'sb1100110000010001010001101100101101;
        end
        1070: begin
            cosine_reg0 <= 36'sb11101010101111111000110001101010100;
            sine_reg0   <= 36'sb1100110000111111010111111000001100;
        end
        1071: begin
            cosine_reg0 <= 36'sb11101010101101011000010010100010011;
            sine_reg0   <= 36'sb1100110001101101011101100100001011;
        end
        1072: begin
            cosine_reg0 <= 36'sb11101010101010110111101010010111001;
            sine_reg0   <= 36'sb1100110010011011100010110000101000;
        end
        1073: begin
            cosine_reg0 <= 36'sb11101010101000010110111001001000111;
            sine_reg0   <= 36'sb1100110011001001100111011101100010;
        end
        1074: begin
            cosine_reg0 <= 36'sb11101010100101110101111110110111110;
            sine_reg0   <= 36'sb1100110011110111101011101010110110;
        end
        1075: begin
            cosine_reg0 <= 36'sb11101010100011010100111011100011110;
            sine_reg0   <= 36'sb1100110100100101101111011000100100;
        end
        1076: begin
            cosine_reg0 <= 36'sb11101010100000110011101111001101000;
            sine_reg0   <= 36'sb1100110101010011110010100110101001;
        end
        1077: begin
            cosine_reg0 <= 36'sb11101010011110010010011001110011101;
            sine_reg0   <= 36'sb1100110110000001110101010101000011;
        end
        1078: begin
            cosine_reg0 <= 36'sb11101010011011110000111011010111110;
            sine_reg0   <= 36'sb1100110110101111110111100011110001;
        end
        1079: begin
            cosine_reg0 <= 36'sb11101010011001001111010011111001011;
            sine_reg0   <= 36'sb1100110111011101111001010010110001;
        end
        1080: begin
            cosine_reg0 <= 36'sb11101010010110101101100011011000101;
            sine_reg0   <= 36'sb1100111000001011111010100010000001;
        end
        1081: begin
            cosine_reg0 <= 36'sb11101010010100001011101001110101110;
            sine_reg0   <= 36'sb1100111000111001111011010001100000;
        end
        1082: begin
            cosine_reg0 <= 36'sb11101010010001101001100111010000101;
            sine_reg0   <= 36'sb1100111001100111111011100001001011;
        end
        1083: begin
            cosine_reg0 <= 36'sb11101010001111000111011011101001100;
            sine_reg0   <= 36'sb1100111010010101111011010001000001;
        end
        1084: begin
            cosine_reg0 <= 36'sb11101010001100100101000111000000011;
            sine_reg0   <= 36'sb1100111011000011111010100001000001;
        end
        1085: begin
            cosine_reg0 <= 36'sb11101010001010000010101001010101011;
            sine_reg0   <= 36'sb1100111011110001111001010001000111;
        end
        1086: begin
            cosine_reg0 <= 36'sb11101010000111100000000010101000101;
            sine_reg0   <= 36'sb1100111100011111110111100001010011;
        end
        1087: begin
            cosine_reg0 <= 36'sb11101010000100111101010010111010010;
            sine_reg0   <= 36'sb1100111101001101110101010001100011;
        end
        1088: begin
            cosine_reg0 <= 36'sb11101010000010011010011010001010011;
            sine_reg0   <= 36'sb1100111101111011110010100001110101;
        end
        1089: begin
            cosine_reg0 <= 36'sb11101001111111110111011000011000111;
            sine_reg0   <= 36'sb1100111110101001101111010010000111;
        end
        1090: begin
            cosine_reg0 <= 36'sb11101001111101010100001101100110001;
            sine_reg0   <= 36'sb1100111111010111101011100010010111;
        end
        1091: begin
            cosine_reg0 <= 36'sb11101001111010110000111001110010001;
            sine_reg0   <= 36'sb1101000000000101100111010010100100;
        end
        1092: begin
            cosine_reg0 <= 36'sb11101001111000001101011100111100111;
            sine_reg0   <= 36'sb1101000000110011100010100010101100;
        end
        1093: begin
            cosine_reg0 <= 36'sb11101001110101101001110111000110101;
            sine_reg0   <= 36'sb1101000001100001011101010010101110;
        end
        1094: begin
            cosine_reg0 <= 36'sb11101001110011000110001000001111010;
            sine_reg0   <= 36'sb1101000010001111010111100010100110;
        end
        1095: begin
            cosine_reg0 <= 36'sb11101001110000100010010000010111001;
            sine_reg0   <= 36'sb1101000010111101010001010010010100;
        end
        1096: begin
            cosine_reg0 <= 36'sb11101001101101111110001111011110010;
            sine_reg0   <= 36'sb1101000011101011001010100001110110;
        end
        1097: begin
            cosine_reg0 <= 36'sb11101001101011011010000101100100101;
            sine_reg0   <= 36'sb1101000100011001000011010001001010;
        end
        1098: begin
            cosine_reg0 <= 36'sb11101001101000110101110010101010100;
            sine_reg0   <= 36'sb1101000101000110111011100000001111;
        end
        1099: begin
            cosine_reg0 <= 36'sb11101001100110010001010110101111111;
            sine_reg0   <= 36'sb1101000101110100110011001111000001;
        end
        1100: begin
            cosine_reg0 <= 36'sb11101001100011101100110001110100111;
            sine_reg0   <= 36'sb1101000110100010101010011101100001;
        end
        1101: begin
            cosine_reg0 <= 36'sb11101001100001001000000011111001100;
            sine_reg0   <= 36'sb1101000111010000100001001011101100;
        end
        1102: begin
            cosine_reg0 <= 36'sb11101001011110100011001100111110000;
            sine_reg0   <= 36'sb1101000111111110010111011001011111;
        end
        1103: begin
            cosine_reg0 <= 36'sb11101001011011111110001101000010100;
            sine_reg0   <= 36'sb1101001000101100001101000110111011;
        end
        1104: begin
            cosine_reg0 <= 36'sb11101001011001011001000100000110111;
            sine_reg0   <= 36'sb1101001001011010000010010011111011;
        end
        1105: begin
            cosine_reg0 <= 36'sb11101001010110110011110010001011100;
            sine_reg0   <= 36'sb1101001010000111110111000000100000;
        end
        1106: begin
            cosine_reg0 <= 36'sb11101001010100001110010111010000010;
            sine_reg0   <= 36'sb1101001010110101101011001100100111;
        end
        1107: begin
            cosine_reg0 <= 36'sb11101001010001101000110011010101011;
            sine_reg0   <= 36'sb1101001011100011011110111000001111;
        end
        1108: begin
            cosine_reg0 <= 36'sb11101001001111000011000110011010111;
            sine_reg0   <= 36'sb1101001100010001010010000011010100;
        end
        1109: begin
            cosine_reg0 <= 36'sb11101001001100011101010000100000111;
            sine_reg0   <= 36'sb1101001100111111000100101101110111;
        end
        1110: begin
            cosine_reg0 <= 36'sb11101001001001110111010001100111100;
            sine_reg0   <= 36'sb1101001101101100110110110111110101;
        end
        1111: begin
            cosine_reg0 <= 36'sb11101001000111010001001001101110111;
            sine_reg0   <= 36'sb1101001110011010101000100001001100;
        end
        1112: begin
            cosine_reg0 <= 36'sb11101001000100101010111000110111001;
            sine_reg0   <= 36'sb1101001111001000011001101001111011;
        end
        1113: begin
            cosine_reg0 <= 36'sb11101001000010000100011111000000001;
            sine_reg0   <= 36'sb1101001111110110001010010010000000;
        end
        1114: begin
            cosine_reg0 <= 36'sb11101000111111011101111100001010010;
            sine_reg0   <= 36'sb1101010000100011111010011001011000;
        end
        1115: begin
            cosine_reg0 <= 36'sb11101000111100110111010000010101100;
            sine_reg0   <= 36'sb1101010001010001101010000000000011;
        end
        1116: begin
            cosine_reg0 <= 36'sb11101000111010010000011011100001111;
            sine_reg0   <= 36'sb1101010001111111011001000101111110;
        end
        1117: begin
            cosine_reg0 <= 36'sb11101000110111101001011101101111101;
            sine_reg0   <= 36'sb1101010010101101000111101011001000;
        end
        1118: begin
            cosine_reg0 <= 36'sb11101000110101000010010110111110111;
            sine_reg0   <= 36'sb1101010011011010110101101111011111;
        end
        1119: begin
            cosine_reg0 <= 36'sb11101000110010011011000111001111100;
            sine_reg0   <= 36'sb1101010100001000100011010011000010;
        end
        1120: begin
            cosine_reg0 <= 36'sb11101000101111110011101110100001111;
            sine_reg0   <= 36'sb1101010100110110010000010101101101;
        end
        1121: begin
            cosine_reg0 <= 36'sb11101000101101001100001100110101111;
            sine_reg0   <= 36'sb1101010101100011111100110111100001;
        end
        1122: begin
            cosine_reg0 <= 36'sb11101000101010100100100010001011110;
            sine_reg0   <= 36'sb1101010110010001101000111000011010;
        end
        1123: begin
            cosine_reg0 <= 36'sb11101000100111111100101110100011100;
            sine_reg0   <= 36'sb1101010110111111010100011000010111;
        end
        1124: begin
            cosine_reg0 <= 36'sb11101000100101010100110001111101010;
            sine_reg0   <= 36'sb1101010111101100111111010111010111;
        end
        1125: begin
            cosine_reg0 <= 36'sb11101000100010101100101100011001001;
            sine_reg0   <= 36'sb1101011000011010101001110101011000;
        end
        1126: begin
            cosine_reg0 <= 36'sb11101000100000000100011101110111011;
            sine_reg0   <= 36'sb1101011001001000010011110010010111;
        end
        1127: begin
            cosine_reg0 <= 36'sb11101000011101011100000110010111110;
            sine_reg0   <= 36'sb1101011001110101111101001110010011;
        end
        1128: begin
            cosine_reg0 <= 36'sb11101000011010110011100101111010110;
            sine_reg0   <= 36'sb1101011010100011100110001001001011;
        end
        1129: begin
            cosine_reg0 <= 36'sb11101000011000001010111100100000001;
            sine_reg0   <= 36'sb1101011011010001001110100010111101;
        end
        1130: begin
            cosine_reg0 <= 36'sb11101000010101100010001010001000001;
            sine_reg0   <= 36'sb1101011011111110110110011011100110;
        end
        1131: begin
            cosine_reg0 <= 36'sb11101000010010111001001110110011000;
            sine_reg0   <= 36'sb1101011100101100011101110011000101;
        end
        1132: begin
            cosine_reg0 <= 36'sb11101000010000010000001010100000101;
            sine_reg0   <= 36'sb1101011101011010000100101001011001;
        end
        1133: begin
            cosine_reg0 <= 36'sb11101000001101100110111101010001001;
            sine_reg0   <= 36'sb1101011110000111101010111110011111;
        end
        1134: begin
            cosine_reg0 <= 36'sb11101000001010111101100111000100110;
            sine_reg0   <= 36'sb1101011110110101010000110010010110;
        end
        1135: begin
            cosine_reg0 <= 36'sb11101000001000010100000111111011100;
            sine_reg0   <= 36'sb1101011111100010110110000100111100;
        end
        1136: begin
            cosine_reg0 <= 36'sb11101000000101101010011111110101100;
            sine_reg0   <= 36'sb1101100000010000011010110110001111;
        end
        1137: begin
            cosine_reg0 <= 36'sb11101000000011000000101110110010110;
            sine_reg0   <= 36'sb1101100000111101111111000110001110;
        end
        1138: begin
            cosine_reg0 <= 36'sb11101000000000010110110100110011101;
            sine_reg0   <= 36'sb1101100001101011100010110100110111;
        end
        1139: begin
            cosine_reg0 <= 36'sb11100111111101101100110001110111111;
            sine_reg0   <= 36'sb1101100010011001000110000010001000;
        end
        1140: begin
            cosine_reg0 <= 36'sb11100111111011000010100101111111111;
            sine_reg0   <= 36'sb1101100011000110101000101101111111;
        end
        1141: begin
            cosine_reg0 <= 36'sb11100111111000011000010001001011101;
            sine_reg0   <= 36'sb1101100011110100001010111000011010;
        end
        1142: begin
            cosine_reg0 <= 36'sb11100111110101101101110011011011001;
            sine_reg0   <= 36'sb1101100100100001101100100001011000;
        end
        1143: begin
            cosine_reg0 <= 36'sb11100111110011000011001100101110110;
            sine_reg0   <= 36'sb1101100101001111001101101000111000;
        end
        1144: begin
            cosine_reg0 <= 36'sb11100111110000011000011101000110011;
            sine_reg0   <= 36'sb1101100101111100101110001110110110;
        end
        1145: begin
            cosine_reg0 <= 36'sb11100111101101101101100100100010001;
            sine_reg0   <= 36'sb1101100110101010001110010011010010;
        end
        1146: begin
            cosine_reg0 <= 36'sb11100111101011000010100011000010001;
            sine_reg0   <= 36'sb1101100111010111101101110110001010;
        end
        1147: begin
            cosine_reg0 <= 36'sb11100111101000010111011000100110100;
            sine_reg0   <= 36'sb1101101000000101001100110111011011;
        end
        1148: begin
            cosine_reg0 <= 36'sb11100111100101101100000101001111100;
            sine_reg0   <= 36'sb1101101000110010101011010111000101;
        end
        1149: begin
            cosine_reg0 <= 36'sb11100111100011000000101000111100111;
            sine_reg0   <= 36'sb1101101001100000001001010101000101;
        end
        1150: begin
            cosine_reg0 <= 36'sb11100111100000010101000011101111000;
            sine_reg0   <= 36'sb1101101010001101100110110001011010;
        end
        1151: begin
            cosine_reg0 <= 36'sb11100111011101101001010101100110000;
            sine_reg0   <= 36'sb1101101010111011000011101100000011;
        end
        1152: begin
            cosine_reg0 <= 36'sb11100111011010111101011110100001110;
            sine_reg0   <= 36'sb1101101011101000100000000100111100;
        end
        1153: begin
            cosine_reg0 <= 36'sb11100111011000010001011110100010101;
            sine_reg0   <= 36'sb1101101100010101111011111100000100;
        end
        1154: begin
            cosine_reg0 <= 36'sb11100111010101100101010101101000100;
            sine_reg0   <= 36'sb1101101101000011010111010001011011;
        end
        1155: begin
            cosine_reg0 <= 36'sb11100111010010111001000011110011101;
            sine_reg0   <= 36'sb1101101101110000110010000100111101;
        end
        1156: begin
            cosine_reg0 <= 36'sb11100111010000001100101001000100000;
            sine_reg0   <= 36'sb1101101110011110001100010110101010;
        end
        1157: begin
            cosine_reg0 <= 36'sb11100111001101100000000101011001110;
            sine_reg0   <= 36'sb1101101111001011100110000110011111;
        end
        1158: begin
            cosine_reg0 <= 36'sb11100111001010110011011000110101001;
            sine_reg0   <= 36'sb1101101111111000111111010100011011;
        end
        1159: begin
            cosine_reg0 <= 36'sb11100111001000000110100011010110000;
            sine_reg0   <= 36'sb1101110000100110011000000000011011;
        end
        1160: begin
            cosine_reg0 <= 36'sb11100111000101011001100100111100110;
            sine_reg0   <= 36'sb1101110001010011110000001010011111;
        end
        1161: begin
            cosine_reg0 <= 36'sb11100111000010101100011101101001001;
            sine_reg0   <= 36'sb1101110010000001000111110010100101;
        end
        1162: begin
            cosine_reg0 <= 36'sb11100110111111111111001101011011100;
            sine_reg0   <= 36'sb1101110010101110011110111000101010;
        end
        1163: begin
            cosine_reg0 <= 36'sb11100110111101010001110100010100000;
            sine_reg0   <= 36'sb1101110011011011110101011100101101;
        end
        1164: begin
            cosine_reg0 <= 36'sb11100110111010100100010010010010100;
            sine_reg0   <= 36'sb1101110100001001001011011110101100;
        end
        1165: begin
            cosine_reg0 <= 36'sb11100110110111110110100111010111011;
            sine_reg0   <= 36'sb1101110100110110100000111110100110;
        end
        1166: begin
            cosine_reg0 <= 36'sb11100110110101001000110011100010100;
            sine_reg0   <= 36'sb1101110101100011110101111100011000;
        end
        1167: begin
            cosine_reg0 <= 36'sb11100110110010011010110110110100001;
            sine_reg0   <= 36'sb1101110110010001001010011000000010;
        end
        1168: begin
            cosine_reg0 <= 36'sb11100110101111101100110001001100010;
            sine_reg0   <= 36'sb1101110110111110011110010001100000;
        end
        1169: begin
            cosine_reg0 <= 36'sb11100110101100111110100010101011000;
            sine_reg0   <= 36'sb1101110111101011110001101000110010;
        end
        1170: begin
            cosine_reg0 <= 36'sb11100110101010010000001011010000101;
            sine_reg0   <= 36'sb1101111000011001000100011101110110;
        end
        1171: begin
            cosine_reg0 <= 36'sb11100110100111100001101010111101000;
            sine_reg0   <= 36'sb1101111001000110010110110000101010;
        end
        1172: begin
            cosine_reg0 <= 36'sb11100110100100110011000001110000100;
            sine_reg0   <= 36'sb1101111001110011101000100001001100;
        end
        1173: begin
            cosine_reg0 <= 36'sb11100110100010000100001111101011000;
            sine_reg0   <= 36'sb1101111010100000111001101111011010;
        end
        1174: begin
            cosine_reg0 <= 36'sb11100110011111010101010100101100101;
            sine_reg0   <= 36'sb1101111011001110001010011011010100;
        end
        1175: begin
            cosine_reg0 <= 36'sb11100110011100100110010000110101101;
            sine_reg0   <= 36'sb1101111011111011011010100100110110;
        end
        1176: begin
            cosine_reg0 <= 36'sb11100110011001110111000100000110000;
            sine_reg0   <= 36'sb1101111100101000101010001100000000;
        end
        1177: begin
            cosine_reg0 <= 36'sb11100110010111000111101110011101111;
            sine_reg0   <= 36'sb1101111101010101111001010000101111;
        end
        1178: begin
            cosine_reg0 <= 36'sb11100110010100011000001111111101010;
            sine_reg0   <= 36'sb1101111110000011000111110011000001;
        end
        1179: begin
            cosine_reg0 <= 36'sb11100110010001101000101000100100100;
            sine_reg0   <= 36'sb1101111110110000010101110010110110;
        end
        1180: begin
            cosine_reg0 <= 36'sb11100110001110111000111000010011100;
            sine_reg0   <= 36'sb1101111111011101100011010000001011;
        end
        1181: begin
            cosine_reg0 <= 36'sb11100110001100001000111111001010011;
            sine_reg0   <= 36'sb1110000000001010110000001010111111;
        end
        1182: begin
            cosine_reg0 <= 36'sb11100110001001011000111101001001011;
            sine_reg0   <= 36'sb1110000000110111111100100011001111;
        end
        1183: begin
            cosine_reg0 <= 36'sb11100110000110101000110010010000100;
            sine_reg0   <= 36'sb1110000001100101001000011000111011;
        end
        1184: begin
            cosine_reg0 <= 36'sb11100110000011111000011110011111110;
            sine_reg0   <= 36'sb1110000010010010010011101100000000;
        end
        1185: begin
            cosine_reg0 <= 36'sb11100110000001001000000001110111100;
            sine_reg0   <= 36'sb1110000010111111011110011100011100;
        end
        1186: begin
            cosine_reg0 <= 36'sb11100101111110010111011100010111101;
            sine_reg0   <= 36'sb1110000011101100101000101010001110;
        end
        1187: begin
            cosine_reg0 <= 36'sb11100101111011100110101110000000010;
            sine_reg0   <= 36'sb1110000100011001110010010101010101;
        end
        1188: begin
            cosine_reg0 <= 36'sb11100101111000110101110110110001101;
            sine_reg0   <= 36'sb1110000101000110111011011101101101;
        end
        1189: begin
            cosine_reg0 <= 36'sb11100101110110000100110110101011110;
            sine_reg0   <= 36'sb1110000101110100000100000011010110;
        end
        1190: begin
            cosine_reg0 <= 36'sb11100101110011010011101101101110111;
            sine_reg0   <= 36'sb1110000110100001001100000110001111;
        end
        1191: begin
            cosine_reg0 <= 36'sb11100101110000100010011011111010111;
            sine_reg0   <= 36'sb1110000111001110010011100110010100;
        end
        1192: begin
            cosine_reg0 <= 36'sb11100101101101110001000001001111111;
            sine_reg0   <= 36'sb1110000111111011011010100011100100;
        end
        1193: begin
            cosine_reg0 <= 36'sb11100101101010111111011101101110010;
            sine_reg0   <= 36'sb1110001000101000100000111101111111;
        end
        1194: begin
            cosine_reg0 <= 36'sb11100101101000001101110001010101111;
            sine_reg0   <= 36'sb1110001001010101100110110101100001;
        end
        1195: begin
            cosine_reg0 <= 36'sb11100101100101011011111100000110111;
            sine_reg0   <= 36'sb1110001010000010101100001010001001;
        end
        1196: begin
            cosine_reg0 <= 36'sb11100101100010101001111110000001011;
            sine_reg0   <= 36'sb1110001010101111110000111011110110;
        end
        1197: begin
            cosine_reg0 <= 36'sb11100101011111110111110111000101100;
            sine_reg0   <= 36'sb1110001011011100110101001010100101;
        end
        1198: begin
            cosine_reg0 <= 36'sb11100101011101000101100111010011100;
            sine_reg0   <= 36'sb1110001100001001111000110110010110;
        end
        1199: begin
            cosine_reg0 <= 36'sb11100101011010010011001110101011010;
            sine_reg0   <= 36'sb1110001100110110111011111111000101;
        end
        1200: begin
            cosine_reg0 <= 36'sb11100101010111100000101101001100111;
            sine_reg0   <= 36'sb1110001101100011111110100100110010;
        end
        1201: begin
            cosine_reg0 <= 36'sb11100101010100101110000010111000101;
            sine_reg0   <= 36'sb1110001110010001000000100111011011;
        end
        1202: begin
            cosine_reg0 <= 36'sb11100101010001111011001111101110101;
            sine_reg0   <= 36'sb1110001110111110000010000110111110;
        end
        1203: begin
            cosine_reg0 <= 36'sb11100101001111001000010011101110110;
            sine_reg0   <= 36'sb1110001111101011000011000011011001;
        end
        1204: begin
            cosine_reg0 <= 36'sb11100101001100010101001110111001011;
            sine_reg0   <= 36'sb1110010000011000000011011100101011;
        end
        1205: begin
            cosine_reg0 <= 36'sb11100101001001100010000001001110100;
            sine_reg0   <= 36'sb1110010001000101000011010010110001;
        end
        1206: begin
            cosine_reg0 <= 36'sb11100101000110101110101010101110001;
            sine_reg0   <= 36'sb1110010001110010000010100101101011;
        end
        1207: begin
            cosine_reg0 <= 36'sb11100101000011111011001011011000100;
            sine_reg0   <= 36'sb1110010010011111000001010101010110;
        end
        1208: begin
            cosine_reg0 <= 36'sb11100101000001000111100011001101110;
            sine_reg0   <= 36'sb1110010011001011111111100001110000;
        end
        1209: begin
            cosine_reg0 <= 36'sb11100100111110010011110010001101110;
            sine_reg0   <= 36'sb1110010011111000111101001010111001;
        end
        1210: begin
            cosine_reg0 <= 36'sb11100100111011011111111000011001000;
            sine_reg0   <= 36'sb1110010100100101111010010000101101;
        end
        1211: begin
            cosine_reg0 <= 36'sb11100100111000101011110101101111010;
            sine_reg0   <= 36'sb1110010101010010110110110011001100;
        end
        1212: begin
            cosine_reg0 <= 36'sb11100100110101110111101010010000110;
            sine_reg0   <= 36'sb1110010101111111110010110010010100;
        end
        1213: begin
            cosine_reg0 <= 36'sb11100100110011000011010101111101101;
            sine_reg0   <= 36'sb1110010110101100101110001110000010;
        end
        1214: begin
            cosine_reg0 <= 36'sb11100100110000001110111000110110000;
            sine_reg0   <= 36'sb1110010111011001101001000110010110;
        end
        1215: begin
            cosine_reg0 <= 36'sb11100100101101011010010010111001111;
            sine_reg0   <= 36'sb1110011000000110100011011011001101;
        end
        1216: begin
            cosine_reg0 <= 36'sb11100100101010100101100100001001100;
            sine_reg0   <= 36'sb1110011000110011011101001100100110;
        end
        1217: begin
            cosine_reg0 <= 36'sb11100100100111110000101100100100111;
            sine_reg0   <= 36'sb1110011001100000010110011010011111;
        end
        1218: begin
            cosine_reg0 <= 36'sb11100100100100111011101100001100010;
            sine_reg0   <= 36'sb1110011010001101001111000100110110;
        end
        1219: begin
            cosine_reg0 <= 36'sb11100100100010000110100010111111100;
            sine_reg0   <= 36'sb1110011010111010000111001011101010;
        end
        1220: begin
            cosine_reg0 <= 36'sb11100100011111010001010000111110111;
            sine_reg0   <= 36'sb1110011011100110111110101110111000;
        end
        1221: begin
            cosine_reg0 <= 36'sb11100100011100011011110110001010101;
            sine_reg0   <= 36'sb1110011100010011110101101110100000;
        end
        1222: begin
            cosine_reg0 <= 36'sb11100100011001100110010010100010100;
            sine_reg0   <= 36'sb1110011101000000101100001010011111;
        end
        1223: begin
            cosine_reg0 <= 36'sb11100100010110110000100110000111000;
            sine_reg0   <= 36'sb1110011101101101100010000010110011;
        end
        1224: begin
            cosine_reg0 <= 36'sb11100100010011111010110000111000000;
            sine_reg0   <= 36'sb1110011110011010010111010111011100;
        end
        1225: begin
            cosine_reg0 <= 36'sb11100100010001000100110010110101101;
            sine_reg0   <= 36'sb1110011111000111001100001000010110;
        end
        1226: begin
            cosine_reg0 <= 36'sb11100100001110001110101100000000000;
            sine_reg0   <= 36'sb1110011111110100000000010101100010;
        end
        1227: begin
            cosine_reg0 <= 36'sb11100100001011011000011100010111011;
            sine_reg0   <= 36'sb1110100000100000110011111110111011;
        end
        1228: begin
            cosine_reg0 <= 36'sb11100100001000100010000011111011101;
            sine_reg0   <= 36'sb1110100001001101100111000100100010;
        end
        1229: begin
            cosine_reg0 <= 36'sb11100100000101101011100010101101000;
            sine_reg0   <= 36'sb1110100001111010011001100110010100;
        end
        1230: begin
            cosine_reg0 <= 36'sb11100100000010110100111000101011101;
            sine_reg0   <= 36'sb1110100010100111001011100100010000;
        end
        1231: begin
            cosine_reg0 <= 36'sb11100011111111111110000101110111101;
            sine_reg0   <= 36'sb1110100011010011111100111110010011;
        end
        1232: begin
            cosine_reg0 <= 36'sb11100011111101000111001010010001000;
            sine_reg0   <= 36'sb1110100100000000101101110100011101;
        end
        1233: begin
            cosine_reg0 <= 36'sb11100011111010010000000101110111111;
            sine_reg0   <= 36'sb1110100100101101011110000110101011;
        end
        1234: begin
            cosine_reg0 <= 36'sb11100011110111011000111000101100100;
            sine_reg0   <= 36'sb1110100101011010001101110100111011;
        end
        1235: begin
            cosine_reg0 <= 36'sb11100011110100100001100010101110111;
            sine_reg0   <= 36'sb1110100110000110111100111111001100;
        end
        1236: begin
            cosine_reg0 <= 36'sb11100011110001101010000011111111000;
            sine_reg0   <= 36'sb1110100110110011101011100101011101;
        end
        1237: begin
            cosine_reg0 <= 36'sb11100011101110110010011100011101010;
            sine_reg0   <= 36'sb1110100111100000011001100111101011;
        end
        1238: begin
            cosine_reg0 <= 36'sb11100011101011111010101100001001100;
            sine_reg0   <= 36'sb1110101000001101000111000101110101;
        end
        1239: begin
            cosine_reg0 <= 36'sb11100011101001000010110011000100000;
            sine_reg0   <= 36'sb1110101000111001110011111111111001;
        end
        1240: begin
            cosine_reg0 <= 36'sb11100011100110001010110001001100111;
            sine_reg0   <= 36'sb1110101001100110100000010101110101;
        end
        1241: begin
            cosine_reg0 <= 36'sb11100011100011010010100110100100001;
            sine_reg0   <= 36'sb1110101010010011001100000111100111;
        end
        1242: begin
            cosine_reg0 <= 36'sb11100011100000011010010011001001111;
            sine_reg0   <= 36'sb1110101010111111110111010101001111;
        end
        1243: begin
            cosine_reg0 <= 36'sb11100011011101100001110110111110011;
            sine_reg0   <= 36'sb1110101011101100100001111110101001;
        end
        1244: begin
            cosine_reg0 <= 36'sb11100011011010101001010010000001100;
            sine_reg0   <= 36'sb1110101100011001001100000011110101;
        end
        1245: begin
            cosine_reg0 <= 36'sb11100011010111110000100100010011101;
            sine_reg0   <= 36'sb1110101101000101110101100100110001;
        end
        1246: begin
            cosine_reg0 <= 36'sb11100011010100110111101101110100101;
            sine_reg0   <= 36'sb1110101101110010011110100001011010;
        end
        1247: begin
            cosine_reg0 <= 36'sb11100011010001111110101110100100110;
            sine_reg0   <= 36'sb1110101110011111000110111001110000;
        end
        1248: begin
            cosine_reg0 <= 36'sb11100011001111000101100110100100001;
            sine_reg0   <= 36'sb1110101111001011101110101101110000;
        end
        1249: begin
            cosine_reg0 <= 36'sb11100011001100001100010101110010111;
            sine_reg0   <= 36'sb1110101111111000010101111101011001;
        end
        1250: begin
            cosine_reg0 <= 36'sb11100011001001010010111100010000111;
            sine_reg0   <= 36'sb1110110000100100111100101000101010;
        end
        1251: begin
            cosine_reg0 <= 36'sb11100011000110011001011001111110101;
            sine_reg0   <= 36'sb1110110001010001100010101111011111;
        end
        1252: begin
            cosine_reg0 <= 36'sb11100011000011011111101110111011111;
            sine_reg0   <= 36'sb1110110001111110001000010001111000;
        end
        1253: begin
            cosine_reg0 <= 36'sb11100011000000100101111011001001000;
            sine_reg0   <= 36'sb1110110010101010101101001111110011;
        end
        1254: begin
            cosine_reg0 <= 36'sb11100010111101101011111110100101111;
            sine_reg0   <= 36'sb1110110011010111010001101001001111;
        end
        1255: begin
            cosine_reg0 <= 36'sb11100010111010110001111001010010111;
            sine_reg0   <= 36'sb1110110100000011110101011110001000;
        end
        1256: begin
            cosine_reg0 <= 36'sb11100010110111110111101011001111111;
            sine_reg0   <= 36'sb1110110100110000011000101110011111;
        end
        1257: begin
            cosine_reg0 <= 36'sb11100010110100111101010100011101001;
            sine_reg0   <= 36'sb1110110101011100111011011010010000;
        end
        1258: begin
            cosine_reg0 <= 36'sb11100010110010000010110100111010101;
            sine_reg0   <= 36'sb1110110110001001011101100001011011;
        end
        1259: begin
            cosine_reg0 <= 36'sb11100010101111001000001100101000101;
            sine_reg0   <= 36'sb1110110110110101111111000011111110;
        end
        1260: begin
            cosine_reg0 <= 36'sb11100010101100001101011011100111010;
            sine_reg0   <= 36'sb1110110111100010100000000001110110;
        end
        1261: begin
            cosine_reg0 <= 36'sb11100010101001010010100001110110100;
            sine_reg0   <= 36'sb1110111000001111000000011011000010;
        end
        1262: begin
            cosine_reg0 <= 36'sb11100010100110010111011111010110100;
            sine_reg0   <= 36'sb1110111000111011100000001111100001;
        end
        1263: begin
            cosine_reg0 <= 36'sb11100010100011011100010100000111011;
            sine_reg0   <= 36'sb1110111001100111111111011111010001;
        end
        1264: begin
            cosine_reg0 <= 36'sb11100010100000100001000000001001010;
            sine_reg0   <= 36'sb1110111010010100011110001010010000;
        end
        1265: begin
            cosine_reg0 <= 36'sb11100010011101100101100011011100010;
            sine_reg0   <= 36'sb1110111011000000111100010000011100;
        end
        1266: begin
            cosine_reg0 <= 36'sb11100010011010101001111110000000100;
            sine_reg0   <= 36'sb1110111011101101011001110001110011;
        end
        1267: begin
            cosine_reg0 <= 36'sb11100010010111101110001111110110000;
            sine_reg0   <= 36'sb1110111100011001110110101110010101;
        end
        1268: begin
            cosine_reg0 <= 36'sb11100010010100110010011000111101001;
            sine_reg0   <= 36'sb1110111101000110010011000101111111;
        end
        1269: begin
            cosine_reg0 <= 36'sb11100010010001110110011001010101101;
            sine_reg0   <= 36'sb1110111101110010101110111000101111;
        end
        1270: begin
            cosine_reg0 <= 36'sb11100010001110111010010000111111111;
            sine_reg0   <= 36'sb1110111110011111001010000110100100;
        end
        1271: begin
            cosine_reg0 <= 36'sb11100010001011111101111111111100000;
            sine_reg0   <= 36'sb1110111111001011100100101111011011;
        end
        1272: begin
            cosine_reg0 <= 36'sb11100010001001000001100110001010000;
            sine_reg0   <= 36'sb1110111111110111111110110011010101;
        end
        1273: begin
            cosine_reg0 <= 36'sb11100010000110000101000011101001111;
            sine_reg0   <= 36'sb1111000000100100011000010010001110;
        end
        1274: begin
            cosine_reg0 <= 36'sb11100010000011001000011000011100000;
            sine_reg0   <= 36'sb1111000001010000110001001100000100;
        end
        1275: begin
            cosine_reg0 <= 36'sb11100010000000001011100100100000011;
            sine_reg0   <= 36'sb1111000001111101001001100000110111;
        end
        1276: begin
            cosine_reg0 <= 36'sb11100001111101001110100111110111001;
            sine_reg0   <= 36'sb1111000010101001100001010000100100;
        end
        1277: begin
            cosine_reg0 <= 36'sb11100001111010010001100010100000011;
            sine_reg0   <= 36'sb1111000011010101111000011011001011;
        end
        1278: begin
            cosine_reg0 <= 36'sb11100001110111010100010100011100001;
            sine_reg0   <= 36'sb1111000100000010001111000000101000;
        end
        1279: begin
            cosine_reg0 <= 36'sb11100001110100010110111101101010101;
            sine_reg0   <= 36'sb1111000100101110100101000000111010;
        end
        1280: begin
            cosine_reg0 <= 36'sb11100001110001011001011110001011111;
            sine_reg0   <= 36'sb1111000101011010111010011100000000;
        end
        1281: begin
            cosine_reg0 <= 36'sb11100001101110011011110110000000001;
            sine_reg0   <= 36'sb1111000110000111001111010001111000;
        end
        1282: begin
            cosine_reg0 <= 36'sb11100001101011011110000101000111011;
            sine_reg0   <= 36'sb1111000110110011100011100010100001;
        end
        1283: begin
            cosine_reg0 <= 36'sb11100001101000100000001011100001111;
            sine_reg0   <= 36'sb1111000111011111110111001101110111;
        end
        1284: begin
            cosine_reg0 <= 36'sb11100001100101100010001001001111101;
            sine_reg0   <= 36'sb1111001000001100001010010011111011;
        end
        1285: begin
            cosine_reg0 <= 36'sb11100001100010100011111110010000101;
            sine_reg0   <= 36'sb1111001000111000011100110100101010;
        end
        1286: begin
            cosine_reg0 <= 36'sb11100001011111100101101010100101010;
            sine_reg0   <= 36'sb1111001001100100101110110000000010;
        end
        1287: begin
            cosine_reg0 <= 36'sb11100001011100100111001110001101100;
            sine_reg0   <= 36'sb1111001010010001000000000110000001;
        end
        1288: begin
            cosine_reg0 <= 36'sb11100001011001101000101001001001100;
            sine_reg0   <= 36'sb1111001010111101010000110110100111;
        end
        1289: begin
            cosine_reg0 <= 36'sb11100001010110101001111011011001010;
            sine_reg0   <= 36'sb1111001011101001100001000001110001;
        end
        1290: begin
            cosine_reg0 <= 36'sb11100001010011101011000100111101000;
            sine_reg0   <= 36'sb1111001100010101110000100111011110;
        end
        1291: begin
            cosine_reg0 <= 36'sb11100001010000101100000101110100111;
            sine_reg0   <= 36'sb1111001101000001111111100111101011;
        end
        1292: begin
            cosine_reg0 <= 36'sb11100001001101101100111110000000111;
            sine_reg0   <= 36'sb1111001101101110001110000010010111;
        end
        1293: begin
            cosine_reg0 <= 36'sb11100001001010101101101101100001010;
            sine_reg0   <= 36'sb1111001110011010011011110111100001;
        end
        1294: begin
            cosine_reg0 <= 36'sb11100001000111101110010100010110000;
            sine_reg0   <= 36'sb1111001111000110101001000111000111;
        end
        1295: begin
            cosine_reg0 <= 36'sb11100001000100101110110010011111010;
            sine_reg0   <= 36'sb1111001111110010110101110001000111;
        end
        1296: begin
            cosine_reg0 <= 36'sb11100001000001101111000111111101001;
            sine_reg0   <= 36'sb1111010000011111000001110101011111;
        end
        1297: begin
            cosine_reg0 <= 36'sb11100000111110101111010100101111111;
            sine_reg0   <= 36'sb1111010001001011001101010100001101;
        end
        1298: begin
            cosine_reg0 <= 36'sb11100000111011101111011000110111100;
            sine_reg0   <= 36'sb1111010001110111011000001101010001;
        end
        1299: begin
            cosine_reg0 <= 36'sb11100000111000101111010100010100001;
            sine_reg0   <= 36'sb1111010010100011100010100000100111;
        end
        1300: begin
            cosine_reg0 <= 36'sb11100000110101101111000111000101110;
            sine_reg0   <= 36'sb1111010011001111101100001110010000;
        end
        1301: begin
            cosine_reg0 <= 36'sb11100000110010101110110001001100110;
            sine_reg0   <= 36'sb1111010011111011110101010110001000;
        end
        1302: begin
            cosine_reg0 <= 36'sb11100000101111101110010010101001000;
            sine_reg0   <= 36'sb1111010100100111111101111000001110;
        end
        1303: begin
            cosine_reg0 <= 36'sb11100000101100101101101011011010110;
            sine_reg0   <= 36'sb1111010101010100000101110100100001;
        end
        1304: begin
            cosine_reg0 <= 36'sb11100000101001101100111011100010001;
            sine_reg0   <= 36'sb1111010110000000001101001010111110;
        end
        1305: begin
            cosine_reg0 <= 36'sb11100000100110101100000010111111001;
            sine_reg0   <= 36'sb1111010110101100010011111011100100;
        end
        1306: begin
            cosine_reg0 <= 36'sb11100000100011101011000001110010000;
            sine_reg0   <= 36'sb1111010111011000011010000110010010;
        end
        1307: begin
            cosine_reg0 <= 36'sb11100000100000101001110111111010110;
            sine_reg0   <= 36'sb1111011000000100011111101011000101;
        end
        1308: begin
            cosine_reg0 <= 36'sb11100000011101101000100101011001100;
            sine_reg0   <= 36'sb1111011000110000100100101001111100;
        end
        1309: begin
            cosine_reg0 <= 36'sb11100000011010100111001010001110100;
            sine_reg0   <= 36'sb1111011001011100101001000010110101;
        end
        1310: begin
            cosine_reg0 <= 36'sb11100000010111100101100110011001110;
            sine_reg0   <= 36'sb1111011010001000101100110101101111;
        end
        1311: begin
            cosine_reg0 <= 36'sb11100000010100100011111001111011011;
            sine_reg0   <= 36'sb1111011010110100110000000010101000;
        end
        1312: begin
            cosine_reg0 <= 36'sb11100000010001100010000100110011100;
            sine_reg0   <= 36'sb1111011011100000110010101001011101;
        end
        1313: begin
            cosine_reg0 <= 36'sb11100000001110100000000111000010010;
            sine_reg0   <= 36'sb1111011100001100110100101010001111;
        end
        1314: begin
            cosine_reg0 <= 36'sb11100000001011011110000000100111110;
            sine_reg0   <= 36'sb1111011100111000110110000100111001;
        end
        1315: begin
            cosine_reg0 <= 36'sb11100000001000011011110001100100001;
            sine_reg0   <= 36'sb1111011101100100110110111001011100;
        end
        1316: begin
            cosine_reg0 <= 36'sb11100000000101011001011001110111100;
            sine_reg0   <= 36'sb1111011110010000110111000111110101;
        end
        1317: begin
            cosine_reg0 <= 36'sb11100000000010010110111001100001111;
            sine_reg0   <= 36'sb1111011110111100110110110000000011;
        end
        1318: begin
            cosine_reg0 <= 36'sb11011111111111010100010000100011100;
            sine_reg0   <= 36'sb1111011111101000110101110010000100;
        end
        1319: begin
            cosine_reg0 <= 36'sb11011111111100010001011110111100100;
            sine_reg0   <= 36'sb1111100000010100110100001101110110;
        end
        1320: begin
            cosine_reg0 <= 36'sb11011111111001001110100100101101000;
            sine_reg0   <= 36'sb1111100001000000110010000011011000;
        end
        1321: begin
            cosine_reg0 <= 36'sb11011111110110001011100001110100111;
            sine_reg0   <= 36'sb1111100001101100101111010010100111;
        end
        1322: begin
            cosine_reg0 <= 36'sb11011111110011001000010110010100101;
            sine_reg0   <= 36'sb1111100010011000101011111011100010;
        end
        1323: begin
            cosine_reg0 <= 36'sb11011111110000000101000010001100001;
            sine_reg0   <= 36'sb1111100011000100100111111110001000;
        end
        1324: begin
            cosine_reg0 <= 36'sb11011111101101000001100101011011100;
            sine_reg0   <= 36'sb1111100011110000100011011010010111;
        end
        1325: begin
            cosine_reg0 <= 36'sb11011111101001111110000000000010111;
            sine_reg0   <= 36'sb1111100100011100011110010000001101;
        end
        1326: begin
            cosine_reg0 <= 36'sb11011111100110111010010010000010011;
            sine_reg0   <= 36'sb1111100101001000011000011111101000;
        end
        1327: begin
            cosine_reg0 <= 36'sb11011111100011110110011011011010010;
            sine_reg0   <= 36'sb1111100101110100010010001000100111;
        end
        1328: begin
            cosine_reg0 <= 36'sb11011111100000110010011100001010100;
            sine_reg0   <= 36'sb1111100110100000001011001011000111;
        end
        1329: begin
            cosine_reg0 <= 36'sb11011111011101101110010100010011010;
            sine_reg0   <= 36'sb1111100111001100000011100111001001;
        end
        1330: begin
            cosine_reg0 <= 36'sb11011111011010101010000011110100101;
            sine_reg0   <= 36'sb1111100111110111111011011100101000;
        end
        1331: begin
            cosine_reg0 <= 36'sb11011111010111100101101010101110101;
            sine_reg0   <= 36'sb1111101000100011110010101011100101;
        end
        1332: begin
            cosine_reg0 <= 36'sb11011111010100100001001001000001101;
            sine_reg0   <= 36'sb1111101001001111101001010011111101;
        end
        1333: begin
            cosine_reg0 <= 36'sb11011111010001011100011110101101101;
            sine_reg0   <= 36'sb1111101001111011011111010101101110;
        end
        1334: begin
            cosine_reg0 <= 36'sb11011111001110010111101011110010101;
            sine_reg0   <= 36'sb1111101010100111010100110000110111;
        end
        1335: begin
            cosine_reg0 <= 36'sb11011111001011010010110000010000111;
            sine_reg0   <= 36'sb1111101011010011001001100101010111;
        end
        1336: begin
            cosine_reg0 <= 36'sb11011111001000001101101100001000011;
            sine_reg0   <= 36'sb1111101011111110111101110011001010;
        end
        1337: begin
            cosine_reg0 <= 36'sb11011111000101001000011111011001100;
            sine_reg0   <= 36'sb1111101100101010110001011010010001;
        end
        1338: begin
            cosine_reg0 <= 36'sb11011111000010000011001010000100001;
            sine_reg0   <= 36'sb1111101101010110100100011010101001;
        end
        1339: begin
            cosine_reg0 <= 36'sb11011110111110111101101100001000011;
            sine_reg0   <= 36'sb1111101110000010010110110100010000;
        end
        1340: begin
            cosine_reg0 <= 36'sb11011110111011111000000101100110100;
            sine_reg0   <= 36'sb1111101110101110001000100111000100;
        end
        1341: begin
            cosine_reg0 <= 36'sb11011110111000110010010110011110100;
            sine_reg0   <= 36'sb1111101111011001111001110011000101;
        end
        1342: begin
            cosine_reg0 <= 36'sb11011110110101101100011110110000101;
            sine_reg0   <= 36'sb1111110000000101101010011000010000;
        end
        1343: begin
            cosine_reg0 <= 36'sb11011110110010100110011110011100111;
            sine_reg0   <= 36'sb1111110000110001011010010110100100;
        end
        1344: begin
            cosine_reg0 <= 36'sb11011110101111100000010101100011011;
            sine_reg0   <= 36'sb1111110001011101001001101101111111;
        end
        1345: begin
            cosine_reg0 <= 36'sb11011110101100011010000100000100011;
            sine_reg0   <= 36'sb1111110010001000111000011110011111;
        end
        1346: begin
            cosine_reg0 <= 36'sb11011110101001010011101001111111110;
            sine_reg0   <= 36'sb1111110010110100100110101000000010;
        end
        1347: begin
            cosine_reg0 <= 36'sb11011110100110001101000111010101111;
            sine_reg0   <= 36'sb1111110011100000010100001010100111;
        end
        1348: begin
            cosine_reg0 <= 36'sb11011110100011000110011100000110110;
            sine_reg0   <= 36'sb1111110100001100000001000110001101;
        end
        1349: begin
            cosine_reg0 <= 36'sb11011110011111111111101000010010100;
            sine_reg0   <= 36'sb1111110100110111101101011010110001;
        end
        1350: begin
            cosine_reg0 <= 36'sb11011110011100111000101011111001010;
            sine_reg0   <= 36'sb1111110101100011011001001000010010;
        end
        1351: begin
            cosine_reg0 <= 36'sb11011110011001110001100110111011001;
            sine_reg0   <= 36'sb1111110110001111000100001110101110;
        end
        1352: begin
            cosine_reg0 <= 36'sb11011110010110101010011001011000010;
            sine_reg0   <= 36'sb1111110110111010101110101110000100;
        end
        1353: begin
            cosine_reg0 <= 36'sb11011110010011100011000011010000110;
            sine_reg0   <= 36'sb1111110111100110011000100110010010;
        end
        1354: begin
            cosine_reg0 <= 36'sb11011110010000011011100100100100110;
            sine_reg0   <= 36'sb1111111000010010000001110111010101;
        end
        1355: begin
            cosine_reg0 <= 36'sb11011110001101010011111101010100011;
            sine_reg0   <= 36'sb1111111000111101101010100001001101;
        end
        1356: begin
            cosine_reg0 <= 36'sb11011110001010001100001101011111101;
            sine_reg0   <= 36'sb1111111001101001010010100011111000;
        end
        1357: begin
            cosine_reg0 <= 36'sb11011110000111000100010101000110110;
            sine_reg0   <= 36'sb1111111010010100111001111111010100;
        end
        1358: begin
            cosine_reg0 <= 36'sb11011110000011111100010100001001111;
            sine_reg0   <= 36'sb1111111011000000100000110011011111;
        end
        1359: begin
            cosine_reg0 <= 36'sb11011110000000110100001010101001001;
            sine_reg0   <= 36'sb1111111011101100000111000000011000;
        end
        1360: begin
            cosine_reg0 <= 36'sb11011101111101101011111000100100100;
            sine_reg0   <= 36'sb1111111100010111101100100101111100;
        end
        1361: begin
            cosine_reg0 <= 36'sb11011101111010100011011101111100010;
            sine_reg0   <= 36'sb1111111101000011010001100100001100;
        end
        1362: begin
            cosine_reg0 <= 36'sb11011101110111011010111010110000011;
            sine_reg0   <= 36'sb1111111101101110110101111011000011;
        end
        1363: begin
            cosine_reg0 <= 36'sb11011101110100010010001111000001001;
            sine_reg0   <= 36'sb1111111110011010011001101010100010;
        end
        1364: begin
            cosine_reg0 <= 36'sb11011101110001001001011010101110101;
            sine_reg0   <= 36'sb1111111111000101111100110010100110;
        end
        1365: begin
            cosine_reg0 <= 36'sb11011101101110000000011101111000111;
            sine_reg0   <= 36'sb1111111111110001011111010011001110;
        end
        1366: begin
            cosine_reg0 <= 36'sb11011101101010110111011000100000000;
            sine_reg0   <= 36'sb10000000000011101000001001100011000;
        end
        1367: begin
            cosine_reg0 <= 36'sb11011101100111101110001010100100010;
            sine_reg0   <= 36'sb10000000001001000100010011110000010;
        end
        1368: begin
            cosine_reg0 <= 36'sb11011101100100100100110100000101101;
            sine_reg0   <= 36'sb10000000001110100000011001000001010;
        end
        1369: begin
            cosine_reg0 <= 36'sb11011101100001011011010101000100010;
            sine_reg0   <= 36'sb10000000010011111100011001010110000;
        end
        1370: begin
            cosine_reg0 <= 36'sb11011101011110010001101101100000011;
            sine_reg0   <= 36'sb10000000011001011000010100101110001;
        end
        1371: begin
            cosine_reg0 <= 36'sb11011101011011000111111101011010000;
            sine_reg0   <= 36'sb10000000011110110100001011001001011;
        end
        1372: begin
            cosine_reg0 <= 36'sb11011101010111111110000100110001011;
            sine_reg0   <= 36'sb10000000100100001111111100100111101;
        end
        1373: begin
            cosine_reg0 <= 36'sb11011101010100110100000011100110011;
            sine_reg0   <= 36'sb10000000101001101011101001001000101;
        end
        1374: begin
            cosine_reg0 <= 36'sb11011101010001101001111001111001011;
            sine_reg0   <= 36'sb10000000101111000111010000101100010;
        end
        1375: begin
            cosine_reg0 <= 36'sb11011101001110011111100111101010011;
            sine_reg0   <= 36'sb10000000110100100010110011010010010;
        end
        1376: begin
            cosine_reg0 <= 36'sb11011101001011010101001100111001101;
            sine_reg0   <= 36'sb10000000111001111110010000111010011;
        end
        1377: begin
            cosine_reg0 <= 36'sb11011101001000001010101001100111000;
            sine_reg0   <= 36'sb10000000111111011001101001100100011;
        end
        1378: begin
            cosine_reg0 <= 36'sb11011101000100111111111101110010110;
            sine_reg0   <= 36'sb10000001000100110100111101010000001;
        end
        1379: begin
            cosine_reg0 <= 36'sb11011101000001110101001001011101001;
            sine_reg0   <= 36'sb10000001001010010000001011111101011;
        end
        1380: begin
            cosine_reg0 <= 36'sb11011100111110101010001100100110001;
            sine_reg0   <= 36'sb10000001001111101011010101101100000;
        end
        1381: begin
            cosine_reg0 <= 36'sb11011100111011011111000111001101110;
            sine_reg0   <= 36'sb10000001010101000110011010011011110;
        end
        1382: begin
            cosine_reg0 <= 36'sb11011100111000010011111001010100011;
            sine_reg0   <= 36'sb10000001011010100001011010001100011;
        end
        1383: begin
            cosine_reg0 <= 36'sb11011100110101001000100010111010000;
            sine_reg0   <= 36'sb10000001011111111100010100111101101;
        end
        1384: begin
            cosine_reg0 <= 36'sb11011100110001111101000011111110101;
            sine_reg0   <= 36'sb10000001100101010111001010101111011;
        end
        1385: begin
            cosine_reg0 <= 36'sb11011100101110110001011100100010101;
            sine_reg0   <= 36'sb10000001101010110001111011100001011;
        end
        1386: begin
            cosine_reg0 <= 36'sb11011100101011100101101100100110000;
            sine_reg0   <= 36'sb10000001110000001100100111010011100;
        end
        1387: begin
            cosine_reg0 <= 36'sb11011100101000011001110100001000110;
            sine_reg0   <= 36'sb10000001110101100111001110000101011;
        end
        1388: begin
            cosine_reg0 <= 36'sb11011100100101001101110011001011010;
            sine_reg0   <= 36'sb10000001111011000001101111110110111;
        end
        1389: begin
            cosine_reg0 <= 36'sb11011100100010000001101001101101011;
            sine_reg0   <= 36'sb10000010000000011100001100100111111;
        end
        1390: begin
            cosine_reg0 <= 36'sb11011100011110110101010111101111011;
            sine_reg0   <= 36'sb10000010000101110110100100011000001;
        end
        1391: begin
            cosine_reg0 <= 36'sb11011100011011101000111101010001011;
            sine_reg0   <= 36'sb10000010001011010000110111000111011;
        end
        1392: begin
            cosine_reg0 <= 36'sb11011100011000011100011010010011100;
            sine_reg0   <= 36'sb10000010010000101011000100110101011;
        end
        1393: begin
            cosine_reg0 <= 36'sb11011100010101001111101110110101111;
            sine_reg0   <= 36'sb10000010010110000101001101100010000;
        end
        1394: begin
            cosine_reg0 <= 36'sb11011100010010000010111010111000101;
            sine_reg0   <= 36'sb10000010011011011111010001001101000;
        end
        1395: begin
            cosine_reg0 <= 36'sb11011100001110110101111110011011110;
            sine_reg0   <= 36'sb10000010100000111001001111110110010;
        end
        1396: begin
            cosine_reg0 <= 36'sb11011100001011101000111001011111100;
            sine_reg0   <= 36'sb10000010100110010011001001011101011;
        end
        1397: begin
            cosine_reg0 <= 36'sb11011100001000011011101100000100000;
            sine_reg0   <= 36'sb10000010101011101100111110000010010;
        end
        1398: begin
            cosine_reg0 <= 36'sb11011100000101001110010110001001011;
            sine_reg0   <= 36'sb10000010110001000110101101100100110;
        end
        1399: begin
            cosine_reg0 <= 36'sb11011100000010000000110111101111110;
            sine_reg0   <= 36'sb10000010110110100000011000000100100;
        end
        1400: begin
            cosine_reg0 <= 36'sb11011011111110110011010000110111001;
            sine_reg0   <= 36'sb10000010111011111001111101100001100;
        end
        1401: begin
            cosine_reg0 <= 36'sb11011011111011100101100001011111110;
            sine_reg0   <= 36'sb10000011000001010011011101111011011;
        end
        1402: begin
            cosine_reg0 <= 36'sb11011011111000010111101001101001110;
            sine_reg0   <= 36'sb10000011000110101100111001010010000;
        end
        1403: begin
            cosine_reg0 <= 36'sb11011011110101001001101001010101001;
            sine_reg0   <= 36'sb10000011001100000110001111100101001;
        end
        1404: begin
            cosine_reg0 <= 36'sb11011011110001111011100000100010010;
            sine_reg0   <= 36'sb10000011010001011111100000110100100;
        end
        1405: begin
            cosine_reg0 <= 36'sb11011011101110101101001111010000111;
            sine_reg0   <= 36'sb10000011010110111000101101000000000;
        end
        1406: begin
            cosine_reg0 <= 36'sb11011011101011011110110101100001100;
            sine_reg0   <= 36'sb10000011011100010001110100000111011;
        end
        1407: begin
            cosine_reg0 <= 36'sb11011011101000010000010011010100000;
            sine_reg0   <= 36'sb10000011100001101010110110001010100;
        end
        1408: begin
            cosine_reg0 <= 36'sb11011011100101000001101000101000101;
            sine_reg0   <= 36'sb10000011100111000011110011001001000;
        end
        1409: begin
            cosine_reg0 <= 36'sb11011011100001110010110101011111100;
            sine_reg0   <= 36'sb10000011101100011100101011000010111;
        end
        1410: begin
            cosine_reg0 <= 36'sb11011011011110100011111001111000110;
            sine_reg0   <= 36'sb10000011110001110101011101110111110;
        end
        1411: begin
            cosine_reg0 <= 36'sb11011011011011010100110101110100011;
            sine_reg0   <= 36'sb10000011110111001110001011100111100;
        end
        1412: begin
            cosine_reg0 <= 36'sb11011011011000000101101001010010101;
            sine_reg0   <= 36'sb10000011111100100110110100010001110;
        end
        1413: begin
            cosine_reg0 <= 36'sb11011011010100110110010100010011100;
            sine_reg0   <= 36'sb10000100000001111111010111110110101;
        end
        1414: begin
            cosine_reg0 <= 36'sb11011011010001100110110110110111010;
            sine_reg0   <= 36'sb10000100000111010111110110010101101;
        end
        1415: begin
            cosine_reg0 <= 36'sb11011011001110010111010000111110000;
            sine_reg0   <= 36'sb10000100001100110000001111101110101;
        end
        1416: begin
            cosine_reg0 <= 36'sb11011011001011000111100010100111111;
            sine_reg0   <= 36'sb10000100010010001000100100000001100;
        end
        1417: begin
            cosine_reg0 <= 36'sb11011011000111110111101011110100111;
            sine_reg0   <= 36'sb10000100010111100000110011001110000;
        end
        1418: begin
            cosine_reg0 <= 36'sb11011011000100100111101100100101010;
            sine_reg0   <= 36'sb10000100011100111000111101010011111;
        end
        1419: begin
            cosine_reg0 <= 36'sb11011011000001010111100100111001000;
            sine_reg0   <= 36'sb10000100100010010001000010010010111;
        end
        1420: begin
            cosine_reg0 <= 36'sb11011010111110000111010100110000100;
            sine_reg0   <= 36'sb10000100100111101001000010001010111;
        end
        1421: begin
            cosine_reg0 <= 36'sb11011010111010110110111100001011101;
            sine_reg0   <= 36'sb10000100101101000000111100111011110;
        end
        1422: begin
            cosine_reg0 <= 36'sb11011010110111100110011011001010100;
            sine_reg0   <= 36'sb10000100110010011000110010100101001;
        end
        1423: begin
            cosine_reg0 <= 36'sb11011010110100010101110001101101100;
            sine_reg0   <= 36'sb10000100110111110000100011000110110;
        end
        1424: begin
            cosine_reg0 <= 36'sb11011010110001000100111111110100100;
            sine_reg0   <= 36'sb10000100111101001000001110100000101;
        end
        1425: begin
            cosine_reg0 <= 36'sb11011010101101110100000101011111101;
            sine_reg0   <= 36'sb10000101000010011111110100110010100;
        end
        1426: begin
            cosine_reg0 <= 36'sb11011010101010100011000010101111010;
            sine_reg0   <= 36'sb10000101000111110111010101111100001;
        end
        1427: begin
            cosine_reg0 <= 36'sb11011010100111010001110111100011010;
            sine_reg0   <= 36'sb10000101001101001110110001111101001;
        end
        1428: begin
            cosine_reg0 <= 36'sb11011010100100000000100011111011111;
            sine_reg0   <= 36'sb10000101010010100110001000110101101;
        end
        1429: begin
            cosine_reg0 <= 36'sb11011010100000101111000111111001010;
            sine_reg0   <= 36'sb10000101010111111101011010100101001;
        end
        1430: begin
            cosine_reg0 <= 36'sb11011010011101011101100011011011011;
            sine_reg0   <= 36'sb10000101011101010100100111001011101;
        end
        1431: begin
            cosine_reg0 <= 36'sb11011010011010001011110110100010101;
            sine_reg0   <= 36'sb10000101100010101011101110101000110;
        end
        1432: begin
            cosine_reg0 <= 36'sb11011010010110111010000001001110111;
            sine_reg0   <= 36'sb10000101101000000010110000111100011;
        end
        1433: begin
            cosine_reg0 <= 36'sb11011010010011101000000011100000011;
            sine_reg0   <= 36'sb10000101101101011001101110000110011;
        end
        1434: begin
            cosine_reg0 <= 36'sb11011010010000010101111101010111001;
            sine_reg0   <= 36'sb10000101110010110000100110000110011;
        end
        1435: begin
            cosine_reg0 <= 36'sb11011010001101000011101110110011100;
            sine_reg0   <= 36'sb10000101111000000111011000111100011;
        end
        1436: begin
            cosine_reg0 <= 36'sb11011010001001110001010111110101011;
            sine_reg0   <= 36'sb10000101111101011110000110100111111;
        end
        1437: begin
            cosine_reg0 <= 36'sb11011010000110011110111000011101000;
            sine_reg0   <= 36'sb10000110000010110100101111001001000;
        end
        1438: begin
            cosine_reg0 <= 36'sb11011010000011001100010000101010100;
            sine_reg0   <= 36'sb10000110001000001011010010011111010;
        end
        1439: begin
            cosine_reg0 <= 36'sb11011001111111111001100000011110000;
            sine_reg0   <= 36'sb10000110001101100001110000101010101;
        end
        1440: begin
            cosine_reg0 <= 36'sb11011001111100100110100111110111100;
            sine_reg0   <= 36'sb10000110010010111000001001101010111;
        end
        1441: begin
            cosine_reg0 <= 36'sb11011001111001010011100110110111011;
            sine_reg0   <= 36'sb10000110011000001110011101011111110;
        end
        1442: begin
            cosine_reg0 <= 36'sb11011001110110000000011101011101101;
            sine_reg0   <= 36'sb10000110011101100100101100001001000;
        end
        1443: begin
            cosine_reg0 <= 36'sb11011001110010101101001011101010010;
            sine_reg0   <= 36'sb10000110100010111010110101100110100;
        end
        1444: begin
            cosine_reg0 <= 36'sb11011001101111011001110001011101100;
            sine_reg0   <= 36'sb10000110101000010000111001111000000;
        end
        1445: begin
            cosine_reg0 <= 36'sb11011001101100000110001110110111101;
            sine_reg0   <= 36'sb10000110101101100110111000111101011;
        end
        1446: begin
            cosine_reg0 <= 36'sb11011001101000110010100011111000100;
            sine_reg0   <= 36'sb10000110110010111100110010110110011;
        end
        1447: begin
            cosine_reg0 <= 36'sb11011001100101011110110000100000100;
            sine_reg0   <= 36'sb10000110111000010010100111100010110;
        end
        1448: begin
            cosine_reg0 <= 36'sb11011001100010001010110100101111100;
            sine_reg0   <= 36'sb10000110111101101000010111000010010;
        end
        1449: begin
            cosine_reg0 <= 36'sb11011001011110110110110000100101110;
            sine_reg0   <= 36'sb10000111000010111110000001010100111;
        end
        1450: begin
            cosine_reg0 <= 36'sb11011001011011100010100100000011100;
            sine_reg0   <= 36'sb10000111001000010011100110011010010;
        end
        1451: begin
            cosine_reg0 <= 36'sb11011001011000001110001111001000110;
            sine_reg0   <= 36'sb10000111001101101001000110010010001;
        end
        1452: begin
            cosine_reg0 <= 36'sb11011001010100111001110001110101100;
            sine_reg0   <= 36'sb10000111010010111110100000111100011;
        end
        1453: begin
            cosine_reg0 <= 36'sb11011001010001100101001100001010001;
            sine_reg0   <= 36'sb10000111011000010011110110011000111;
        end
        1454: begin
            cosine_reg0 <= 36'sb11011001001110010000011110000110101;
            sine_reg0   <= 36'sb10000111011101101001000110100111011;
        end
        1455: begin
            cosine_reg0 <= 36'sb11011001001010111011100111101011010;
            sine_reg0   <= 36'sb10000111100010111110010001100111100;
        end
        1456: begin
            cosine_reg0 <= 36'sb11011001000111100110101000110111111;
            sine_reg0   <= 36'sb10000111101000010011010111011001010;
        end
        1457: begin
            cosine_reg0 <= 36'sb11011001000100010001100001101100111;
            sine_reg0   <= 36'sb10000111101101101000010111111100011;
        end
        1458: begin
            cosine_reg0 <= 36'sb11011001000000111100010010001010010;
            sine_reg0   <= 36'sb10000111110010111101010011010000101;
        end
        1459: begin
            cosine_reg0 <= 36'sb11011000111101100110111010010000001;
            sine_reg0   <= 36'sb10000111111000010010001001010101110;
        end
        1460: begin
            cosine_reg0 <= 36'sb11011000111010010001011001111110110;
            sine_reg0   <= 36'sb10000111111101100110111010001011101;
        end
        1461: begin
            cosine_reg0 <= 36'sb11011000110110111011110001010110001;
            sine_reg0   <= 36'sb10001000000010111011100101110010001;
        end
        1462: begin
            cosine_reg0 <= 36'sb11011000110011100110000000010110011;
            sine_reg0   <= 36'sb10001000001000010000001100001000111;
        end
        1463: begin
            cosine_reg0 <= 36'sb11011000110000010000000110111111110;
            sine_reg0   <= 36'sb10001000001101100100101101001111101;
        end
        1464: begin
            cosine_reg0 <= 36'sb11011000101100111010000101010010010;
            sine_reg0   <= 36'sb10001000010010111001001001000110100;
        end
        1465: begin
            cosine_reg0 <= 36'sb11011000101001100011111011001110001;
            sine_reg0   <= 36'sb10001000011000001101011111101100111;
        end
        1466: begin
            cosine_reg0 <= 36'sb11011000100110001101101000110011011;
            sine_reg0   <= 36'sb10001000011101100001110001000010111;
        end
        1467: begin
            cosine_reg0 <= 36'sb11011000100010110111001110000010010;
            sine_reg0   <= 36'sb10001000100010110101111101001000001;
        end
        1468: begin
            cosine_reg0 <= 36'sb11011000011111100000101010111010110;
            sine_reg0   <= 36'sb10001000101000001010000011111100100;
        end
        1469: begin
            cosine_reg0 <= 36'sb11011000011100001001111111011101001;
            sine_reg0   <= 36'sb10001000101101011110000101011111110;
        end
        1470: begin
            cosine_reg0 <= 36'sb11011000011000110011001011101001100;
            sine_reg0   <= 36'sb10001000110010110010000001110001110;
        end
        1471: begin
            cosine_reg0 <= 36'sb11011000010101011100001111011111111;
            sine_reg0   <= 36'sb10001000111000000101111000110010001;
        end
        1472: begin
            cosine_reg0 <= 36'sb11011000010010000101001011000000100;
            sine_reg0   <= 36'sb10001000111101011001101010100000110;
        end
        1473: begin
            cosine_reg0 <= 36'sb11011000001110101101111110001011100;
            sine_reg0   <= 36'sb10001001000010101101010110111101100;
        end
        1474: begin
            cosine_reg0 <= 36'sb11011000001011010110101001000001000;
            sine_reg0   <= 36'sb10001001001000000000111110001000001;
        end
        1475: begin
            cosine_reg0 <= 36'sb11011000000111111111001011100001000;
            sine_reg0   <= 36'sb10001001001101010100100000000000011;
        end
        1476: begin
            cosine_reg0 <= 36'sb11011000000100100111100101101011110;
            sine_reg0   <= 36'sb10001001010010100111111100100110001;
        end
        1477: begin
            cosine_reg0 <= 36'sb11011000000001001111110111100001100;
            sine_reg0   <= 36'sb10001001010111111011010011111001000;
        end
        1478: begin
            cosine_reg0 <= 36'sb11010111111101111000000001000010001;
            sine_reg0   <= 36'sb10001001011101001110100101111001000;
        end
        1479: begin
            cosine_reg0 <= 36'sb11010111111010100000000010001101111;
            sine_reg0   <= 36'sb10001001100010100001110010100101111;
        end
        1480: begin
            cosine_reg0 <= 36'sb11010111110111000111111011000100111;
            sine_reg0   <= 36'sb10001001100111110100111001111111011;
        end
        1481: begin
            cosine_reg0 <= 36'sb11010111110011101111101011100111010;
            sine_reg0   <= 36'sb10001001101101000111111100000101010;
        end
        1482: begin
            cosine_reg0 <= 36'sb11010111110000010111010011110101010;
            sine_reg0   <= 36'sb10001001110010011010111000110111011;
        end
        1483: begin
            cosine_reg0 <= 36'sb11010111101100111110110011101110110;
            sine_reg0   <= 36'sb10001001110111101101110000010101101;
        end
        1484: begin
            cosine_reg0 <= 36'sb11010111101001100110001011010100001;
            sine_reg0   <= 36'sb10001001111101000000100010011111100;
        end
        1485: begin
            cosine_reg0 <= 36'sb11010111100110001101011010100101011;
            sine_reg0   <= 36'sb10001010000010010011001111010101001;
        end
        1486: begin
            cosine_reg0 <= 36'sb11010111100010110100100001100010101;
            sine_reg0   <= 36'sb10001010000111100101110110110110001;
        end
        1487: begin
            cosine_reg0 <= 36'sb11010111011111011011100000001100000;
            sine_reg0   <= 36'sb10001010001100111000011001000010011;
        end
        1488: begin
            cosine_reg0 <= 36'sb11010111011100000010010110100001110;
            sine_reg0   <= 36'sb10001010010010001010110101111001100;
        end
        1489: begin
            cosine_reg0 <= 36'sb11010111011000101001000100100100000;
            sine_reg0   <= 36'sb10001010010111011101001101011011100;
        end
        1490: begin
            cosine_reg0 <= 36'sb11010111010101001111101010010010101;
            sine_reg0   <= 36'sb10001010011100101111011111101000001;
        end
        1491: begin
            cosine_reg0 <= 36'sb11010111010001110110000111101110001;
            sine_reg0   <= 36'sb10001010100010000001101100011111001;
        end
        1492: begin
            cosine_reg0 <= 36'sb11010111001110011100011100110110010;
            sine_reg0   <= 36'sb10001010100111010011110100000000010;
        end
        1493: begin
            cosine_reg0 <= 36'sb11010111001011000010101001101011100;
            sine_reg0   <= 36'sb10001010101100100101110110001011100;
        end
        1494: begin
            cosine_reg0 <= 36'sb11010111000111101000101110001101110;
            sine_reg0   <= 36'sb10001010110001110111110011000000011;
        end
        1495: begin
            cosine_reg0 <= 36'sb11010111000100001110101010011101010;
            sine_reg0   <= 36'sb10001010110111001001101010011110111;
        end
        1496: begin
            cosine_reg0 <= 36'sb11010111000000110100011110011010001;
            sine_reg0   <= 36'sb10001010111100011011011100100110110;
        end
        1497: begin
            cosine_reg0 <= 36'sb11010110111101011010001010000100011;
            sine_reg0   <= 36'sb10001011000001101101001001010111111;
        end
        1498: begin
            cosine_reg0 <= 36'sb11010110111001111111101101011100010;
            sine_reg0   <= 36'sb10001011000110111110110000110001111;
        end
        1499: begin
            cosine_reg0 <= 36'sb11010110110110100101001000100010000;
            sine_reg0   <= 36'sb10001011001100010000010010110100101;
        end
        1500: begin
            cosine_reg0 <= 36'sb11010110110011001010011011010101100;
            sine_reg0   <= 36'sb10001011010001100001101111100000000;
        end
        1501: begin
            cosine_reg0 <= 36'sb11010110101111101111100101110111000;
            sine_reg0   <= 36'sb10001011010110110011000110110011110;
        end
        1502: begin
            cosine_reg0 <= 36'sb11010110101100010100101000000110101;
            sine_reg0   <= 36'sb10001011011100000100011000101111100;
        end
        1503: begin
            cosine_reg0 <= 36'sb11010110101000111001100010000100101;
            sine_reg0   <= 36'sb10001011100001010101100101010011011;
        end
        1504: begin
            cosine_reg0 <= 36'sb11010110100101011110010011110001000;
            sine_reg0   <= 36'sb10001011100110100110101100011110111;
        end
        1505: begin
            cosine_reg0 <= 36'sb11010110100010000010111101001011111;
            sine_reg0   <= 36'sb10001011101011110111101110010010000;
        end
        1506: begin
            cosine_reg0 <= 36'sb11010110011110100111011110010101011;
            sine_reg0   <= 36'sb10001011110001001000101010101100011;
        end
        1507: begin
            cosine_reg0 <= 36'sb11010110011011001011110111001101101;
            sine_reg0   <= 36'sb10001011110110011001100001101110000;
        end
        1508: begin
            cosine_reg0 <= 36'sb11010110010111110000000111110100111;
            sine_reg0   <= 36'sb10001011111011101010010011010110100;
        end
        1509: begin
            cosine_reg0 <= 36'sb11010110010100010100010000001011010;
            sine_reg0   <= 36'sb10001100000000111010111111100101110;
        end
        1510: begin
            cosine_reg0 <= 36'sb11010110010000111000010000010000110;
            sine_reg0   <= 36'sb10001100000110001011100110011011100;
        end
        1511: begin
            cosine_reg0 <= 36'sb11010110001101011100001000000101101;
            sine_reg0   <= 36'sb10001100001011011100000111110111100;
        end
        1512: begin
            cosine_reg0 <= 36'sb11010110001001111111110111101001111;
            sine_reg0   <= 36'sb10001100010000101100100011111001110;
        end
        1513: begin
            cosine_reg0 <= 36'sb11010110000110100011011110111101110;
            sine_reg0   <= 36'sb10001100010101111100111010100001111;
        end
        1514: begin
            cosine_reg0 <= 36'sb11010110000011000110111110000001011;
            sine_reg0   <= 36'sb10001100011011001101001011101111110;
        end
        1515: begin
            cosine_reg0 <= 36'sb11010101111111101010010100110100110;
            sine_reg0   <= 36'sb10001100100000011101010111100011001;
        end
        1516: begin
            cosine_reg0 <= 36'sb11010101111100001101100011011000010;
            sine_reg0   <= 36'sb10001100100101101101011101111011110;
        end
        1517: begin
            cosine_reg0 <= 36'sb11010101111000110000101001101011111;
            sine_reg0   <= 36'sb10001100101010111101011110111001100;
        end
        1518: begin
            cosine_reg0 <= 36'sb11010101110101010011100111101111101;
            sine_reg0   <= 36'sb10001100110000001101011010011100010;
        end
        1519: begin
            cosine_reg0 <= 36'sb11010101110001110110011101100011111;
            sine_reg0   <= 36'sb10001100110101011101010000100011101;
        end
        1520: begin
            cosine_reg0 <= 36'sb11010101101110011001001011001000101;
            sine_reg0   <= 36'sb10001100111010101101000001001111100;
        end
        1521: begin
            cosine_reg0 <= 36'sb11010101101010111011110000011110000;
            sine_reg0   <= 36'sb10001100111111111100101100011111110;
        end
        1522: begin
            cosine_reg0 <= 36'sb11010101100111011110001101100100001;
            sine_reg0   <= 36'sb10001101000101001100010010010100000;
        end
        1523: begin
            cosine_reg0 <= 36'sb11010101100100000000100010011011010;
            sine_reg0   <= 36'sb10001101001010011011110010101100010;
        end
        1524: begin
            cosine_reg0 <= 36'sb11010101100000100010101111000011100;
            sine_reg0   <= 36'sb10001101001111101011001101101000001;
        end
        1525: begin
            cosine_reg0 <= 36'sb11010101011101000100110011011100110;
            sine_reg0   <= 36'sb10001101010100111010100011000111100;
        end
        1526: begin
            cosine_reg0 <= 36'sb11010101011001100110101111100111100;
            sine_reg0   <= 36'sb10001101011010001001110011001010001;
        end
        1527: begin
            cosine_reg0 <= 36'sb11010101010110001000100011100011101;
            sine_reg0   <= 36'sb10001101011111011000111101101111111;
        end
        1528: begin
            cosine_reg0 <= 36'sb11010101010010101010001111010001010;
            sine_reg0   <= 36'sb10001101100100101000000010111000100;
        end
        1529: begin
            cosine_reg0 <= 36'sb11010101001111001011110010110000110;
            sine_reg0   <= 36'sb10001101101001110111000010100011111;
        end
        1530: begin
            cosine_reg0 <= 36'sb11010101001011101101001110000010000;
            sine_reg0   <= 36'sb10001101101111000101111100110001101;
        end
        1531: begin
            cosine_reg0 <= 36'sb11010101001000001110100001000101011;
            sine_reg0   <= 36'sb10001101110100010100110001100001110;
        end
        1532: begin
            cosine_reg0 <= 36'sb11010101000100101111101011111010110;
            sine_reg0   <= 36'sb10001101111001100011100000110100000;
        end
        1533: begin
            cosine_reg0 <= 36'sb11010101000001010000101110100010011;
            sine_reg0   <= 36'sb10001101111110110010001010101000000;
        end
        1534: begin
            cosine_reg0 <= 36'sb11010100111101110001101000111100100;
            sine_reg0   <= 36'sb10001110000100000000101110111101110;
        end
        1535: begin
            cosine_reg0 <= 36'sb11010100111010010010011011001001001;
            sine_reg0   <= 36'sb10001110001001001111001101110100111;
        end
        1536: begin
            cosine_reg0 <= 36'sb11010100110110110011000101001000011;
            sine_reg0   <= 36'sb10001110001110011101100111001101011;
        end
        1537: begin
            cosine_reg0 <= 36'sb11010100110011010011100110111010011;
            sine_reg0   <= 36'sb10001110010011101011111011000110111;
        end
        1538: begin
            cosine_reg0 <= 36'sb11010100101111110100000000011111011;
            sine_reg0   <= 36'sb10001110011000111010001001100001011;
        end
        1539: begin
            cosine_reg0 <= 36'sb11010100101100010100010001110111100;
            sine_reg0   <= 36'sb10001110011110001000010010011100011;
        end
        1540: begin
            cosine_reg0 <= 36'sb11010100101000110100011011000010110;
            sine_reg0   <= 36'sb10001110100011010110010101111000000;
        end
        1541: begin
            cosine_reg0 <= 36'sb11010100100101010100011100000001011;
            sine_reg0   <= 36'sb10001110101000100100010011110011110;
        end
        1542: begin
            cosine_reg0 <= 36'sb11010100100001110100010100110011011;
            sine_reg0   <= 36'sb10001110101101110010001100001111101;
        end
        1543: begin
            cosine_reg0 <= 36'sb11010100011110010100000101011001001;
            sine_reg0   <= 36'sb10001110110010111111111111001011011;
        end
        1544: begin
            cosine_reg0 <= 36'sb11010100011010110011101101110010100;
            sine_reg0   <= 36'sb10001110111000001101101100100110111;
        end
        1545: begin
            cosine_reg0 <= 36'sb11010100010111010011001101111111111;
            sine_reg0   <= 36'sb10001110111101011011010100100001101;
        end
        1546: begin
            cosine_reg0 <= 36'sb11010100010011110010100110000001001;
            sine_reg0   <= 36'sb10001111000010101000110110111011111;
        end
        1547: begin
            cosine_reg0 <= 36'sb11010100010000010001110101110110101;
            sine_reg0   <= 36'sb10001111000111110110010011110101000;
        end
        1548: begin
            cosine_reg0 <= 36'sb11010100001100110000111101100000011;
            sine_reg0   <= 36'sb10001111001101000011101011001101000;
        end
        1549: begin
            cosine_reg0 <= 36'sb11010100001001001111111100111110100;
            sine_reg0   <= 36'sb10001111010010010000111101000011110;
        end
        1550: begin
            cosine_reg0 <= 36'sb11010100000101101110110100010001010;
            sine_reg0   <= 36'sb10001111010111011110001001011000111;
        end
        1551: begin
            cosine_reg0 <= 36'sb11010100000010001101100011011000101;
            sine_reg0   <= 36'sb10001111011100101011010000001100011;
        end
        1552: begin
            cosine_reg0 <= 36'sb11010011111110101100001010010100111;
            sine_reg0   <= 36'sb10001111100001111000010001011101111;
        end
        1553: begin
            cosine_reg0 <= 36'sb11010011111011001010101001000110001;
            sine_reg0   <= 36'sb10001111100111000101001101001101001;
        end
        1554: begin
            cosine_reg0 <= 36'sb11010011110111101000111111101100011;
            sine_reg0   <= 36'sb10001111101100010010000011011010001;
        end
        1555: begin
            cosine_reg0 <= 36'sb11010011110100000111001110000111111;
            sine_reg0   <= 36'sb10001111110001011110110100000100101;
        end
        1556: begin
            cosine_reg0 <= 36'sb11010011110000100101010100011000110;
            sine_reg0   <= 36'sb10001111110110101011011111001100010;
        end
        1557: begin
            cosine_reg0 <= 36'sb11010011101101000011010010011111010;
            sine_reg0   <= 36'sb10001111111011111000000100110001000;
        end
        1558: begin
            cosine_reg0 <= 36'sb11010011101001100001001000011011010;
            sine_reg0   <= 36'sb10010000000001000100100100110010101;
        end
        1559: begin
            cosine_reg0 <= 36'sb11010011100101111110110110001101001;
            sine_reg0   <= 36'sb10010000000110010000111111010000111;
        end
        1560: begin
            cosine_reg0 <= 36'sb11010011100010011100011011110100111;
            sine_reg0   <= 36'sb10010000001011011101010100001011101;
        end
        1561: begin
            cosine_reg0 <= 36'sb11010011011110111001111001010010101;
            sine_reg0   <= 36'sb10010000010000101001100011100010100;
        end
        1562: begin
            cosine_reg0 <= 36'sb11010011011011010111001110100110101;
            sine_reg0   <= 36'sb10010000010101110101101101010101101;
        end
        1563: begin
            cosine_reg0 <= 36'sb11010011010111110100011011110000111;
            sine_reg0   <= 36'sb10010000011011000001110001100100100;
        end
        1564: begin
            cosine_reg0 <= 36'sb11010011010100010001100000110001101;
            sine_reg0   <= 36'sb10010000100000001101110000001111000;
        end
        1565: begin
            cosine_reg0 <= 36'sb11010011010000101110011101101001000;
            sine_reg0   <= 36'sb10010000100101011001101001010100111;
        end
        1566: begin
            cosine_reg0 <= 36'sb11010011001101001011010010010111001;
            sine_reg0   <= 36'sb10010000101010100101011100110110001;
        end
        1567: begin
            cosine_reg0 <= 36'sb11010011001001100111111110111100000;
            sine_reg0   <= 36'sb10010000101111110001001010110010011;
        end
        1568: begin
            cosine_reg0 <= 36'sb11010011000110000100100011011000000;
            sine_reg0   <= 36'sb10010000110100111100110011001001100;
        end
        1569: begin
            cosine_reg0 <= 36'sb11010011000010100000111111101011001;
            sine_reg0   <= 36'sb10010000111010001000010101111011011;
        end
        1570: begin
            cosine_reg0 <= 36'sb11010010111110111101010011110101100;
            sine_reg0   <= 36'sb10010000111111010011110011000111101;
        end
        1571: begin
            cosine_reg0 <= 36'sb11010010111011011001011111110111010;
            sine_reg0   <= 36'sb10010001000100011111001010101110000;
        end
        1572: begin
            cosine_reg0 <= 36'sb11010010110111110101100011110000101;
            sine_reg0   <= 36'sb10010001001001101010011100101110101;
        end
        1573: begin
            cosine_reg0 <= 36'sb11010010110100010001011111100001110;
            sine_reg0   <= 36'sb10010001001110110101101001001001000;
        end
        1574: begin
            cosine_reg0 <= 36'sb11010010110000101101010011001010101;
            sine_reg0   <= 36'sb10010001010100000000101111111101000;
        end
        1575: begin
            cosine_reg0 <= 36'sb11010010101101001000111110101011100;
            sine_reg0   <= 36'sb10010001011001001011110001001010100;
        end
        1576: begin
            cosine_reg0 <= 36'sb11010010101001100100100010000100011;
            sine_reg0   <= 36'sb10010001011110010110101100110001010;
        end
        1577: begin
            cosine_reg0 <= 36'sb11010010100101111111111101010101101;
            sine_reg0   <= 36'sb10010001100011100001100010110001001;
        end
        1578: begin
            cosine_reg0 <= 36'sb11010010100010011011010000011111010;
            sine_reg0   <= 36'sb10010001101000101100010011001001110;
        end
        1579: begin
            cosine_reg0 <= 36'sb11010010011110110110011011100001011;
            sine_reg0   <= 36'sb10010001101101110110111101111011001;
        end
        1580: begin
            cosine_reg0 <= 36'sb11010010011011010001011110011100001;
            sine_reg0   <= 36'sb10010001110011000001100011000100111;
        end
        1581: begin
            cosine_reg0 <= 36'sb11010010010111101100011001001111101;
            sine_reg0   <= 36'sb10010001111000001100000010100111000;
        end
        1582: begin
            cosine_reg0 <= 36'sb11010010010100000111001011111100001;
            sine_reg0   <= 36'sb10010001111101010110011100100001001;
        end
        1583: begin
            cosine_reg0 <= 36'sb11010010010000100001110110100001101;
            sine_reg0   <= 36'sb10010010000010100000110000110011001;
        end
        1584: begin
            cosine_reg0 <= 36'sb11010010001100111100011001000000100;
            sine_reg0   <= 36'sb10010010000111101010111111011100110;
        end
        1585: begin
            cosine_reg0 <= 36'sb11010010001001010110110011011000100;
            sine_reg0   <= 36'sb10010010001100110101001000011101110;
        end
        1586: begin
            cosine_reg0 <= 36'sb11010010000101110001000101101010001;
            sine_reg0   <= 36'sb10010010010001111111001011110110001;
        end
        1587: begin
            cosine_reg0 <= 36'sb11010010000010001011001111110101011;
            sine_reg0   <= 36'sb10010010010111001001001001100101101;
        end
        1588: begin
            cosine_reg0 <= 36'sb11010001111110100101010001111010011;
            sine_reg0   <= 36'sb10010010011100010011000001101011111;
        end
        1589: begin
            cosine_reg0 <= 36'sb11010001111010111111001011111001010;
            sine_reg0   <= 36'sb10010010100001011100110100001000111;
        end
        1590: begin
            cosine_reg0 <= 36'sb11010001110111011000111101110010001;
            sine_reg0   <= 36'sb10010010100110100110100000111100010;
        end
        1591: begin
            cosine_reg0 <= 36'sb11010001110011110010100111100101010;
            sine_reg0   <= 36'sb10010010101011110000001000000110000;
        end
        1592: begin
            cosine_reg0 <= 36'sb11010001110000001100001001010010101;
            sine_reg0   <= 36'sb10010010110000111001101001100101110;
        end
        1593: begin
            cosine_reg0 <= 36'sb11010001101100100101100010111010100;
            sine_reg0   <= 36'sb10010010110110000011000101011011100;
        end
        1594: begin
            cosine_reg0 <= 36'sb11010001101000111110110100011101000;
            sine_reg0   <= 36'sb10010010111011001100011011100110110;
        end
        1595: begin
            cosine_reg0 <= 36'sb11010001100101010111111101111010010;
            sine_reg0   <= 36'sb10010011000000010101101100000111101;
        end
        1596: begin
            cosine_reg0 <= 36'sb11010001100001110000111111010010010;
            sine_reg0   <= 36'sb10010011000101011110110110111101101;
        end
        1597: begin
            cosine_reg0 <= 36'sb11010001011110001001111000100101011;
            sine_reg0   <= 36'sb10010011001010100111111100001000111;
        end
        1598: begin
            cosine_reg0 <= 36'sb11010001011010100010101001110011101;
            sine_reg0   <= 36'sb10010011001111110000111011101000111;
        end
        1599: begin
            cosine_reg0 <= 36'sb11010001010110111011010010111101001;
            sine_reg0   <= 36'sb10010011010100111001110101011101101;
        end
        1600: begin
            cosine_reg0 <= 36'sb11010001010011010011110100000010001;
            sine_reg0   <= 36'sb10010011011010000010101001100110111;
        end
        1601: begin
            cosine_reg0 <= 36'sb11010001001111101100001101000010101;
            sine_reg0   <= 36'sb10010011011111001011011000000100011;
        end
        1602: begin
            cosine_reg0 <= 36'sb11010001001100000100011101111110111;
            sine_reg0   <= 36'sb10010011100100010100000000110110000;
        end
        1603: begin
            cosine_reg0 <= 36'sb11010001001000011100100110110110111;
            sine_reg0   <= 36'sb10010011101001011100100011111011011;
        end
        1604: begin
            cosine_reg0 <= 36'sb11010001000100110100100111101011000;
            sine_reg0   <= 36'sb10010011101110100101000001010100101;
        end
        1605: begin
            cosine_reg0 <= 36'sb11010001000001001100100000011011001;
            sine_reg0   <= 36'sb10010011110011101101011001000001010;
        end
        1606: begin
            cosine_reg0 <= 36'sb11010000111101100100010001000111101;
            sine_reg0   <= 36'sb10010011111000110101101011000001010;
        end
        1607: begin
            cosine_reg0 <= 36'sb11010000111001111011111001110000100;
            sine_reg0   <= 36'sb10010011111101111101110111010100011;
        end
        1608: begin
            cosine_reg0 <= 36'sb11010000110110010011011010010101111;
            sine_reg0   <= 36'sb10010100000011000101111101111010011;
        end
        1609: begin
            cosine_reg0 <= 36'sb11010000110010101010110010111000000;
            sine_reg0   <= 36'sb10010100001000001101111110110011000;
        end
        1610: begin
            cosine_reg0 <= 36'sb11010000101111000010000011010111000;
            sine_reg0   <= 36'sb10010100001101010101111001111110010;
        end
        1611: begin
            cosine_reg0 <= 36'sb11010000101011011001001011110010111;
            sine_reg0   <= 36'sb10010100010010011101101111011011110;
        end
        1612: begin
            cosine_reg0 <= 36'sb11010000100111110000001100001011111;
            sine_reg0   <= 36'sb10010100010111100101011111001011011;
        end
        1613: begin
            cosine_reg0 <= 36'sb11010000100100000111000100100010001;
            sine_reg0   <= 36'sb10010100011100101101001001001100111;
        end
        1614: begin
            cosine_reg0 <= 36'sb11010000100000011101110100110101110;
            sine_reg0   <= 36'sb10010100100001110100101101100000001;
        end
        1615: begin
            cosine_reg0 <= 36'sb11010000011100110100011101000110111;
            sine_reg0   <= 36'sb10010100100110111100001100000100111;
        end
        1616: begin
            cosine_reg0 <= 36'sb11010000011001001010111101010101110;
            sine_reg0   <= 36'sb10010100101100000011100100111011000;
        end
        1617: begin
            cosine_reg0 <= 36'sb11010000010101100001010101100010011;
            sine_reg0   <= 36'sb10010100110001001010111000000010010;
        end
        1618: begin
            cosine_reg0 <= 36'sb11010000010001110111100101101101000;
            sine_reg0   <= 36'sb10010100110110010010000101011010011;
        end
        1619: begin
            cosine_reg0 <= 36'sb11010000001110001101101101110101101;
            sine_reg0   <= 36'sb10010100111011011001001101000011010;
        end
        1620: begin
            cosine_reg0 <= 36'sb11010000001010100011101101111100101;
            sine_reg0   <= 36'sb10010101000000100000001110111100101;
        end
        1621: begin
            cosine_reg0 <= 36'sb11010000000110111001100110000001111;
            sine_reg0   <= 36'sb10010101000101100111001011000110100;
        end
        1622: begin
            cosine_reg0 <= 36'sb11010000000011001111010110000101110;
            sine_reg0   <= 36'sb10010101001010101110000001100000011;
        end
        1623: begin
            cosine_reg0 <= 36'sb11001111111111100100111110001000001;
            sine_reg0   <= 36'sb10010101001111110100110010001010001;
        end
        1624: begin
            cosine_reg0 <= 36'sb11001111111011111010011110001001100;
            sine_reg0   <= 36'sb10010101010100111011011101000011110;
        end
        1625: begin
            cosine_reg0 <= 36'sb11001111111000001111110110001001101;
            sine_reg0   <= 36'sb10010101011010000010000010001100111;
        end
        1626: begin
            cosine_reg0 <= 36'sb11001111110100100101000110001000111;
            sine_reg0   <= 36'sb10010101011111001000100001100101011;
        end
        1627: begin
            cosine_reg0 <= 36'sb11001111110000111010001110000111011;
            sine_reg0   <= 36'sb10010101100100001110111011001101000;
        end
        1628: begin
            cosine_reg0 <= 36'sb11001111101101001111001110000101010;
            sine_reg0   <= 36'sb10010101101001010101001111000011101;
        end
        1629: begin
            cosine_reg0 <= 36'sb11001111101001100100000110000010101;
            sine_reg0   <= 36'sb10010101101110011011011101001001000;
        end
        1630: begin
            cosine_reg0 <= 36'sb11001111100101111000110101111111101;
            sine_reg0   <= 36'sb10010101110011100001100101011101000;
        end
        1631: begin
            cosine_reg0 <= 36'sb11001111100010001101011101111100100;
            sine_reg0   <= 36'sb10010101111000100111100111111111010;
        end
        1632: begin
            cosine_reg0 <= 36'sb11001111011110100001111101111001010;
            sine_reg0   <= 36'sb10010101111101101101100100101111110;
        end
        1633: begin
            cosine_reg0 <= 36'sb11001111011010110110010101110110000;
            sine_reg0   <= 36'sb10010110000010110011011011101110010;
        end
        1634: begin
            cosine_reg0 <= 36'sb11001111010111001010100101110011000;
            sine_reg0   <= 36'sb10010110000111111001001100111010100;
        end
        1635: begin
            cosine_reg0 <= 36'sb11001111010011011110101101110000011;
            sine_reg0   <= 36'sb10010110001100111110111000010100010;
        end
        1636: begin
            cosine_reg0 <= 36'sb11001111001111110010101101101110010;
            sine_reg0   <= 36'sb10010110010010000100011101111011100;
        end
        1637: begin
            cosine_reg0 <= 36'sb11001111001100000110100101101100110;
            sine_reg0   <= 36'sb10010110010111001001111101110000000;
        end
        1638: begin
            cosine_reg0 <= 36'sb11001111001000011010010101101100000;
            sine_reg0   <= 36'sb10010110011100001111010111110001011;
        end
        1639: begin
            cosine_reg0 <= 36'sb11001111000100101101111101101100010;
            sine_reg0   <= 36'sb10010110100001010100101011111111101;
        end
        1640: begin
            cosine_reg0 <= 36'sb11001111000001000001011101101101100;
            sine_reg0   <= 36'sb10010110100110011001111010011010011;
        end
        1641: begin
            cosine_reg0 <= 36'sb11001110111101010100110101110000000;
            sine_reg0   <= 36'sb10010110101011011111000011000001101;
        end
        1642: begin
            cosine_reg0 <= 36'sb11001110111001101000000101110011111;
            sine_reg0   <= 36'sb10010110110000100100000101110101000;
        end
        1643: begin
            cosine_reg0 <= 36'sb11001110110101111011001101111001001;
            sine_reg0   <= 36'sb10010110110101101001000010110100100;
        end
        1644: begin
            cosine_reg0 <= 36'sb11001110110010001110001110000000001;
            sine_reg0   <= 36'sb10010110111010101101111001111111110;
        end
        1645: begin
            cosine_reg0 <= 36'sb11001110101110100001000110001000111;
            sine_reg0   <= 36'sb10010110111111110010101011010110110;
        end
        1646: begin
            cosine_reg0 <= 36'sb11001110101010110011110110010011100;
            sine_reg0   <= 36'sb10010111000100110111010110111001000;
        end
        1647: begin
            cosine_reg0 <= 36'sb11001110100111000110011110100000010;
            sine_reg0   <= 36'sb10010111001001111011111100100110101;
        end
        1648: begin
            cosine_reg0 <= 36'sb11001110100011011000111110101111010;
            sine_reg0   <= 36'sb10010111001111000000011100011111010;
        end
        1649: begin
            cosine_reg0 <= 36'sb11001110011111101011010111000000100;
            sine_reg0   <= 36'sb10010111010100000100110110100010101;
        end
        1650: begin
            cosine_reg0 <= 36'sb11001110011011111101100111010100010;
            sine_reg0   <= 36'sb10010111011001001001001010110000110;
        end
        1651: begin
            cosine_reg0 <= 36'sb11001110011000001111101111101010110;
            sine_reg0   <= 36'sb10010111011110001101011001001001011;
        end
        1652: begin
            cosine_reg0 <= 36'sb11001110010100100001110000000011111;
            sine_reg0   <= 36'sb10010111100011010001100001101100001;
        end
        1653: begin
            cosine_reg0 <= 36'sb11001110010000110011101000100000000;
            sine_reg0   <= 36'sb10010111101000010101100100011001000;
        end
        1654: begin
            cosine_reg0 <= 36'sb11001110001101000101011000111111010;
            sine_reg0   <= 36'sb10010111101101011001100001001111110;
        end
        1655: begin
            cosine_reg0 <= 36'sb11001110001001010111000001100001101;
            sine_reg0   <= 36'sb10010111110010011101011000010000001;
        end
        1656: begin
            cosine_reg0 <= 36'sb11001110000101101000100010000111011;
            sine_reg0   <= 36'sb10010111110111100001001001011010000;
        end
        1657: begin
            cosine_reg0 <= 36'sb11001110000001111001111010110000101;
            sine_reg0   <= 36'sb10010111111100100100110100101101010;
        end
        1658: begin
            cosine_reg0 <= 36'sb11001101111110001011001011011101101;
            sine_reg0   <= 36'sb10011000000001101000011010001001100;
        end
        1659: begin
            cosine_reg0 <= 36'sb11001101111010011100010100001110010;
            sine_reg0   <= 36'sb10011000000110101011111001101110101;
        end
        1660: begin
            cosine_reg0 <= 36'sb11001101110110101101010101000010111;
            sine_reg0   <= 36'sb10011000001011101111010011011100100;
        end
        1661: begin
            cosine_reg0 <= 36'sb11001101110010111110001101111011100;
            sine_reg0   <= 36'sb10011000010000110010100111010010111;
        end
        1662: begin
            cosine_reg0 <= 36'sb11001101101111001110111110111000100;
            sine_reg0   <= 36'sb10011000010101110101110101010001100;
        end
        1663: begin
            cosine_reg0 <= 36'sb11001101101011011111100111111001110;
            sine_reg0   <= 36'sb10011000011010111000111101011000010;
        end
        1664: begin
            cosine_reg0 <= 36'sb11001101100111110000001000111111100;
            sine_reg0   <= 36'sb10011000011111111011111111100111000;
        end
        1665: begin
            cosine_reg0 <= 36'sb11001101100100000000100010001001111;
            sine_reg0   <= 36'sb10011000100100111110111011111101011;
        end
        1666: begin
            cosine_reg0 <= 36'sb11001101100000010000110011011001001;
            sine_reg0   <= 36'sb10011000101010000001110010011011011;
        end
        1667: begin
            cosine_reg0 <= 36'sb11001101011100100000111100101101010;
            sine_reg0   <= 36'sb10011000101111000100100011000000101;
        end
        1668: begin
            cosine_reg0 <= 36'sb11001101011000110000111110000110100;
            sine_reg0   <= 36'sb10011000110100000111001101101101000;
        end
        1669: begin
            cosine_reg0 <= 36'sb11001101010101000000110111100101000;
            sine_reg0   <= 36'sb10011000111001001001110010100000011;
        end
        1670: begin
            cosine_reg0 <= 36'sb11001101010001010000101001001000111;
            sine_reg0   <= 36'sb10011000111110001100010001011010100;
        end
        1671: begin
            cosine_reg0 <= 36'sb11001101001101100000010010110010010;
            sine_reg0   <= 36'sb10011001000011001110101010011011010;
        end
        1672: begin
            cosine_reg0 <= 36'sb11001101001001101111110100100001010;
            sine_reg0   <= 36'sb10011001001000010000111101100010010;
        end
        1673: begin
            cosine_reg0 <= 36'sb11001101000101111111001110010110001;
            sine_reg0   <= 36'sb10011001001101010011001010101111011;
        end
        1674: begin
            cosine_reg0 <= 36'sb11001101000010001110100000010000111;
            sine_reg0   <= 36'sb10011001010010010101010010000010101;
        end
        1675: begin
            cosine_reg0 <= 36'sb11001100111110011101101010010001110;
            sine_reg0   <= 36'sb10011001010111010111010011011011101;
        end
        1676: begin
            cosine_reg0 <= 36'sb11001100111010101100101100011000111;
            sine_reg0   <= 36'sb10011001011100011001001110111010001;
        end
        1677: begin
            cosine_reg0 <= 36'sb11001100110110111011100110100110011;
            sine_reg0   <= 36'sb10011001100001011011000100011110001;
        end
        1678: begin
            cosine_reg0 <= 36'sb11001100110011001010011000111010011;
            sine_reg0   <= 36'sb10011001100110011100110100000111010;
        end
        1679: begin
            cosine_reg0 <= 36'sb11001100101111011001000011010101001;
            sine_reg0   <= 36'sb10011001101011011110011101110101011;
        end
        1680: begin
            cosine_reg0 <= 36'sb11001100101011100111100101110110101;
            sine_reg0   <= 36'sb10011001110000100000000001101000011;
        end
        1681: begin
            cosine_reg0 <= 36'sb11001100100111110110000000011111001;
            sine_reg0   <= 36'sb10011001110101100001011111011111111;
        end
        1682: begin
            cosine_reg0 <= 36'sb11001100100100000100010011001110110;
            sine_reg0   <= 36'sb10011001111010100010110111011011111;
        end
        1683: begin
            cosine_reg0 <= 36'sb11001100100000010010011110000101101;
            sine_reg0   <= 36'sb10011001111111100100001001011100001;
        end
        1684: begin
            cosine_reg0 <= 36'sb11001100011100100000100001000100000;
            sine_reg0   <= 36'sb10011010000100100101010101100000011;
        end
        1685: begin
            cosine_reg0 <= 36'sb11001100011000101110011100001001110;
            sine_reg0   <= 36'sb10011010001001100110011011101000100;
        end
        1686: begin
            cosine_reg0 <= 36'sb11001100010100111100001111010111011;
            sine_reg0   <= 36'sb10011010001110100111011011110100010;
        end
        1687: begin
            cosine_reg0 <= 36'sb11001100010001001001111010101100110;
            sine_reg0   <= 36'sb10011010010011101000010110000011100;
        end
        1688: begin
            cosine_reg0 <= 36'sb11001100001101010111011110001010001;
            sine_reg0   <= 36'sb10011010011000101001001010010110000;
        end
        1689: begin
            cosine_reg0 <= 36'sb11001100001001100100111001101111101;
            sine_reg0   <= 36'sb10011010011101101001111000101011100;
        end
        1690: begin
            cosine_reg0 <= 36'sb11001100000101110010001101011101011;
            sine_reg0   <= 36'sb10011010100010101010100001000100000;
        end
        1691: begin
            cosine_reg0 <= 36'sb11001100000001111111011001010011101;
            sine_reg0   <= 36'sb10011010100111101011000011011111000;
        end
        1692: begin
            cosine_reg0 <= 36'sb11001011111110001100011101010010011;
            sine_reg0   <= 36'sb10011010101100101011011111111100101;
        end
        1693: begin
            cosine_reg0 <= 36'sb11001011111010011001011001011001111;
            sine_reg0   <= 36'sb10011010110001101011110110011100101;
        end
        1694: begin
            cosine_reg0 <= 36'sb11001011110110100110001101101010010;
            sine_reg0   <= 36'sb10011010110110101100000110111110101;
        end
        1695: begin
            cosine_reg0 <= 36'sb11001011110010110010111010000011101;
            sine_reg0   <= 36'sb10011010111011101100010001100010100;
        end
        1696: begin
            cosine_reg0 <= 36'sb11001011101110111111011110100110001;
            sine_reg0   <= 36'sb10011011000000101100010110001000001;
        end
        1697: begin
            cosine_reg0 <= 36'sb11001011101011001011111011010010000;
            sine_reg0   <= 36'sb10011011000101101100010100101111010;
        end
        1698: begin
            cosine_reg0 <= 36'sb11001011100111011000010000000111010;
            sine_reg0   <= 36'sb10011011001010101100001101010111110;
        end
        1699: begin
            cosine_reg0 <= 36'sb11001011100011100100011101000110010;
            sine_reg0   <= 36'sb10011011001111101100000000000001011;
        end
        1700: begin
            cosine_reg0 <= 36'sb11001011011111110000100010001110111;
            sine_reg0   <= 36'sb10011011010100101011101100101100000;
        end
        1701: begin
            cosine_reg0 <= 36'sb11001011011011111100011111100001011;
            sine_reg0   <= 36'sb10011011011001101011010011010111011;
        end
        1702: begin
            cosine_reg0 <= 36'sb11001011011000001000010100111110000;
            sine_reg0   <= 36'sb10011011011110101010110100000011010;
        end
        1703: begin
            cosine_reg0 <= 36'sb11001011010100010100000010100100110;
            sine_reg0   <= 36'sb10011011100011101010001110101111100;
        end
        1704: begin
            cosine_reg0 <= 36'sb11001011010000011111101000010101111;
            sine_reg0   <= 36'sb10011011101000101001100011011100000;
        end
        1705: begin
            cosine_reg0 <= 36'sb11001011001100101011000110010001011;
            sine_reg0   <= 36'sb10011011101101101000110010001000011;
        end
        1706: begin
            cosine_reg0 <= 36'sb11001011001000110110011100010111101;
            sine_reg0   <= 36'sb10011011110010100111111010110100101;
        end
        1707: begin
            cosine_reg0 <= 36'sb11001011000101000001101010101000101;
            sine_reg0   <= 36'sb10011011110111100110111101100000100;
        end
        1708: begin
            cosine_reg0 <= 36'sb11001011000001001100110001000100100;
            sine_reg0   <= 36'sb10011011111100100101111010001011110;
        end
        1709: begin
            cosine_reg0 <= 36'sb11001010111101010111101111101011100;
            sine_reg0   <= 36'sb10011100000001100100110000110110001;
        end
        1710: begin
            cosine_reg0 <= 36'sb11001010111001100010100110011101110;
            sine_reg0   <= 36'sb10011100000110100011100001011111101;
        end
        1711: begin
            cosine_reg0 <= 36'sb11001010110101101101010101011011010;
            sine_reg0   <= 36'sb10011100001011100010001100001000000;
        end
        1712: begin
            cosine_reg0 <= 36'sb11001010110001110111111100100100011;
            sine_reg0   <= 36'sb10011100010000100000110000101110111;
        end
        1713: begin
            cosine_reg0 <= 36'sb11001010101110000010011011111001001;
            sine_reg0   <= 36'sb10011100010101011111001111010100011;
        end
        1714: begin
            cosine_reg0 <= 36'sb11001010101010001100110011011001101;
            sine_reg0   <= 36'sb10011100011010011101100111111000000;
        end
        1715: begin
            cosine_reg0 <= 36'sb11001010100110010111000011000110001;
            sine_reg0   <= 36'sb10011100011111011011111010011001110;
        end
        1716: begin
            cosine_reg0 <= 36'sb11001010100010100001001010111110110;
            sine_reg0   <= 36'sb10011100100100011010000110111001011;
        end
        1717: begin
            cosine_reg0 <= 36'sb11001010011110101011001011000011101;
            sine_reg0   <= 36'sb10011100101001011000001101010110101;
        end
        1718: begin
            cosine_reg0 <= 36'sb11001010011010110101000011010100111;
            sine_reg0   <= 36'sb10011100101110010110001101110001011;
        end
        1719: begin
            cosine_reg0 <= 36'sb11001010010110111110110011110010110;
            sine_reg0   <= 36'sb10011100110011010100001000001001100;
        end
        1720: begin
            cosine_reg0 <= 36'sb11001010010011001000011100011101010;
            sine_reg0   <= 36'sb10011100111000010001111100011110101;
        end
        1721: begin
            cosine_reg0 <= 36'sb11001010001111010001111101010100101;
            sine_reg0   <= 36'sb10011100111101001111101010110000110;
        end
        1722: begin
            cosine_reg0 <= 36'sb11001010001011011011010110011001000;
            sine_reg0   <= 36'sb10011101000010001101010010111111100;
        end
        1723: begin
            cosine_reg0 <= 36'sb11001010000111100100100111101010100;
            sine_reg0   <= 36'sb10011101000111001010110101001010111;
        end
        1724: begin
            cosine_reg0 <= 36'sb11001010000011101101110001001001011;
            sine_reg0   <= 36'sb10011101001100001000010001010010101;
        end
        1725: begin
            cosine_reg0 <= 36'sb11001001111111110110110010110101101;
            sine_reg0   <= 36'sb10011101010001000101100111010110011;
        end
        1726: begin
            cosine_reg0 <= 36'sb11001001111011111111101100101111011;
            sine_reg0   <= 36'sb10011101010110000010110111010110010;
        end
        1727: begin
            cosine_reg0 <= 36'sb11001001111000001000011110110111000;
            sine_reg0   <= 36'sb10011101011011000000000001010001110;
        end
        1728: begin
            cosine_reg0 <= 36'sb11001001110100010001001001001100100;
            sine_reg0   <= 36'sb10011101011111111101000101001000111;
        end
        1729: begin
            cosine_reg0 <= 36'sb11001001110000011001101011110000000;
            sine_reg0   <= 36'sb10011101100100111010000010111011100;
        end
        1730: begin
            cosine_reg0 <= 36'sb11001001101100100010000110100001101;
            sine_reg0   <= 36'sb10011101101001110110111010101001010;
        end
        1731: begin
            cosine_reg0 <= 36'sb11001001101000101010011001100001110;
            sine_reg0   <= 36'sb10011101101110110011101100010001111;
        end
        1732: begin
            cosine_reg0 <= 36'sb11001001100100110010100100110000010;
            sine_reg0   <= 36'sb10011101110011110000010111110101100;
        end
        1733: begin
            cosine_reg0 <= 36'sb11001001100000111010101000001101011;
            sine_reg0   <= 36'sb10011101111000101100111101010011101;
        end
        1734: begin
            cosine_reg0 <= 36'sb11001001011101000010100011111001010;
            sine_reg0   <= 36'sb10011101111101101001011100101100010;
        end
        1735: begin
            cosine_reg0 <= 36'sb11001001011001001010010111110100001;
            sine_reg0   <= 36'sb10011110000010100101110101111111001;
        end
        1736: begin
            cosine_reg0 <= 36'sb11001001010101010010000011111110001;
            sine_reg0   <= 36'sb10011110000111100010001001001100000;
        end
        1737: begin
            cosine_reg0 <= 36'sb11001001010001011001101000010111010;
            sine_reg0   <= 36'sb10011110001100011110010110010010110;
        end
        1738: begin
            cosine_reg0 <= 36'sb11001001001101100001000100111111110;
            sine_reg0   <= 36'sb10011110010001011010011101010011001;
        end
        1739: begin
            cosine_reg0 <= 36'sb11001001001001101000011001110111111;
            sine_reg0   <= 36'sb10011110010110010110011110001101000;
        end
        1740: begin
            cosine_reg0 <= 36'sb11001001000101101111100110111111101;
            sine_reg0   <= 36'sb10011110011011010010011001000000010;
        end
        1741: begin
            cosine_reg0 <= 36'sb11001001000001110110101100010111010;
            sine_reg0   <= 36'sb10011110100000001110001101101100100;
        end
        1742: begin
            cosine_reg0 <= 36'sb11001000111101111101101001111110111;
            sine_reg0   <= 36'sb10011110100101001001111100010001110;
        end
        1743: begin
            cosine_reg0 <= 36'sb11001000111010000100011111110110100;
            sine_reg0   <= 36'sb10011110101010000101100100101111101;
        end
        1744: begin
            cosine_reg0 <= 36'sb11001000110110001011001101111110100;
            sine_reg0   <= 36'sb10011110101111000001000111000110001;
        end
        1745: begin
            cosine_reg0 <= 36'sb11001000110010010001110100010111000;
            sine_reg0   <= 36'sb10011110110011111100100011010100111;
        end
        1746: begin
            cosine_reg0 <= 36'sb11001000101110011000010011000000000;
            sine_reg0   <= 36'sb10011110111000110111111001011011110;
        end
        1747: begin
            cosine_reg0 <= 36'sb11001000101010011110101001111001110;
            sine_reg0   <= 36'sb10011110111101110011001001011010110;
        end
        1748: begin
            cosine_reg0 <= 36'sb11001000100110100100111001000100011;
            sine_reg0   <= 36'sb10011111000010101110010011010001011;
        end
        1749: begin
            cosine_reg0 <= 36'sb11001000100010101011000000100000000;
            sine_reg0   <= 36'sb10011111000111101001010110111111101;
        end
        1750: begin
            cosine_reg0 <= 36'sb11001000011110110001000000001100111;
            sine_reg0   <= 36'sb10011111001100100100010100100101010;
        end
        1751: begin
            cosine_reg0 <= 36'sb11001000011010110110111000001011000;
            sine_reg0   <= 36'sb10011111010001011111001100000010000;
        end
        1752: begin
            cosine_reg0 <= 36'sb11001000010110111100101000011010101;
            sine_reg0   <= 36'sb10011111010110011001111101010101111;
        end
        1753: begin
            cosine_reg0 <= 36'sb11001000010011000010010000111011111;
            sine_reg0   <= 36'sb10011111011011010100101000100000100;
        end
        1754: begin
            cosine_reg0 <= 36'sb11001000001111000111110001101111000;
            sine_reg0   <= 36'sb10011111100000001111001101100001110;
        end
        1755: begin
            cosine_reg0 <= 36'sb11001000001011001101001010110100000;
            sine_reg0   <= 36'sb10011111100101001001101100011001100;
        end
        1756: begin
            cosine_reg0 <= 36'sb11001000000111010010011100001011001;
            sine_reg0   <= 36'sb10011111101010000100000101000111100;
        end
        1757: begin
            cosine_reg0 <= 36'sb11001000000011010111100101110100011;
            sine_reg0   <= 36'sb10011111101110111110010111101011100;
        end
        1758: begin
            cosine_reg0 <= 36'sb11000111111111011100100111110000001;
            sine_reg0   <= 36'sb10011111110011111000100100000101011;
        end
        1759: begin
            cosine_reg0 <= 36'sb11000111111011100001100001111110011;
            sine_reg0   <= 36'sb10011111111000110010101010010101000;
        end
        1760: begin
            cosine_reg0 <= 36'sb11000111110111100110010100011111011;
            sine_reg0   <= 36'sb10011111111101101100101010011010001;
        end
        1761: begin
            cosine_reg0 <= 36'sb11000111110011101010111111010011010;
            sine_reg0   <= 36'sb10100000000010100110100100010100100;
        end
        1762: begin
            cosine_reg0 <= 36'sb11000111101111101111100010011010000;
            sine_reg0   <= 36'sb10100000000111100000011000000100000;
        end
        1763: begin
            cosine_reg0 <= 36'sb11000111101011110011111101110011111;
            sine_reg0   <= 36'sb10100000001100011010000101101000011;
        end
        1764: begin
            cosine_reg0 <= 36'sb11000111100111111000010001100001001;
            sine_reg0   <= 36'sb10100000010001010011101101000001101;
        end
        1765: begin
            cosine_reg0 <= 36'sb11000111100011111100011101100001111;
            sine_reg0   <= 36'sb10100000010110001101001110001111010;
        end
        1766: begin
            cosine_reg0 <= 36'sb11000111100000000000100001110110001;
            sine_reg0   <= 36'sb10100000011011000110101001010001011;
        end
        1767: begin
            cosine_reg0 <= 36'sb11000111011100000100011110011110010;
            sine_reg0   <= 36'sb10100000011111111111111110000111101;
        end
        1768: begin
            cosine_reg0 <= 36'sb11000111011000001000010011011010001;
            sine_reg0   <= 36'sb10100000100100111001001100110001111;
        end
        1769: begin
            cosine_reg0 <= 36'sb11000111010100001100000000101010001;
            sine_reg0   <= 36'sb10100000101001110010010101001111111;
        end
        1770: begin
            cosine_reg0 <= 36'sb11000111010000001111100110001110011;
            sine_reg0   <= 36'sb10100000101110101011010111100001100;
        end
        1771: begin
            cosine_reg0 <= 36'sb11000111001100010011000100000111000;
            sine_reg0   <= 36'sb10100000110011100100010011100110100;
        end
        1772: begin
            cosine_reg0 <= 36'sb11000111001000010110011010010100001;
            sine_reg0   <= 36'sb10100000111000011101001001011110110;
        end
        1773: begin
            cosine_reg0 <= 36'sb11000111000100011001101000110101111;
            sine_reg0   <= 36'sb10100000111101010101111001001010001;
        end
        1774: begin
            cosine_reg0 <= 36'sb11000111000000011100101111101100011;
            sine_reg0   <= 36'sb10100001000010001110100010101000010;
        end
        1775: begin
            cosine_reg0 <= 36'sb11000110111100011111101110111000000;
            sine_reg0   <= 36'sb10100001000111000111000101111001001;
        end
        1776: begin
            cosine_reg0 <= 36'sb11000110111000100010100110011000101;
            sine_reg0   <= 36'sb10100001001011111111100010111100011;
        end
        1777: begin
            cosine_reg0 <= 36'sb11000110110100100101010110001110100;
            sine_reg0   <= 36'sb10100001010000110111111001110010000;
        end
        1778: begin
            cosine_reg0 <= 36'sb11000110110000100111111110011001111;
            sine_reg0   <= 36'sb10100001010101110000001010011001101;
        end
        1779: begin
            cosine_reg0 <= 36'sb11000110101100101010011110111010111;
            sine_reg0   <= 36'sb10100001011010101000010100110011010;
        end
        1780: begin
            cosine_reg0 <= 36'sb11000110101000101100110111110001100;
            sine_reg0   <= 36'sb10100001011111100000011000111110100;
        end
        1781: begin
            cosine_reg0 <= 36'sb11000110100100101111001000111110001;
            sine_reg0   <= 36'sb10100001100100011000010110111011011;
        end
        1782: begin
            cosine_reg0 <= 36'sb11000110100000110001010010100000110;
            sine_reg0   <= 36'sb10100001101001010000001110101001101;
        end
        1783: begin
            cosine_reg0 <= 36'sb11000110011100110011010100011001100;
            sine_reg0   <= 36'sb10100001101110001000000000001000111;
        end
        1784: begin
            cosine_reg0 <= 36'sb11000110011000110101001110101000101;
            sine_reg0   <= 36'sb10100001110010111111101011011001010;
        end
        1785: begin
            cosine_reg0 <= 36'sb11000110010100110111000001001110010;
            sine_reg0   <= 36'sb10100001110111110111010000011010011;
        end
        1786: begin
            cosine_reg0 <= 36'sb11000110010000111000101100001010101;
            sine_reg0   <= 36'sb10100001111100101110101111001100000;
        end
        1787: begin
            cosine_reg0 <= 36'sb11000110001100111010001111011101101;
            sine_reg0   <= 36'sb10100010000001100110000111101110001;
        end
        1788: begin
            cosine_reg0 <= 36'sb11000110001000111011101011000111110;
            sine_reg0   <= 36'sb10100010000110011101011010000000100;
        end
        1789: begin
            cosine_reg0 <= 36'sb11000110000100111100111111001000111;
            sine_reg0   <= 36'sb10100010001011010100100110000010111;
        end
        1790: begin
            cosine_reg0 <= 36'sb11000110000000111110001011100001010;
            sine_reg0   <= 36'sb10100010010000001011101011110101000;
        end
        1791: begin
            cosine_reg0 <= 36'sb11000101111100111111010000010001001;
            sine_reg0   <= 36'sb10100010010101000010101011010110111;
        end
        1792: begin
            cosine_reg0 <= 36'sb11000101111001000000001101011000100;
            sine_reg0   <= 36'sb10100010011001111001100100101000010;
        end
        1793: begin
            cosine_reg0 <= 36'sb11000101110101000001000010110111110;
            sine_reg0   <= 36'sb10100010011110110000010111101000111;
        end
        1794: begin
            cosine_reg0 <= 36'sb11000101110001000001110000101110110;
            sine_reg0   <= 36'sb10100010100011100111000100011000100;
        end
        1795: begin
            cosine_reg0 <= 36'sb11000101101101000010010110111101110;
            sine_reg0   <= 36'sb10100010101000011101101010110111001;
        end
        1796: begin
            cosine_reg0 <= 36'sb11000101101001000010110101100101000;
            sine_reg0   <= 36'sb10100010101101010100001011000100100;
        end
        1797: begin
            cosine_reg0 <= 36'sb11000101100101000011001100100100100;
            sine_reg0   <= 36'sb10100010110010001010100101000000011;
        end
        1798: begin
            cosine_reg0 <= 36'sb11000101100001000011011011111100101;
            sine_reg0   <= 36'sb10100010110111000000111000101010100;
        end
        1799: begin
            cosine_reg0 <= 36'sb11000101011101000011100011101101011;
            sine_reg0   <= 36'sb10100010111011110111000110000010111;
        end
        1800: begin
            cosine_reg0 <= 36'sb11000101011001000011100011110110111;
            sine_reg0   <= 36'sb10100011000000101101001101001001010;
        end
        1801: begin
            cosine_reg0 <= 36'sb11000101010101000011011100011001011;
            sine_reg0   <= 36'sb10100011000101100011001101111101011;
        end
        1802: begin
            cosine_reg0 <= 36'sb11000101010001000011001101010100111;
            sine_reg0   <= 36'sb10100011001010011001001000011111001;
        end
        1803: begin
            cosine_reg0 <= 36'sb11000101001101000010110110101001110;
            sine_reg0   <= 36'sb10100011001111001110111100101110010;
        end
        1804: begin
            cosine_reg0 <= 36'sb11000101001001000010011000011000000;
            sine_reg0   <= 36'sb10100011010100000100101010101010101;
        end
        1805: begin
            cosine_reg0 <= 36'sb11000101000101000001110010011111111;
            sine_reg0   <= 36'sb10100011011000111010010010010100001;
        end
        1806: begin
            cosine_reg0 <= 36'sb11000101000001000001000101000001011;
            sine_reg0   <= 36'sb10100011011101101111110011101010011;
        end
        1807: begin
            cosine_reg0 <= 36'sb11000100111101000000001111111100111;
            sine_reg0   <= 36'sb10100011100010100101001110101101010;
        end
        1808: begin
            cosine_reg0 <= 36'sb11000100111000111111010011010010011;
            sine_reg0   <= 36'sb10100011100111011010100011011100101;
        end
        1809: begin
            cosine_reg0 <= 36'sb11000100110100111110001111000010000;
            sine_reg0   <= 36'sb10100011101100001111110001111000011;
        end
        1810: begin
            cosine_reg0 <= 36'sb11000100110000111101000011001100000;
            sine_reg0   <= 36'sb10100011110001000100111010000000010;
        end
        1811: begin
            cosine_reg0 <= 36'sb11000100101100111011101111110000101;
            sine_reg0   <= 36'sb10100011110101111001111011110100000;
        end
        1812: begin
            cosine_reg0 <= 36'sb11000100101000111010010100101111110;
            sine_reg0   <= 36'sb10100011111010101110110111010011011;
        end
        1813: begin
            cosine_reg0 <= 36'sb11000100100100111000110010001001110;
            sine_reg0   <= 36'sb10100011111111100011101100011110011;
        end
        1814: begin
            cosine_reg0 <= 36'sb11000100100000110111000111111110110;
            sine_reg0   <= 36'sb10100100000100011000011011010100111;
        end
        1815: begin
            cosine_reg0 <= 36'sb11000100011100110101010110001110110;
            sine_reg0   <= 36'sb10100100001001001101000011110110011;
        end
        1816: begin
            cosine_reg0 <= 36'sb11000100011000110011011100111010001;
            sine_reg0   <= 36'sb10100100001110000001100110000011000;
        end
        1817: begin
            cosine_reg0 <= 36'sb11000100010100110001011100000001000;
            sine_reg0   <= 36'sb10100100010010110110000001111010010;
        end
        1818: begin
            cosine_reg0 <= 36'sb11000100010000101111010011100011011;
            sine_reg0   <= 36'sb10100100010111101010010111011100010;
        end
        1819: begin
            cosine_reg0 <= 36'sb11000100001100101101000011100001100;
            sine_reg0   <= 36'sb10100100011100011110100110101000110;
        end
        1820: begin
            cosine_reg0 <= 36'sb11000100001000101010101011111011100;
            sine_reg0   <= 36'sb10100100100001010010101111011111011;
        end
        1821: begin
            cosine_reg0 <= 36'sb11000100000100101000001100110001101;
            sine_reg0   <= 36'sb10100100100110000110110010000000001;
        end
        1822: begin
            cosine_reg0 <= 36'sb11000100000000100101100110000011111;
            sine_reg0   <= 36'sb10100100101010111010101110001010101;
        end
        1823: begin
            cosine_reg0 <= 36'sb11000011111100100010110111110010100;
            sine_reg0   <= 36'sb10100100101111101110100011111111000;
        end
        1824: begin
            cosine_reg0 <= 36'sb11000011111000100000000001111101110;
            sine_reg0   <= 36'sb10100100110100100010010011011100110;
        end
        1825: begin
            cosine_reg0 <= 36'sb11000011110100011101000100100101101;
            sine_reg0   <= 36'sb10100100111001010101111100100011111;
        end
        1826: begin
            cosine_reg0 <= 36'sb11000011110000011001111111101010010;
            sine_reg0   <= 36'sb10100100111110001001011111010100001;
        end
        1827: begin
            cosine_reg0 <= 36'sb11000011101100010110110011001100000;
            sine_reg0   <= 36'sb10100101000010111100111011101101011;
        end
        1828: begin
            cosine_reg0 <= 36'sb11000011101000010011011111001010110;
            sine_reg0   <= 36'sb10100101000111110000010001101111011;
        end
        1829: begin
            cosine_reg0 <= 36'sb11000011100100010000000011100111000;
            sine_reg0   <= 36'sb10100101001100100011100001011001111;
        end
        1830: begin
            cosine_reg0 <= 36'sb11000011100000001100100000100000100;
            sine_reg0   <= 36'sb10100101010001010110101010101100110;
        end
        1831: begin
            cosine_reg0 <= 36'sb11000011011100001000110101110111110;
            sine_reg0   <= 36'sb10100101010110001001101101101000000;
        end
        1832: begin
            cosine_reg0 <= 36'sb11000011011000000101000011101100110;
            sine_reg0   <= 36'sb10100101011010111100101010001011001;
        end
        1833: begin
            cosine_reg0 <= 36'sb11000011010100000001001001111111101;
            sine_reg0   <= 36'sb10100101011111101111100000010110001;
        end
        1834: begin
            cosine_reg0 <= 36'sb11000011001111111101001000110000101;
            sine_reg0   <= 36'sb10100101100100100010010000001000111;
        end
        1835: begin
            cosine_reg0 <= 36'sb11000011001011111000111111111111111;
            sine_reg0   <= 36'sb10100101101001010100111001100011000;
        end
        1836: begin
            cosine_reg0 <= 36'sb11000011000111110100101111101101100;
            sine_reg0   <= 36'sb10100101101110000111011100100100011;
        end
        1837: begin
            cosine_reg0 <= 36'sb11000011000011110000010111111001110;
            sine_reg0   <= 36'sb10100101110010111001111001001101000;
        end
        1838: begin
            cosine_reg0 <= 36'sb11000010111111101011111000100100101;
            sine_reg0   <= 36'sb10100101110111101100001111011100011;
        end
        1839: begin
            cosine_reg0 <= 36'sb11000010111011100111010001101110011;
            sine_reg0   <= 36'sb10100101111100011110011111010010101;
        end
        1840: begin
            cosine_reg0 <= 36'sb11000010110111100010100011010111010;
            sine_reg0   <= 36'sb10100110000001010000101000101111010;
        end
        1841: begin
            cosine_reg0 <= 36'sb11000010110011011101101101011111001;
            sine_reg0   <= 36'sb10100110000110000010101011110010011;
        end
        1842: begin
            cosine_reg0 <= 36'sb11000010101111011000110000000110100;
            sine_reg0   <= 36'sb10100110001010110100101000011011101;
        end
        1843: begin
            cosine_reg0 <= 36'sb11000010101011010011101011001101011;
            sine_reg0   <= 36'sb10100110001111100110011110101010111;
        end
        1844: begin
            cosine_reg0 <= 36'sb11000010100111001110011110110011110;
            sine_reg0   <= 36'sb10100110010100011000001110100000000;
        end
        1845: begin
            cosine_reg0 <= 36'sb11000010100011001001001010111010001;
            sine_reg0   <= 36'sb10100110011001001001110111111010101;
        end
        1846: begin
            cosine_reg0 <= 36'sb11000010011111000011101111100000011;
            sine_reg0   <= 36'sb10100110011101111011011010111010111;
        end
        1847: begin
            cosine_reg0 <= 36'sb11000010011010111110001100100110110;
            sine_reg0   <= 36'sb10100110100010101100110111100000010;
        end
        1848: begin
            cosine_reg0 <= 36'sb11000010010110111000100010001101011;
            sine_reg0   <= 36'sb10100110100111011110001101101010110;
        end
        1849: begin
            cosine_reg0 <= 36'sb11000010010010110010110000010100100;
            sine_reg0   <= 36'sb10100110101100001111011101011010000;
        end
        1850: begin
            cosine_reg0 <= 36'sb11000010001110101100110110111100010;
            sine_reg0   <= 36'sb10100110110001000000100110101110001;
        end
        1851: begin
            cosine_reg0 <= 36'sb11000010001010100110110110000100101;
            sine_reg0   <= 36'sb10100110110101110001101001100110110;
        end
        1852: begin
            cosine_reg0 <= 36'sb11000010000110100000101101101110000;
            sine_reg0   <= 36'sb10100110111010100010100110000011101;
        end
        1853: begin
            cosine_reg0 <= 36'sb11000010000010011010011101111000100;
            sine_reg0   <= 36'sb10100110111111010011011100000100110;
        end
        1854: begin
            cosine_reg0 <= 36'sb11000001111110010100000110100100010;
            sine_reg0   <= 36'sb10100111000100000100001011101001110;
        end
        1855: begin
            cosine_reg0 <= 36'sb11000001111010001101100111110001010;
            sine_reg0   <= 36'sb10100111001000110100110100110010101;
        end
        1856: begin
            cosine_reg0 <= 36'sb11000001110110000111000001011111111;
            sine_reg0   <= 36'sb10100111001101100101010111011111000;
        end
        1857: begin
            cosine_reg0 <= 36'sb11000001110010000000010011110000010;
            sine_reg0   <= 36'sb10100111010010010101110011101110111;
        end
        1858: begin
            cosine_reg0 <= 36'sb11000001101101111001011110100010011;
            sine_reg0   <= 36'sb10100111010111000110001001100010000;
        end
        1859: begin
            cosine_reg0 <= 36'sb11000001101001110010100001110110101;
            sine_reg0   <= 36'sb10100111011011110110011000111000001;
        end
        1860: begin
            cosine_reg0 <= 36'sb11000001100101101011011101101101000;
            sine_reg0   <= 36'sb10100111100000100110100001110001001;
        end
        1861: begin
            cosine_reg0 <= 36'sb11000001100001100100010010000101110;
            sine_reg0   <= 36'sb10100111100101010110100100001100111;
        end
        1862: begin
            cosine_reg0 <= 36'sb11000001011101011100111111000001000;
            sine_reg0   <= 36'sb10100111101010000110100000001011001;
        end
        1863: begin
            cosine_reg0 <= 36'sb11000001011001010101100100011110111;
            sine_reg0   <= 36'sb10100111101110110110010101101011101;
        end
        1864: begin
            cosine_reg0 <= 36'sb11000001010101001110000010011111101;
            sine_reg0   <= 36'sb10100111110011100110000100101110011;
        end
        1865: begin
            cosine_reg0 <= 36'sb11000001010001000110011001000011010;
            sine_reg0   <= 36'sb10100111111000010101101101010011000;
        end
        1866: begin
            cosine_reg0 <= 36'sb11000001001100111110101000001010000;
            sine_reg0   <= 36'sb10100111111101000101001111011001011;
        end
        1867: begin
            cosine_reg0 <= 36'sb11000001001000110110101111110100001;
            sine_reg0   <= 36'sb10101000000001110100101011000001011;
        end
        1868: begin
            cosine_reg0 <= 36'sb11000001000100101110110000000001110;
            sine_reg0   <= 36'sb10101000000110100100000000001010110;
        end
        1869: begin
            cosine_reg0 <= 36'sb11000001000000100110101000110010111;
            sine_reg0   <= 36'sb10101000001011010011001110110101011;
        end
        1870: begin
            cosine_reg0 <= 36'sb11000000111100011110011010000111110;
            sine_reg0   <= 36'sb10101000010000000010010111000001000;
        end
        1871: begin
            cosine_reg0 <= 36'sb11000000111000010110000100000000101;
            sine_reg0   <= 36'sb10101000010100110001011000101101100;
        end
        1872: begin
            cosine_reg0 <= 36'sb11000000110100001101100110011101101;
            sine_reg0   <= 36'sb10101000011001100000010011111010110;
        end
        1873: begin
            cosine_reg0 <= 36'sb11000000110000000101000001011110110;
            sine_reg0   <= 36'sb10101000011110001111001000101000011;
        end
        1874: begin
            cosine_reg0 <= 36'sb11000000101011111100010101000100011;
            sine_reg0   <= 36'sb10101000100010111101110110110110011;
        end
        1875: begin
            cosine_reg0 <= 36'sb11000000100111110011100001001110100;
            sine_reg0   <= 36'sb10101000100111101100011110100100100;
        end
        1876: begin
            cosine_reg0 <= 36'sb11000000100011101010100101111101011;
            sine_reg0   <= 36'sb10101000101100011010111111110010101;
        end
        1877: begin
            cosine_reg0 <= 36'sb11000000011111100001100011010001001;
            sine_reg0   <= 36'sb10101000110001001001011010100000100;
        end
        1878: begin
            cosine_reg0 <= 36'sb11000000011011011000011001001010000;
            sine_reg0   <= 36'sb10101000110101110111101110101101111;
        end
        1879: begin
            cosine_reg0 <= 36'sb11000000010111001111000111101000000;
            sine_reg0   <= 36'sb10101000111010100101111100011010101;
        end
        1880: begin
            cosine_reg0 <= 36'sb11000000010011000101101110101011011;
            sine_reg0   <= 36'sb10101000111111010100000011100110110;
        end
        1881: begin
            cosine_reg0 <= 36'sb11000000001110111100001110010100010;
            sine_reg0   <= 36'sb10101001000100000010000100010001110;
        end
        1882: begin
            cosine_reg0 <= 36'sb11000000001010110010100110100010111;
            sine_reg0   <= 36'sb10101001001000101111111110011011110;
        end
        1883: begin
            cosine_reg0 <= 36'sb11000000000110101000110111010111010;
            sine_reg0   <= 36'sb10101001001101011101110010000100011;
        end
        1884: begin
            cosine_reg0 <= 36'sb11000000000010011111000000110001101;
            sine_reg0   <= 36'sb10101001010010001011011111001011011;
        end
        1885: begin
            cosine_reg0 <= 36'sb10111111111110010101000010110010010;
            sine_reg0   <= 36'sb10101001010110111001000101110000110;
        end
        1886: begin
            cosine_reg0 <= 36'sb10111111111010001010111101011001010;
            sine_reg0   <= 36'sb10101001011011100110100101110100011;
        end
        1887: begin
            cosine_reg0 <= 36'sb10111111110110000000110000100110101;
            sine_reg0   <= 36'sb10101001100000010011111111010101110;
        end
        1888: begin
            cosine_reg0 <= 36'sb10111111110001110110011100011010101;
            sine_reg0   <= 36'sb10101001100101000001010010010101000;
        end
        1889: begin
            cosine_reg0 <= 36'sb10111111101101101100000000110101100;
            sine_reg0   <= 36'sb10101001101001101110011110110001111;
        end
        1890: begin
            cosine_reg0 <= 36'sb10111111101001100001011101110111010;
            sine_reg0   <= 36'sb10101001101110011011100100101100000;
        end
        1891: begin
            cosine_reg0 <= 36'sb10111111100101010110110011100000010;
            sine_reg0   <= 36'sb10101001110011001000100100000011100;
        end
        1892: begin
            cosine_reg0 <= 36'sb10111111100001001100000001110000100;
            sine_reg0   <= 36'sb10101001110111110101011100111000000;
        end
        1893: begin
            cosine_reg0 <= 36'sb10111111011101000001001000101000001;
            sine_reg0   <= 36'sb10101001111100100010001111001001010;
        end
        1894: begin
            cosine_reg0 <= 36'sb10111111011000110110001000000111011;
            sine_reg0   <= 36'sb10101010000001001110111010110111010;
        end
        1895: begin
            cosine_reg0 <= 36'sb10111111010100101011000000001110100;
            sine_reg0   <= 36'sb10101010000101111011100000000001110;
        end
        1896: begin
            cosine_reg0 <= 36'sb10111111010000011111110000111101011;
            sine_reg0   <= 36'sb10101010001010100111111110101000101;
        end
        1897: begin
            cosine_reg0 <= 36'sb10111111001100010100011010010100100;
            sine_reg0   <= 36'sb10101010001111010100010110101011100;
        end
        1898: begin
            cosine_reg0 <= 36'sb10111111001000001000111100010011110;
            sine_reg0   <= 36'sb10101010010100000000101000001010011;
        end
        1899: begin
            cosine_reg0 <= 36'sb10111111000011111101010110111011100;
            sine_reg0   <= 36'sb10101010011000101100110011000101001;
        end
        1900: begin
            cosine_reg0 <= 36'sb10111110111111110001101010001011111;
            sine_reg0   <= 36'sb10101010011101011000110111011011011;
        end
        1901: begin
            cosine_reg0 <= 36'sb10111110111011100101110110000100111;
            sine_reg0   <= 36'sb10101010100010000100110101001101000;
        end
        1902: begin
            cosine_reg0 <= 36'sb10111110110111011001111010100110110;
            sine_reg0   <= 36'sb10101010100110110000101100011001111;
        end
        1903: begin
            cosine_reg0 <= 36'sb10111110110011001101110111110001110;
            sine_reg0   <= 36'sb10101010101011011100011101000001111;
        end
        1904: begin
            cosine_reg0 <= 36'sb10111110101111000001101101100110000;
            sine_reg0   <= 36'sb10101010110000001000000111000100101;
        end
        1905: begin
            cosine_reg0 <= 36'sb10111110101010110101011100000011101;
            sine_reg0   <= 36'sb10101010110100110011101010100010001;
        end
        1906: begin
            cosine_reg0 <= 36'sb10111110100110101001000011001010110;
            sine_reg0   <= 36'sb10101010111001011111000111011010001;
        end
        1907: begin
            cosine_reg0 <= 36'sb10111110100010011100100010111011101;
            sine_reg0   <= 36'sb10101010111110001010011101101100100;
        end
        1908: begin
            cosine_reg0 <= 36'sb10111110011110001111111011010110010;
            sine_reg0   <= 36'sb10101011000010110101101101011000111;
        end
        1909: begin
            cosine_reg0 <= 36'sb10111110011010000011001100011011000;
            sine_reg0   <= 36'sb10101011000111100000110110011111011;
        end
        1910: begin
            cosine_reg0 <= 36'sb10111110010101110110010110001001111;
            sine_reg0   <= 36'sb10101011001100001011111000111111101;
        end
        1911: begin
            cosine_reg0 <= 36'sb10111110010001101001011000100011010;
            sine_reg0   <= 36'sb10101011010000110110110100111001011;
        end
        1912: begin
            cosine_reg0 <= 36'sb10111110001101011100010011100111000;
            sine_reg0   <= 36'sb10101011010101100001101010001100101;
        end
        1913: begin
            cosine_reg0 <= 36'sb10111110001001001111000111010101100;
            sine_reg0   <= 36'sb10101011011010001100011000111001001;
        end
        1914: begin
            cosine_reg0 <= 36'sb10111110000101000001110011101110110;
            sine_reg0   <= 36'sb10101011011110110111000000111110110;
        end
        1915: begin
            cosine_reg0 <= 36'sb10111110000000110100011000110011000;
            sine_reg0   <= 36'sb10101011100011100001100010011101001;
        end
        1916: begin
            cosine_reg0 <= 36'sb10111101111100100110110110100010100;
            sine_reg0   <= 36'sb10101011101000001011111101010100010;
        end
        1917: begin
            cosine_reg0 <= 36'sb10111101111000011001001100111101010;
            sine_reg0   <= 36'sb10101011101100110110010001100100000;
        end
        1918: begin
            cosine_reg0 <= 36'sb10111101110100001011011100000011101;
            sine_reg0   <= 36'sb10101011110001100000011111001100000;
        end
        1919: begin
            cosine_reg0 <= 36'sb10111101101111111101100011110101100;
            sine_reg0   <= 36'sb10101011110110001010100110001100001;
        end
        1920: begin
            cosine_reg0 <= 36'sb10111101101011101111100100010011010;
            sine_reg0   <= 36'sb10101011111010110100100110100100011;
        end
        1921: begin
            cosine_reg0 <= 36'sb10111101100111100001011101011101000;
            sine_reg0   <= 36'sb10101011111111011110100000010100010;
        end
        1922: begin
            cosine_reg0 <= 36'sb10111101100011010011001111010010110;
            sine_reg0   <= 36'sb10101100000100001000010011011011111;
        end
        1923: begin
            cosine_reg0 <= 36'sb10111101011111000100111001110101000;
            sine_reg0   <= 36'sb10101100001000110001111111111011000;
        end
        1924: begin
            cosine_reg0 <= 36'sb10111101011010110110011101000011100;
            sine_reg0   <= 36'sb10101100001101011011100101110001010;
        end
        1925: begin
            cosine_reg0 <= 36'sb10111101010110100111111000111110110;
            sine_reg0   <= 36'sb10101100010010000101000100111110101;
        end
        1926: begin
            cosine_reg0 <= 36'sb10111101010010011001001101100110111;
            sine_reg0   <= 36'sb10101100010110101110011101100011000;
        end
        1927: begin
            cosine_reg0 <= 36'sb10111101001110001010011010111011110;
            sine_reg0   <= 36'sb10101100011011010111101111011110000;
        end
        1928: begin
            cosine_reg0 <= 36'sb10111101001001111011100000111101111;
            sine_reg0   <= 36'sb10101100100000000000111010101111101;
        end
        1929: begin
            cosine_reg0 <= 36'sb10111101000101101100011111101101010;
            sine_reg0   <= 36'sb10101100100100101001111111010111101;
        end
        1930: begin
            cosine_reg0 <= 36'sb10111101000001011101010111001010001;
            sine_reg0   <= 36'sb10101100101001010010111101010101110;
        end
        1931: begin
            cosine_reg0 <= 36'sb10111100111101001110000111010100100;
            sine_reg0   <= 36'sb10101100101101111011110100101010000;
        end
        1932: begin
            cosine_reg0 <= 36'sb10111100111000111110110000001100101;
            sine_reg0   <= 36'sb10101100110010100100100101010100000;
        end
        1933: begin
            cosine_reg0 <= 36'sb10111100110100101111010001110010110;
            sine_reg0   <= 36'sb10101100110111001101001111010011101;
        end
        1934: begin
            cosine_reg0 <= 36'sb10111100110000011111101100000111000;
            sine_reg0   <= 36'sb10101100111011110101110010101000110;
        end
        1935: begin
            cosine_reg0 <= 36'sb10111100101100001111111111001001100;
            sine_reg0   <= 36'sb10101101000000011110001111010011010;
        end
        1936: begin
            cosine_reg0 <= 36'sb10111100101000000000001010111010011;
            sine_reg0   <= 36'sb10101101000101000110100101010010111;
        end
        1937: begin
            cosine_reg0 <= 36'sb10111100100011110000001111011001111;
            sine_reg0   <= 36'sb10101101001001101110110100100111011;
        end
        1938: begin
            cosine_reg0 <= 36'sb10111100011111100000001100101000001;
            sine_reg0   <= 36'sb10101101001110010110111101010000101;
        end
        1939: begin
            cosine_reg0 <= 36'sb10111100011011010000000010100101010;
            sine_reg0   <= 36'sb10101101010010111110111111001110100;
        end
        1940: begin
            cosine_reg0 <= 36'sb10111100010110111111110001010001100;
            sine_reg0   <= 36'sb10101101010111100110111010100000110;
        end
        1941: begin
            cosine_reg0 <= 36'sb10111100010010101111011000101101000;
            sine_reg0   <= 36'sb10101101011100001110101111000111010;
        end
        1942: begin
            cosine_reg0 <= 36'sb10111100001110011110111000110111110;
            sine_reg0   <= 36'sb10101101100000110110011101000001111;
        end
        1943: begin
            cosine_reg0 <= 36'sb10111100001010001110010001110010010;
            sine_reg0   <= 36'sb10101101100101011110000100010000010;
        end
        1944: begin
            cosine_reg0 <= 36'sb10111100000101111101100011011100011;
            sine_reg0   <= 36'sb10101101101010000101100100110010011;
        end
        1945: begin
            cosine_reg0 <= 36'sb10111100000001101100101101110110100;
            sine_reg0   <= 36'sb10101101101110101100111110101000000;
        end
        1946: begin
            cosine_reg0 <= 36'sb10111011111101011011110001000000101;
            sine_reg0   <= 36'sb10101101110011010100010001110001000;
        end
        1947: begin
            cosine_reg0 <= 36'sb10111011111001001010101100111011000;
            sine_reg0   <= 36'sb10101101110111111011011110001101001;
        end
        1948: begin
            cosine_reg0 <= 36'sb10111011110100111001100001100101110;
            sine_reg0   <= 36'sb10101101111100100010100011111100010;
        end
        1949: begin
            cosine_reg0 <= 36'sb10111011110000101000001111000001001;
            sine_reg0   <= 36'sb10101110000001001001100010111110010;
        end
        1950: begin
            cosine_reg0 <= 36'sb10111011101100010110110101001101001;
            sine_reg0   <= 36'sb10101110000101110000011011010010110;
        end
        1951: begin
            cosine_reg0 <= 36'sb10111011101000000101010100001010000;
            sine_reg0   <= 36'sb10101110001010010111001100111001110;
        end
        1952: begin
            cosine_reg0 <= 36'sb10111011100011110011101011111000000;
            sine_reg0   <= 36'sb10101110001110111101110111110011001;
        end
        1953: begin
            cosine_reg0 <= 36'sb10111011011111100001111100010111010;
            sine_reg0   <= 36'sb10101110010011100100011011111110100;
        end
        1954: begin
            cosine_reg0 <= 36'sb10111011011011010000000101100111110;
            sine_reg0   <= 36'sb10101110011000001010111001011011110;
        end
        1955: begin
            cosine_reg0 <= 36'sb10111011010110111110000111101001111;
            sine_reg0   <= 36'sb10101110011100110001010000001010110;
        end
        1956: begin
            cosine_reg0 <= 36'sb10111011010010101100000010011101110;
            sine_reg0   <= 36'sb10101110100001010111100000001011011;
        end
        1957: begin
            cosine_reg0 <= 36'sb10111011001110011001110110000011011;
            sine_reg0   <= 36'sb10101110100101111101101001011101011;
        end
        1958: begin
            cosine_reg0 <= 36'sb10111011001010000111100010011011001;
            sine_reg0   <= 36'sb10101110101010100011101100000000100;
        end
        1959: begin
            cosine_reg0 <= 36'sb10111011000101110101000111100101001;
            sine_reg0   <= 36'sb10101110101111001001100111110100110;
        end
        1960: begin
            cosine_reg0 <= 36'sb10111011000001100010100101100001011;
            sine_reg0   <= 36'sb10101110110011101111011100111001111;
        end
        1961: begin
            cosine_reg0 <= 36'sb10111010111101001111111100010000010;
            sine_reg0   <= 36'sb10101110111000010101001011001111101;
        end
        1962: begin
            cosine_reg0 <= 36'sb10111010111000111101001011110001111;
            sine_reg0   <= 36'sb10101110111100111010110010110101111;
        end
        1963: begin
            cosine_reg0 <= 36'sb10111010110100101010010100000110010;
            sine_reg0   <= 36'sb10101111000001100000010011101100100;
        end
        1964: begin
            cosine_reg0 <= 36'sb10111010110000010111010101001101110;
            sine_reg0   <= 36'sb10101111000110000101101101110011001;
        end
        1965: begin
            cosine_reg0 <= 36'sb10111010101100000100001111001000011;
            sine_reg0   <= 36'sb10101111001010101011000001001001111;
        end
        1966: begin
            cosine_reg0 <= 36'sb10111010100111110001000001110110011;
            sine_reg0   <= 36'sb10101111001111010000001101110000011;
        end
        1967: begin
            cosine_reg0 <= 36'sb10111010100011011101101101011000000;
            sine_reg0   <= 36'sb10101111010011110101010011100110100;
        end
        1968: begin
            cosine_reg0 <= 36'sb10111010011111001010010001101101001;
            sine_reg0   <= 36'sb10101111011000011010010010101100000;
        end
        1969: begin
            cosine_reg0 <= 36'sb10111010011010110110101110110110010;
            sine_reg0   <= 36'sb10101111011100111111001011000000111;
        end
        1970: begin
            cosine_reg0 <= 36'sb10111010010110100011000100110011011;
            sine_reg0   <= 36'sb10101111100001100011111100100100110;
        end
        1971: begin
            cosine_reg0 <= 36'sb10111010010010001111010011100100110;
            sine_reg0   <= 36'sb10101111100110001000100111010111100;
        end
        1972: begin
            cosine_reg0 <= 36'sb10111010001101111011011011001010100;
            sine_reg0   <= 36'sb10101111101010101101001011011001001;
        end
        1973: begin
            cosine_reg0 <= 36'sb10111010001001100111011011100100101;
            sine_reg0   <= 36'sb10101111101111010001101000101001001;
        end
        1974: begin
            cosine_reg0 <= 36'sb10111010000101010011010100110011101;
            sine_reg0   <= 36'sb10101111110011110101111111000111101;
        end
        1975: begin
            cosine_reg0 <= 36'sb10111010000000111111000110110111011;
            sine_reg0   <= 36'sb10101111111000011010001110110100011;
        end
        1976: begin
            cosine_reg0 <= 36'sb10111001111100101010110001110000001;
            sine_reg0   <= 36'sb10101111111100111110010111101111001;
        end
        1977: begin
            cosine_reg0 <= 36'sb10111001111000010110010101011110001;
            sine_reg0   <= 36'sb10110000000001100010011001110111101;
        end
        1978: begin
            cosine_reg0 <= 36'sb10111001110100000001110010000001100;
            sine_reg0   <= 36'sb10110000000110000110010101001101111;
        end
        1979: begin
            cosine_reg0 <= 36'sb10111001101111101101000111011010011;
            sine_reg0   <= 36'sb10110000001010101010001001110001101;
        end
        1980: begin
            cosine_reg0 <= 36'sb10111001101011011000010101101000111;
            sine_reg0   <= 36'sb10110000001111001101110111100010110;
        end
        1981: begin
            cosine_reg0 <= 36'sb10111001100111000011011100101101011;
            sine_reg0   <= 36'sb10110000010011110001011110100001000;
        end
        1982: begin
            cosine_reg0 <= 36'sb10111001100010101110011100100111110;
            sine_reg0   <= 36'sb10110000011000010100111110101100010;
        end
        1983: begin
            cosine_reg0 <= 36'sb10111001011110011001010101011000011;
            sine_reg0   <= 36'sb10110000011100111000011000000100010;
        end
        1984: begin
            cosine_reg0 <= 36'sb10111001011010000100000110111111011;
            sine_reg0   <= 36'sb10110000100001011011101010101000111;
        end
        1985: begin
            cosine_reg0 <= 36'sb10111001010101101110110001011100111;
            sine_reg0   <= 36'sb10110000100101111110110110011001111;
        end
        1986: begin
            cosine_reg0 <= 36'sb10111001010001011001010100110001001;
            sine_reg0   <= 36'sb10110000101010100001111011010111010;
        end
        1987: begin
            cosine_reg0 <= 36'sb10111001001101000011110000111100010;
            sine_reg0   <= 36'sb10110000101111000100111001100000110;
        end
        1988: begin
            cosine_reg0 <= 36'sb10111001001000101110000101111110011;
            sine_reg0   <= 36'sb10110000110011100111110000110110001;
        end
        1989: begin
            cosine_reg0 <= 36'sb10111001000100011000010011110111101;
            sine_reg0   <= 36'sb10110000111000001010100001010111010;
        end
        1990: begin
            cosine_reg0 <= 36'sb10111001000000000010011010101000010;
            sine_reg0   <= 36'sb10110000111100101101001011000011111;
        end
        1991: begin
            cosine_reg0 <= 36'sb10111000111011101100011010010000100;
            sine_reg0   <= 36'sb10110001000001001111101101111100000;
        end
        1992: begin
            cosine_reg0 <= 36'sb10111000110111010110010010110000011;
            sine_reg0   <= 36'sb10110001000101110010001001111111010;
        end
        1993: begin
            cosine_reg0 <= 36'sb10111000110011000000000100001000001;
            sine_reg0   <= 36'sb10110001001010010100011111001101101;
        end
        1994: begin
            cosine_reg0 <= 36'sb10111000101110101001101110010111111;
            sine_reg0   <= 36'sb10110001001110110110101101100110111;
        end
        1995: begin
            cosine_reg0 <= 36'sb10111000101010010011010001011111111;
            sine_reg0   <= 36'sb10110001010011011000110101001010110;
        end
        1996: begin
            cosine_reg0 <= 36'sb10111000100101111100101101100000010;
            sine_reg0   <= 36'sb10110001010111111010110101111001010;
        end
        1997: begin
            cosine_reg0 <= 36'sb10111000100001100110000010011001001;
            sine_reg0   <= 36'sb10110001011100011100101111110010000;
        end
        1998: begin
            cosine_reg0 <= 36'sb10111000011101001111010000001010101;
            sine_reg0   <= 36'sb10110001100000111110100010110101000;
        end
        1999: begin
            cosine_reg0 <= 36'sb10111000011000111000010110110101001;
            sine_reg0   <= 36'sb10110001100101100000001111000010000;
        end
        2000: begin
            cosine_reg0 <= 36'sb10111000010100100001010110011000101;
            sine_reg0   <= 36'sb10110001101010000001110100011000110;
        end
        2001: begin
            cosine_reg0 <= 36'sb10111000010000001010001110110101011;
            sine_reg0   <= 36'sb10110001101110100011010010111001010;
        end
        2002: begin
            cosine_reg0 <= 36'sb10111000001011110011000000001011011;
            sine_reg0   <= 36'sb10110001110011000100101010100011001;
        end
        2003: begin
            cosine_reg0 <= 36'sb10111000000111011011101010011011000;
            sine_reg0   <= 36'sb10110001110111100101111011010110011;
        end
        2004: begin
            cosine_reg0 <= 36'sb10111000000011000100001101100100011;
            sine_reg0   <= 36'sb10110001111100000111000101010010110;
        end
        2005: begin
            cosine_reg0 <= 36'sb10110111111110101100101001100111101;
            sine_reg0   <= 36'sb10110010000000101000001000011000000;
        end
        2006: begin
            cosine_reg0 <= 36'sb10110111111010010100111110100100111;
            sine_reg0   <= 36'sb10110010000101001001000100100110001;
        end
        2007: begin
            cosine_reg0 <= 36'sb10110111110101111101001100011100011;
            sine_reg0   <= 36'sb10110010001001101001111001111100110;
        end
        2008: begin
            cosine_reg0 <= 36'sb10110111110001100101010011001110010;
            sine_reg0   <= 36'sb10110010001110001010101000011011111;
        end
        2009: begin
            cosine_reg0 <= 36'sb10110111101101001101010010111010101;
            sine_reg0   <= 36'sb10110010010010101011010000000011010;
        end
        2010: begin
            cosine_reg0 <= 36'sb10110111101000110101001011100001110;
            sine_reg0   <= 36'sb10110010010111001011110000110010110;
        end
        2011: begin
            cosine_reg0 <= 36'sb10110111100100011100111101000011110;
            sine_reg0   <= 36'sb10110010011011101100001010101010001;
        end
        2012: begin
            cosine_reg0 <= 36'sb10110111100000000100100111100000111;
            sine_reg0   <= 36'sb10110010100000001100011101101001001;
        end
        2013: begin
            cosine_reg0 <= 36'sb10110111011011101100001010111001010;
            sine_reg0   <= 36'sb10110010100100101100101001101111111;
        end
        2014: begin
            cosine_reg0 <= 36'sb10110111010111010011100111001100111;
            sine_reg0   <= 36'sb10110010101001001100101110111101111;
        end
        2015: begin
            cosine_reg0 <= 36'sb10110111010010111010111100011100010;
            sine_reg0   <= 36'sb10110010101101101100101101010011001;
        end
        2016: begin
            cosine_reg0 <= 36'sb10110111001110100010001010100111010;
            sine_reg0   <= 36'sb10110010110010001100100100101111011;
        end
        2017: begin
            cosine_reg0 <= 36'sb10110111001010001001010001101110001;
            sine_reg0   <= 36'sb10110010110110101100010101010010101;
        end
        2018: begin
            cosine_reg0 <= 36'sb10110111000101110000010001110001001;
            sine_reg0   <= 36'sb10110010111011001011111110111100100;
        end
        2019: begin
            cosine_reg0 <= 36'sb10110111000001010111001010110000011;
            sine_reg0   <= 36'sb10110010111111101011100001101100111;
        end
        2020: begin
            cosine_reg0 <= 36'sb10110110111100111101111100101100001;
            sine_reg0   <= 36'sb10110011000100001010111101100011101;
        end
        2021: begin
            cosine_reg0 <= 36'sb10110110111000100100100111100100011;
            sine_reg0   <= 36'sb10110011001000101010010010100000100;
        end
        2022: begin
            cosine_reg0 <= 36'sb10110110110100001011001011011001011;
            sine_reg0   <= 36'sb10110011001101001001100000100011011;
        end
        2023: begin
            cosine_reg0 <= 36'sb10110110101111110001101000001011010;
            sine_reg0   <= 36'sb10110011010001101000100111101100001;
        end
        2024: begin
            cosine_reg0 <= 36'sb10110110101011010111111101111010010;
            sine_reg0   <= 36'sb10110011010110000111100111111010100;
        end
        2025: begin
            cosine_reg0 <= 36'sb10110110100110111110001100100110100;
            sine_reg0   <= 36'sb10110011011010100110100001001110011;
        end
        2026: begin
            cosine_reg0 <= 36'sb10110110100010100100010100010000010;
            sine_reg0   <= 36'sb10110011011111000101010011100111100;
        end
        2027: begin
            cosine_reg0 <= 36'sb10110110011110001010010100110111100;
            sine_reg0   <= 36'sb10110011100011100011111111000101111;
        end
        2028: begin
            cosine_reg0 <= 36'sb10110110011001110000001110011100101;
            sine_reg0   <= 36'sb10110011101000000010100011101001001;
        end
        2029: begin
            cosine_reg0 <= 36'sb10110110010101010110000000111111101;
            sine_reg0   <= 36'sb10110011101100100001000001010001010;
        end
        2030: begin
            cosine_reg0 <= 36'sb10110110010000111011101100100000110;
            sine_reg0   <= 36'sb10110011110000111111010111111101111;
        end
        2031: begin
            cosine_reg0 <= 36'sb10110110001100100001010001000000001;
            sine_reg0   <= 36'sb10110011110101011101100111101111000;
        end
        2032: begin
            cosine_reg0 <= 36'sb10110110001000000110101110011110000;
            sine_reg0   <= 36'sb10110011111001111011110000100100100;
        end
        2033: begin
            cosine_reg0 <= 36'sb10110110000011101100000100111010011;
            sine_reg0   <= 36'sb10110011111110011001110010011110000;
        end
        2034: begin
            cosine_reg0 <= 36'sb10110101111111010001010100010101110;
            sine_reg0   <= 36'sb10110100000010110111101101011011011;
        end
        2035: begin
            cosine_reg0 <= 36'sb10110101111010110110011100101111111;
            sine_reg0   <= 36'sb10110100000111010101100001011100101;
        end
        2036: begin
            cosine_reg0 <= 36'sb10110101110110011011011110001001010;
            sine_reg0   <= 36'sb10110100001011110011001110100001011;
        end
        2037: begin
            cosine_reg0 <= 36'sb10110101110010000000011000100001111;
            sine_reg0   <= 36'sb10110100010000010000110100101001101;
        end
        2038: begin
            cosine_reg0 <= 36'sb10110101101101100101001011111010000;
            sine_reg0   <= 36'sb10110100010100101110010011110101000;
        end
        2039: begin
            cosine_reg0 <= 36'sb10110101101001001001111000010001111;
            sine_reg0   <= 36'sb10110100011001001011101100000011100;
        end
        2040: begin
            cosine_reg0 <= 36'sb10110101100100101110011101101001011;
            sine_reg0   <= 36'sb10110100011101101000111101010101000;
        end
        2041: begin
            cosine_reg0 <= 36'sb10110101100000010010111100000001000;
            sine_reg0   <= 36'sb10110100100010000110000111101001001;
        end
        2042: begin
            cosine_reg0 <= 36'sb10110101011011110111010011011000110;
            sine_reg0   <= 36'sb10110100100110100011001010111111110;
        end
        2043: begin
            cosine_reg0 <= 36'sb10110101010111011011100011110000110;
            sine_reg0   <= 36'sb10110100101011000000000111011000111;
        end
        2044: begin
            cosine_reg0 <= 36'sb10110101010010111111101101001001010;
            sine_reg0   <= 36'sb10110100101111011100111100110100001;
        end
        2045: begin
            cosine_reg0 <= 36'sb10110101001110100011101111100010100;
            sine_reg0   <= 36'sb10110100110011111001101011010001011;
        end
        2046: begin
            cosine_reg0 <= 36'sb10110101001010000111101010111100101;
            sine_reg0   <= 36'sb10110100111000010110010010110000101;
        end
        2047: begin
            cosine_reg0 <= 36'sb10110101000101101011011111010111101;
            sine_reg0   <= 36'sb10110100111100110010110011010001100;
        end
        2048: begin
            cosine_reg0 <= 36'sb10110101000001001111001100110011111;
            sine_reg0   <= 36'sb10110101000001001111001100110011111;
        end
        2049: begin
            cosine_reg0 <= 36'sb10110100111100110010110011010001100;
            sine_reg0   <= 36'sb10110101000101101011011111010111101;
        end
        2050: begin
            cosine_reg0 <= 36'sb10110100111000010110010010110000101;
            sine_reg0   <= 36'sb10110101001010000111101010111100101;
        end
        2051: begin
            cosine_reg0 <= 36'sb10110100110011111001101011010001011;
            sine_reg0   <= 36'sb10110101001110100011101111100010100;
        end
        2052: begin
            cosine_reg0 <= 36'sb10110100101111011100111100110100001;
            sine_reg0   <= 36'sb10110101010010111111101101001001010;
        end
        2053: begin
            cosine_reg0 <= 36'sb10110100101011000000000111011000111;
            sine_reg0   <= 36'sb10110101010111011011100011110000110;
        end
        2054: begin
            cosine_reg0 <= 36'sb10110100100110100011001010111111110;
            sine_reg0   <= 36'sb10110101011011110111010011011000110;
        end
        2055: begin
            cosine_reg0 <= 36'sb10110100100010000110000111101001001;
            sine_reg0   <= 36'sb10110101100000010010111100000001000;
        end
        2056: begin
            cosine_reg0 <= 36'sb10110100011101101000111101010101000;
            sine_reg0   <= 36'sb10110101100100101110011101101001011;
        end
        2057: begin
            cosine_reg0 <= 36'sb10110100011001001011101100000011100;
            sine_reg0   <= 36'sb10110101101001001001111000010001111;
        end
        2058: begin
            cosine_reg0 <= 36'sb10110100010100101110010011110101000;
            sine_reg0   <= 36'sb10110101101101100101001011111010000;
        end
        2059: begin
            cosine_reg0 <= 36'sb10110100010000010000110100101001101;
            sine_reg0   <= 36'sb10110101110010000000011000100001111;
        end
        2060: begin
            cosine_reg0 <= 36'sb10110100001011110011001110100001011;
            sine_reg0   <= 36'sb10110101110110011011011110001001010;
        end
        2061: begin
            cosine_reg0 <= 36'sb10110100000111010101100001011100101;
            sine_reg0   <= 36'sb10110101111010110110011100101111111;
        end
        2062: begin
            cosine_reg0 <= 36'sb10110100000010110111101101011011011;
            sine_reg0   <= 36'sb10110101111111010001010100010101110;
        end
        2063: begin
            cosine_reg0 <= 36'sb10110011111110011001110010011110000;
            sine_reg0   <= 36'sb10110110000011101100000100111010011;
        end
        2064: begin
            cosine_reg0 <= 36'sb10110011111001111011110000100100100;
            sine_reg0   <= 36'sb10110110001000000110101110011110000;
        end
        2065: begin
            cosine_reg0 <= 36'sb10110011110101011101100111101111000;
            sine_reg0   <= 36'sb10110110001100100001010001000000001;
        end
        2066: begin
            cosine_reg0 <= 36'sb10110011110000111111010111111101111;
            sine_reg0   <= 36'sb10110110010000111011101100100000110;
        end
        2067: begin
            cosine_reg0 <= 36'sb10110011101100100001000001010001010;
            sine_reg0   <= 36'sb10110110010101010110000000111111101;
        end
        2068: begin
            cosine_reg0 <= 36'sb10110011101000000010100011101001001;
            sine_reg0   <= 36'sb10110110011001110000001110011100101;
        end
        2069: begin
            cosine_reg0 <= 36'sb10110011100011100011111111000101111;
            sine_reg0   <= 36'sb10110110011110001010010100110111100;
        end
        2070: begin
            cosine_reg0 <= 36'sb10110011011111000101010011100111100;
            sine_reg0   <= 36'sb10110110100010100100010100010000010;
        end
        2071: begin
            cosine_reg0 <= 36'sb10110011011010100110100001001110011;
            sine_reg0   <= 36'sb10110110100110111110001100100110100;
        end
        2072: begin
            cosine_reg0 <= 36'sb10110011010110000111100111111010100;
            sine_reg0   <= 36'sb10110110101011010111111101111010010;
        end
        2073: begin
            cosine_reg0 <= 36'sb10110011010001101000100111101100001;
            sine_reg0   <= 36'sb10110110101111110001101000001011010;
        end
        2074: begin
            cosine_reg0 <= 36'sb10110011001101001001100000100011011;
            sine_reg0   <= 36'sb10110110110100001011001011011001011;
        end
        2075: begin
            cosine_reg0 <= 36'sb10110011001000101010010010100000100;
            sine_reg0   <= 36'sb10110110111000100100100111100100011;
        end
        2076: begin
            cosine_reg0 <= 36'sb10110011000100001010111101100011101;
            sine_reg0   <= 36'sb10110110111100111101111100101100001;
        end
        2077: begin
            cosine_reg0 <= 36'sb10110010111111101011100001101100111;
            sine_reg0   <= 36'sb10110111000001010111001010110000011;
        end
        2078: begin
            cosine_reg0 <= 36'sb10110010111011001011111110111100100;
            sine_reg0   <= 36'sb10110111000101110000010001110001001;
        end
        2079: begin
            cosine_reg0 <= 36'sb10110010110110101100010101010010101;
            sine_reg0   <= 36'sb10110111001010001001010001101110001;
        end
        2080: begin
            cosine_reg0 <= 36'sb10110010110010001100100100101111011;
            sine_reg0   <= 36'sb10110111001110100010001010100111010;
        end
        2081: begin
            cosine_reg0 <= 36'sb10110010101101101100101101010011001;
            sine_reg0   <= 36'sb10110111010010111010111100011100010;
        end
        2082: begin
            cosine_reg0 <= 36'sb10110010101001001100101110111101111;
            sine_reg0   <= 36'sb10110111010111010011100111001100111;
        end
        2083: begin
            cosine_reg0 <= 36'sb10110010100100101100101001101111111;
            sine_reg0   <= 36'sb10110111011011101100001010111001010;
        end
        2084: begin
            cosine_reg0 <= 36'sb10110010100000001100011101101001001;
            sine_reg0   <= 36'sb10110111100000000100100111100000111;
        end
        2085: begin
            cosine_reg0 <= 36'sb10110010011011101100001010101010001;
            sine_reg0   <= 36'sb10110111100100011100111101000011110;
        end
        2086: begin
            cosine_reg0 <= 36'sb10110010010111001011110000110010110;
            sine_reg0   <= 36'sb10110111101000110101001011100001110;
        end
        2087: begin
            cosine_reg0 <= 36'sb10110010010010101011010000000011010;
            sine_reg0   <= 36'sb10110111101101001101010010111010101;
        end
        2088: begin
            cosine_reg0 <= 36'sb10110010001110001010101000011011111;
            sine_reg0   <= 36'sb10110111110001100101010011001110010;
        end
        2089: begin
            cosine_reg0 <= 36'sb10110010001001101001111001111100110;
            sine_reg0   <= 36'sb10110111110101111101001100011100011;
        end
        2090: begin
            cosine_reg0 <= 36'sb10110010000101001001000100100110001;
            sine_reg0   <= 36'sb10110111111010010100111110100100111;
        end
        2091: begin
            cosine_reg0 <= 36'sb10110010000000101000001000011000000;
            sine_reg0   <= 36'sb10110111111110101100101001100111101;
        end
        2092: begin
            cosine_reg0 <= 36'sb10110001111100000111000101010010110;
            sine_reg0   <= 36'sb10111000000011000100001101100100011;
        end
        2093: begin
            cosine_reg0 <= 36'sb10110001110111100101111011010110011;
            sine_reg0   <= 36'sb10111000000111011011101010011011000;
        end
        2094: begin
            cosine_reg0 <= 36'sb10110001110011000100101010100011001;
            sine_reg0   <= 36'sb10111000001011110011000000001011011;
        end
        2095: begin
            cosine_reg0 <= 36'sb10110001101110100011010010111001010;
            sine_reg0   <= 36'sb10111000010000001010001110110101011;
        end
        2096: begin
            cosine_reg0 <= 36'sb10110001101010000001110100011000110;
            sine_reg0   <= 36'sb10111000010100100001010110011000101;
        end
        2097: begin
            cosine_reg0 <= 36'sb10110001100101100000001111000010000;
            sine_reg0   <= 36'sb10111000011000111000010110110101001;
        end
        2098: begin
            cosine_reg0 <= 36'sb10110001100000111110100010110101000;
            sine_reg0   <= 36'sb10111000011101001111010000001010101;
        end
        2099: begin
            cosine_reg0 <= 36'sb10110001011100011100101111110010000;
            sine_reg0   <= 36'sb10111000100001100110000010011001001;
        end
        2100: begin
            cosine_reg0 <= 36'sb10110001010111111010110101111001010;
            sine_reg0   <= 36'sb10111000100101111100101101100000010;
        end
        2101: begin
            cosine_reg0 <= 36'sb10110001010011011000110101001010110;
            sine_reg0   <= 36'sb10111000101010010011010001011111111;
        end
        2102: begin
            cosine_reg0 <= 36'sb10110001001110110110101101100110111;
            sine_reg0   <= 36'sb10111000101110101001101110010111111;
        end
        2103: begin
            cosine_reg0 <= 36'sb10110001001010010100011111001101101;
            sine_reg0   <= 36'sb10111000110011000000000100001000001;
        end
        2104: begin
            cosine_reg0 <= 36'sb10110001000101110010001001111111010;
            sine_reg0   <= 36'sb10111000110111010110010010110000011;
        end
        2105: begin
            cosine_reg0 <= 36'sb10110001000001001111101101111100000;
            sine_reg0   <= 36'sb10111000111011101100011010010000100;
        end
        2106: begin
            cosine_reg0 <= 36'sb10110000111100101101001011000011111;
            sine_reg0   <= 36'sb10111001000000000010011010101000010;
        end
        2107: begin
            cosine_reg0 <= 36'sb10110000111000001010100001010111010;
            sine_reg0   <= 36'sb10111001000100011000010011110111101;
        end
        2108: begin
            cosine_reg0 <= 36'sb10110000110011100111110000110110001;
            sine_reg0   <= 36'sb10111001001000101110000101111110011;
        end
        2109: begin
            cosine_reg0 <= 36'sb10110000101111000100111001100000110;
            sine_reg0   <= 36'sb10111001001101000011110000111100010;
        end
        2110: begin
            cosine_reg0 <= 36'sb10110000101010100001111011010111010;
            sine_reg0   <= 36'sb10111001010001011001010100110001001;
        end
        2111: begin
            cosine_reg0 <= 36'sb10110000100101111110110110011001111;
            sine_reg0   <= 36'sb10111001010101101110110001011100111;
        end
        2112: begin
            cosine_reg0 <= 36'sb10110000100001011011101010101000111;
            sine_reg0   <= 36'sb10111001011010000100000110111111011;
        end
        2113: begin
            cosine_reg0 <= 36'sb10110000011100111000011000000100010;
            sine_reg0   <= 36'sb10111001011110011001010101011000011;
        end
        2114: begin
            cosine_reg0 <= 36'sb10110000011000010100111110101100010;
            sine_reg0   <= 36'sb10111001100010101110011100100111110;
        end
        2115: begin
            cosine_reg0 <= 36'sb10110000010011110001011110100001000;
            sine_reg0   <= 36'sb10111001100111000011011100101101011;
        end
        2116: begin
            cosine_reg0 <= 36'sb10110000001111001101110111100010110;
            sine_reg0   <= 36'sb10111001101011011000010101101000111;
        end
        2117: begin
            cosine_reg0 <= 36'sb10110000001010101010001001110001101;
            sine_reg0   <= 36'sb10111001101111101101000111011010011;
        end
        2118: begin
            cosine_reg0 <= 36'sb10110000000110000110010101001101111;
            sine_reg0   <= 36'sb10111001110100000001110010000001100;
        end
        2119: begin
            cosine_reg0 <= 36'sb10110000000001100010011001110111101;
            sine_reg0   <= 36'sb10111001111000010110010101011110001;
        end
        2120: begin
            cosine_reg0 <= 36'sb10101111111100111110010111101111001;
            sine_reg0   <= 36'sb10111001111100101010110001110000001;
        end
        2121: begin
            cosine_reg0 <= 36'sb10101111111000011010001110110100011;
            sine_reg0   <= 36'sb10111010000000111111000110110111011;
        end
        2122: begin
            cosine_reg0 <= 36'sb10101111110011110101111111000111101;
            sine_reg0   <= 36'sb10111010000101010011010100110011101;
        end
        2123: begin
            cosine_reg0 <= 36'sb10101111101111010001101000101001001;
            sine_reg0   <= 36'sb10111010001001100111011011100100101;
        end
        2124: begin
            cosine_reg0 <= 36'sb10101111101010101101001011011001001;
            sine_reg0   <= 36'sb10111010001101111011011011001010100;
        end
        2125: begin
            cosine_reg0 <= 36'sb10101111100110001000100111010111100;
            sine_reg0   <= 36'sb10111010010010001111010011100100110;
        end
        2126: begin
            cosine_reg0 <= 36'sb10101111100001100011111100100100110;
            sine_reg0   <= 36'sb10111010010110100011000100110011011;
        end
        2127: begin
            cosine_reg0 <= 36'sb10101111011100111111001011000000111;
            sine_reg0   <= 36'sb10111010011010110110101110110110010;
        end
        2128: begin
            cosine_reg0 <= 36'sb10101111011000011010010010101100000;
            sine_reg0   <= 36'sb10111010011111001010010001101101001;
        end
        2129: begin
            cosine_reg0 <= 36'sb10101111010011110101010011100110100;
            sine_reg0   <= 36'sb10111010100011011101101101011000000;
        end
        2130: begin
            cosine_reg0 <= 36'sb10101111001111010000001101110000011;
            sine_reg0   <= 36'sb10111010100111110001000001110110011;
        end
        2131: begin
            cosine_reg0 <= 36'sb10101111001010101011000001001001111;
            sine_reg0   <= 36'sb10111010101100000100001111001000011;
        end
        2132: begin
            cosine_reg0 <= 36'sb10101111000110000101101101110011001;
            sine_reg0   <= 36'sb10111010110000010111010101001101110;
        end
        2133: begin
            cosine_reg0 <= 36'sb10101111000001100000010011101100100;
            sine_reg0   <= 36'sb10111010110100101010010100000110010;
        end
        2134: begin
            cosine_reg0 <= 36'sb10101110111100111010110010110101111;
            sine_reg0   <= 36'sb10111010111000111101001011110001111;
        end
        2135: begin
            cosine_reg0 <= 36'sb10101110111000010101001011001111101;
            sine_reg0   <= 36'sb10111010111101001111111100010000010;
        end
        2136: begin
            cosine_reg0 <= 36'sb10101110110011101111011100111001111;
            sine_reg0   <= 36'sb10111011000001100010100101100001011;
        end
        2137: begin
            cosine_reg0 <= 36'sb10101110101111001001100111110100110;
            sine_reg0   <= 36'sb10111011000101110101000111100101001;
        end
        2138: begin
            cosine_reg0 <= 36'sb10101110101010100011101100000000100;
            sine_reg0   <= 36'sb10111011001010000111100010011011001;
        end
        2139: begin
            cosine_reg0 <= 36'sb10101110100101111101101001011101011;
            sine_reg0   <= 36'sb10111011001110011001110110000011011;
        end
        2140: begin
            cosine_reg0 <= 36'sb10101110100001010111100000001011011;
            sine_reg0   <= 36'sb10111011010010101100000010011101110;
        end
        2141: begin
            cosine_reg0 <= 36'sb10101110011100110001010000001010110;
            sine_reg0   <= 36'sb10111011010110111110000111101001111;
        end
        2142: begin
            cosine_reg0 <= 36'sb10101110011000001010111001011011110;
            sine_reg0   <= 36'sb10111011011011010000000101100111110;
        end
        2143: begin
            cosine_reg0 <= 36'sb10101110010011100100011011111110100;
            sine_reg0   <= 36'sb10111011011111100001111100010111010;
        end
        2144: begin
            cosine_reg0 <= 36'sb10101110001110111101110111110011001;
            sine_reg0   <= 36'sb10111011100011110011101011111000000;
        end
        2145: begin
            cosine_reg0 <= 36'sb10101110001010010111001100111001110;
            sine_reg0   <= 36'sb10111011101000000101010100001010000;
        end
        2146: begin
            cosine_reg0 <= 36'sb10101110000101110000011011010010110;
            sine_reg0   <= 36'sb10111011101100010110110101001101001;
        end
        2147: begin
            cosine_reg0 <= 36'sb10101110000001001001100010111110010;
            sine_reg0   <= 36'sb10111011110000101000001111000001001;
        end
        2148: begin
            cosine_reg0 <= 36'sb10101101111100100010100011111100010;
            sine_reg0   <= 36'sb10111011110100111001100001100101110;
        end
        2149: begin
            cosine_reg0 <= 36'sb10101101110111111011011110001101001;
            sine_reg0   <= 36'sb10111011111001001010101100111011000;
        end
        2150: begin
            cosine_reg0 <= 36'sb10101101110011010100010001110001000;
            sine_reg0   <= 36'sb10111011111101011011110001000000101;
        end
        2151: begin
            cosine_reg0 <= 36'sb10101101101110101100111110101000000;
            sine_reg0   <= 36'sb10111100000001101100101101110110100;
        end
        2152: begin
            cosine_reg0 <= 36'sb10101101101010000101100100110010011;
            sine_reg0   <= 36'sb10111100000101111101100011011100011;
        end
        2153: begin
            cosine_reg0 <= 36'sb10101101100101011110000100010000010;
            sine_reg0   <= 36'sb10111100001010001110010001110010010;
        end
        2154: begin
            cosine_reg0 <= 36'sb10101101100000110110011101000001111;
            sine_reg0   <= 36'sb10111100001110011110111000110111110;
        end
        2155: begin
            cosine_reg0 <= 36'sb10101101011100001110101111000111010;
            sine_reg0   <= 36'sb10111100010010101111011000101101000;
        end
        2156: begin
            cosine_reg0 <= 36'sb10101101010111100110111010100000110;
            sine_reg0   <= 36'sb10111100010110111111110001010001100;
        end
        2157: begin
            cosine_reg0 <= 36'sb10101101010010111110111111001110100;
            sine_reg0   <= 36'sb10111100011011010000000010100101010;
        end
        2158: begin
            cosine_reg0 <= 36'sb10101101001110010110111101010000101;
            sine_reg0   <= 36'sb10111100011111100000001100101000001;
        end
        2159: begin
            cosine_reg0 <= 36'sb10101101001001101110110100100111011;
            sine_reg0   <= 36'sb10111100100011110000001111011001111;
        end
        2160: begin
            cosine_reg0 <= 36'sb10101101000101000110100101010010111;
            sine_reg0   <= 36'sb10111100101000000000001010111010011;
        end
        2161: begin
            cosine_reg0 <= 36'sb10101101000000011110001111010011010;
            sine_reg0   <= 36'sb10111100101100001111111111001001100;
        end
        2162: begin
            cosine_reg0 <= 36'sb10101100111011110101110010101000110;
            sine_reg0   <= 36'sb10111100110000011111101100000111000;
        end
        2163: begin
            cosine_reg0 <= 36'sb10101100110111001101001111010011101;
            sine_reg0   <= 36'sb10111100110100101111010001110010110;
        end
        2164: begin
            cosine_reg0 <= 36'sb10101100110010100100100101010100000;
            sine_reg0   <= 36'sb10111100111000111110110000001100101;
        end
        2165: begin
            cosine_reg0 <= 36'sb10101100101101111011110100101010000;
            sine_reg0   <= 36'sb10111100111101001110000111010100100;
        end
        2166: begin
            cosine_reg0 <= 36'sb10101100101001010010111101010101110;
            sine_reg0   <= 36'sb10111101000001011101010111001010001;
        end
        2167: begin
            cosine_reg0 <= 36'sb10101100100100101001111111010111101;
            sine_reg0   <= 36'sb10111101000101101100011111101101010;
        end
        2168: begin
            cosine_reg0 <= 36'sb10101100100000000000111010101111101;
            sine_reg0   <= 36'sb10111101001001111011100000111101111;
        end
        2169: begin
            cosine_reg0 <= 36'sb10101100011011010111101111011110000;
            sine_reg0   <= 36'sb10111101001110001010011010111011110;
        end
        2170: begin
            cosine_reg0 <= 36'sb10101100010110101110011101100011000;
            sine_reg0   <= 36'sb10111101010010011001001101100110111;
        end
        2171: begin
            cosine_reg0 <= 36'sb10101100010010000101000100111110101;
            sine_reg0   <= 36'sb10111101010110100111111000111110110;
        end
        2172: begin
            cosine_reg0 <= 36'sb10101100001101011011100101110001010;
            sine_reg0   <= 36'sb10111101011010110110011101000011100;
        end
        2173: begin
            cosine_reg0 <= 36'sb10101100001000110001111111111011000;
            sine_reg0   <= 36'sb10111101011111000100111001110101000;
        end
        2174: begin
            cosine_reg0 <= 36'sb10101100000100001000010011011011111;
            sine_reg0   <= 36'sb10111101100011010011001111010010110;
        end
        2175: begin
            cosine_reg0 <= 36'sb10101011111111011110100000010100010;
            sine_reg0   <= 36'sb10111101100111100001011101011101000;
        end
        2176: begin
            cosine_reg0 <= 36'sb10101011111010110100100110100100011;
            sine_reg0   <= 36'sb10111101101011101111100100010011010;
        end
        2177: begin
            cosine_reg0 <= 36'sb10101011110110001010100110001100001;
            sine_reg0   <= 36'sb10111101101111111101100011110101100;
        end
        2178: begin
            cosine_reg0 <= 36'sb10101011110001100000011111001100000;
            sine_reg0   <= 36'sb10111101110100001011011100000011101;
        end
        2179: begin
            cosine_reg0 <= 36'sb10101011101100110110010001100100000;
            sine_reg0   <= 36'sb10111101111000011001001100111101010;
        end
        2180: begin
            cosine_reg0 <= 36'sb10101011101000001011111101010100010;
            sine_reg0   <= 36'sb10111101111100100110110110100010100;
        end
        2181: begin
            cosine_reg0 <= 36'sb10101011100011100001100010011101001;
            sine_reg0   <= 36'sb10111110000000110100011000110011000;
        end
        2182: begin
            cosine_reg0 <= 36'sb10101011011110110111000000111110110;
            sine_reg0   <= 36'sb10111110000101000001110011101110110;
        end
        2183: begin
            cosine_reg0 <= 36'sb10101011011010001100011000111001001;
            sine_reg0   <= 36'sb10111110001001001111000111010101100;
        end
        2184: begin
            cosine_reg0 <= 36'sb10101011010101100001101010001100101;
            sine_reg0   <= 36'sb10111110001101011100010011100111000;
        end
        2185: begin
            cosine_reg0 <= 36'sb10101011010000110110110100111001011;
            sine_reg0   <= 36'sb10111110010001101001011000100011010;
        end
        2186: begin
            cosine_reg0 <= 36'sb10101011001100001011111000111111101;
            sine_reg0   <= 36'sb10111110010101110110010110001001111;
        end
        2187: begin
            cosine_reg0 <= 36'sb10101011000111100000110110011111011;
            sine_reg0   <= 36'sb10111110011010000011001100011011000;
        end
        2188: begin
            cosine_reg0 <= 36'sb10101011000010110101101101011000111;
            sine_reg0   <= 36'sb10111110011110001111111011010110010;
        end
        2189: begin
            cosine_reg0 <= 36'sb10101010111110001010011101101100100;
            sine_reg0   <= 36'sb10111110100010011100100010111011101;
        end
        2190: begin
            cosine_reg0 <= 36'sb10101010111001011111000111011010001;
            sine_reg0   <= 36'sb10111110100110101001000011001010110;
        end
        2191: begin
            cosine_reg0 <= 36'sb10101010110100110011101010100010001;
            sine_reg0   <= 36'sb10111110101010110101011100000011101;
        end
        2192: begin
            cosine_reg0 <= 36'sb10101010110000001000000111000100101;
            sine_reg0   <= 36'sb10111110101111000001101101100110000;
        end
        2193: begin
            cosine_reg0 <= 36'sb10101010101011011100011101000001111;
            sine_reg0   <= 36'sb10111110110011001101110111110001110;
        end
        2194: begin
            cosine_reg0 <= 36'sb10101010100110110000101100011001111;
            sine_reg0   <= 36'sb10111110110111011001111010100110110;
        end
        2195: begin
            cosine_reg0 <= 36'sb10101010100010000100110101001101000;
            sine_reg0   <= 36'sb10111110111011100101110110000100111;
        end
        2196: begin
            cosine_reg0 <= 36'sb10101010011101011000110111011011011;
            sine_reg0   <= 36'sb10111110111111110001101010001011111;
        end
        2197: begin
            cosine_reg0 <= 36'sb10101010011000101100110011000101001;
            sine_reg0   <= 36'sb10111111000011111101010110111011100;
        end
        2198: begin
            cosine_reg0 <= 36'sb10101010010100000000101000001010011;
            sine_reg0   <= 36'sb10111111001000001000111100010011110;
        end
        2199: begin
            cosine_reg0 <= 36'sb10101010001111010100010110101011100;
            sine_reg0   <= 36'sb10111111001100010100011010010100100;
        end
        2200: begin
            cosine_reg0 <= 36'sb10101010001010100111111110101000101;
            sine_reg0   <= 36'sb10111111010000011111110000111101011;
        end
        2201: begin
            cosine_reg0 <= 36'sb10101010000101111011100000000001110;
            sine_reg0   <= 36'sb10111111010100101011000000001110100;
        end
        2202: begin
            cosine_reg0 <= 36'sb10101010000001001110111010110111010;
            sine_reg0   <= 36'sb10111111011000110110001000000111011;
        end
        2203: begin
            cosine_reg0 <= 36'sb10101001111100100010001111001001010;
            sine_reg0   <= 36'sb10111111011101000001001000101000001;
        end
        2204: begin
            cosine_reg0 <= 36'sb10101001110111110101011100111000000;
            sine_reg0   <= 36'sb10111111100001001100000001110000100;
        end
        2205: begin
            cosine_reg0 <= 36'sb10101001110011001000100100000011100;
            sine_reg0   <= 36'sb10111111100101010110110011100000010;
        end
        2206: begin
            cosine_reg0 <= 36'sb10101001101110011011100100101100000;
            sine_reg0   <= 36'sb10111111101001100001011101110111010;
        end
        2207: begin
            cosine_reg0 <= 36'sb10101001101001101110011110110001111;
            sine_reg0   <= 36'sb10111111101101101100000000110101100;
        end
        2208: begin
            cosine_reg0 <= 36'sb10101001100101000001010010010101000;
            sine_reg0   <= 36'sb10111111110001110110011100011010101;
        end
        2209: begin
            cosine_reg0 <= 36'sb10101001100000010011111111010101110;
            sine_reg0   <= 36'sb10111111110110000000110000100110101;
        end
        2210: begin
            cosine_reg0 <= 36'sb10101001011011100110100101110100011;
            sine_reg0   <= 36'sb10111111111010001010111101011001010;
        end
        2211: begin
            cosine_reg0 <= 36'sb10101001010110111001000101110000110;
            sine_reg0   <= 36'sb10111111111110010101000010110010010;
        end
        2212: begin
            cosine_reg0 <= 36'sb10101001010010001011011111001011011;
            sine_reg0   <= 36'sb11000000000010011111000000110001101;
        end
        2213: begin
            cosine_reg0 <= 36'sb10101001001101011101110010000100011;
            sine_reg0   <= 36'sb11000000000110101000110111010111010;
        end
        2214: begin
            cosine_reg0 <= 36'sb10101001001000101111111110011011110;
            sine_reg0   <= 36'sb11000000001010110010100110100010111;
        end
        2215: begin
            cosine_reg0 <= 36'sb10101001000100000010000100010001110;
            sine_reg0   <= 36'sb11000000001110111100001110010100010;
        end
        2216: begin
            cosine_reg0 <= 36'sb10101000111111010100000011100110110;
            sine_reg0   <= 36'sb11000000010011000101101110101011011;
        end
        2217: begin
            cosine_reg0 <= 36'sb10101000111010100101111100011010101;
            sine_reg0   <= 36'sb11000000010111001111000111101000000;
        end
        2218: begin
            cosine_reg0 <= 36'sb10101000110101110111101110101101111;
            sine_reg0   <= 36'sb11000000011011011000011001001010000;
        end
        2219: begin
            cosine_reg0 <= 36'sb10101000110001001001011010100000100;
            sine_reg0   <= 36'sb11000000011111100001100011010001001;
        end
        2220: begin
            cosine_reg0 <= 36'sb10101000101100011010111111110010101;
            sine_reg0   <= 36'sb11000000100011101010100101111101011;
        end
        2221: begin
            cosine_reg0 <= 36'sb10101000100111101100011110100100100;
            sine_reg0   <= 36'sb11000000100111110011100001001110100;
        end
        2222: begin
            cosine_reg0 <= 36'sb10101000100010111101110110110110011;
            sine_reg0   <= 36'sb11000000101011111100010101000100011;
        end
        2223: begin
            cosine_reg0 <= 36'sb10101000011110001111001000101000011;
            sine_reg0   <= 36'sb11000000110000000101000001011110110;
        end
        2224: begin
            cosine_reg0 <= 36'sb10101000011001100000010011111010110;
            sine_reg0   <= 36'sb11000000110100001101100110011101101;
        end
        2225: begin
            cosine_reg0 <= 36'sb10101000010100110001011000101101100;
            sine_reg0   <= 36'sb11000000111000010110000100000000101;
        end
        2226: begin
            cosine_reg0 <= 36'sb10101000010000000010010111000001000;
            sine_reg0   <= 36'sb11000000111100011110011010000111110;
        end
        2227: begin
            cosine_reg0 <= 36'sb10101000001011010011001110110101011;
            sine_reg0   <= 36'sb11000001000000100110101000110010111;
        end
        2228: begin
            cosine_reg0 <= 36'sb10101000000110100100000000001010110;
            sine_reg0   <= 36'sb11000001000100101110110000000001110;
        end
        2229: begin
            cosine_reg0 <= 36'sb10101000000001110100101011000001011;
            sine_reg0   <= 36'sb11000001001000110110101111110100001;
        end
        2230: begin
            cosine_reg0 <= 36'sb10100111111101000101001111011001011;
            sine_reg0   <= 36'sb11000001001100111110101000001010000;
        end
        2231: begin
            cosine_reg0 <= 36'sb10100111111000010101101101010011000;
            sine_reg0   <= 36'sb11000001010001000110011001000011010;
        end
        2232: begin
            cosine_reg0 <= 36'sb10100111110011100110000100101110011;
            sine_reg0   <= 36'sb11000001010101001110000010011111101;
        end
        2233: begin
            cosine_reg0 <= 36'sb10100111101110110110010101101011101;
            sine_reg0   <= 36'sb11000001011001010101100100011110111;
        end
        2234: begin
            cosine_reg0 <= 36'sb10100111101010000110100000001011001;
            sine_reg0   <= 36'sb11000001011101011100111111000001000;
        end
        2235: begin
            cosine_reg0 <= 36'sb10100111100101010110100100001100111;
            sine_reg0   <= 36'sb11000001100001100100010010000101110;
        end
        2236: begin
            cosine_reg0 <= 36'sb10100111100000100110100001110001001;
            sine_reg0   <= 36'sb11000001100101101011011101101101000;
        end
        2237: begin
            cosine_reg0 <= 36'sb10100111011011110110011000111000001;
            sine_reg0   <= 36'sb11000001101001110010100001110110101;
        end
        2238: begin
            cosine_reg0 <= 36'sb10100111010111000110001001100010000;
            sine_reg0   <= 36'sb11000001101101111001011110100010011;
        end
        2239: begin
            cosine_reg0 <= 36'sb10100111010010010101110011101110111;
            sine_reg0   <= 36'sb11000001110010000000010011110000010;
        end
        2240: begin
            cosine_reg0 <= 36'sb10100111001101100101010111011111000;
            sine_reg0   <= 36'sb11000001110110000111000001011111111;
        end
        2241: begin
            cosine_reg0 <= 36'sb10100111001000110100110100110010101;
            sine_reg0   <= 36'sb11000001111010001101100111110001010;
        end
        2242: begin
            cosine_reg0 <= 36'sb10100111000100000100001011101001110;
            sine_reg0   <= 36'sb11000001111110010100000110100100010;
        end
        2243: begin
            cosine_reg0 <= 36'sb10100110111111010011011100000100110;
            sine_reg0   <= 36'sb11000010000010011010011101111000100;
        end
        2244: begin
            cosine_reg0 <= 36'sb10100110111010100010100110000011101;
            sine_reg0   <= 36'sb11000010000110100000101101101110000;
        end
        2245: begin
            cosine_reg0 <= 36'sb10100110110101110001101001100110110;
            sine_reg0   <= 36'sb11000010001010100110110110000100101;
        end
        2246: begin
            cosine_reg0 <= 36'sb10100110110001000000100110101110001;
            sine_reg0   <= 36'sb11000010001110101100110110111100010;
        end
        2247: begin
            cosine_reg0 <= 36'sb10100110101100001111011101011010000;
            sine_reg0   <= 36'sb11000010010010110010110000010100100;
        end
        2248: begin
            cosine_reg0 <= 36'sb10100110100111011110001101101010110;
            sine_reg0   <= 36'sb11000010010110111000100010001101011;
        end
        2249: begin
            cosine_reg0 <= 36'sb10100110100010101100110111100000010;
            sine_reg0   <= 36'sb11000010011010111110001100100110110;
        end
        2250: begin
            cosine_reg0 <= 36'sb10100110011101111011011010111010111;
            sine_reg0   <= 36'sb11000010011111000011101111100000011;
        end
        2251: begin
            cosine_reg0 <= 36'sb10100110011001001001110111111010101;
            sine_reg0   <= 36'sb11000010100011001001001010111010001;
        end
        2252: begin
            cosine_reg0 <= 36'sb10100110010100011000001110100000000;
            sine_reg0   <= 36'sb11000010100111001110011110110011110;
        end
        2253: begin
            cosine_reg0 <= 36'sb10100110001111100110011110101010111;
            sine_reg0   <= 36'sb11000010101011010011101011001101011;
        end
        2254: begin
            cosine_reg0 <= 36'sb10100110001010110100101000011011101;
            sine_reg0   <= 36'sb11000010101111011000110000000110100;
        end
        2255: begin
            cosine_reg0 <= 36'sb10100110000110000010101011110010011;
            sine_reg0   <= 36'sb11000010110011011101101101011111001;
        end
        2256: begin
            cosine_reg0 <= 36'sb10100110000001010000101000101111010;
            sine_reg0   <= 36'sb11000010110111100010100011010111010;
        end
        2257: begin
            cosine_reg0 <= 36'sb10100101111100011110011111010010101;
            sine_reg0   <= 36'sb11000010111011100111010001101110011;
        end
        2258: begin
            cosine_reg0 <= 36'sb10100101110111101100001111011100011;
            sine_reg0   <= 36'sb11000010111111101011111000100100101;
        end
        2259: begin
            cosine_reg0 <= 36'sb10100101110010111001111001001101000;
            sine_reg0   <= 36'sb11000011000011110000010111111001110;
        end
        2260: begin
            cosine_reg0 <= 36'sb10100101101110000111011100100100011;
            sine_reg0   <= 36'sb11000011000111110100101111101101100;
        end
        2261: begin
            cosine_reg0 <= 36'sb10100101101001010100111001100011000;
            sine_reg0   <= 36'sb11000011001011111000111111111111111;
        end
        2262: begin
            cosine_reg0 <= 36'sb10100101100100100010010000001000111;
            sine_reg0   <= 36'sb11000011001111111101001000110000101;
        end
        2263: begin
            cosine_reg0 <= 36'sb10100101011111101111100000010110001;
            sine_reg0   <= 36'sb11000011010100000001001001111111101;
        end
        2264: begin
            cosine_reg0 <= 36'sb10100101011010111100101010001011001;
            sine_reg0   <= 36'sb11000011011000000101000011101100110;
        end
        2265: begin
            cosine_reg0 <= 36'sb10100101010110001001101101101000000;
            sine_reg0   <= 36'sb11000011011100001000110101110111110;
        end
        2266: begin
            cosine_reg0 <= 36'sb10100101010001010110101010101100110;
            sine_reg0   <= 36'sb11000011100000001100100000100000100;
        end
        2267: begin
            cosine_reg0 <= 36'sb10100101001100100011100001011001111;
            sine_reg0   <= 36'sb11000011100100010000000011100111000;
        end
        2268: begin
            cosine_reg0 <= 36'sb10100101000111110000010001101111011;
            sine_reg0   <= 36'sb11000011101000010011011111001010110;
        end
        2269: begin
            cosine_reg0 <= 36'sb10100101000010111100111011101101011;
            sine_reg0   <= 36'sb11000011101100010110110011001100000;
        end
        2270: begin
            cosine_reg0 <= 36'sb10100100111110001001011111010100001;
            sine_reg0   <= 36'sb11000011110000011001111111101010010;
        end
        2271: begin
            cosine_reg0 <= 36'sb10100100111001010101111100100011111;
            sine_reg0   <= 36'sb11000011110100011101000100100101101;
        end
        2272: begin
            cosine_reg0 <= 36'sb10100100110100100010010011011100110;
            sine_reg0   <= 36'sb11000011111000100000000001111101110;
        end
        2273: begin
            cosine_reg0 <= 36'sb10100100101111101110100011111111000;
            sine_reg0   <= 36'sb11000011111100100010110111110010100;
        end
        2274: begin
            cosine_reg0 <= 36'sb10100100101010111010101110001010101;
            sine_reg0   <= 36'sb11000100000000100101100110000011111;
        end
        2275: begin
            cosine_reg0 <= 36'sb10100100100110000110110010000000001;
            sine_reg0   <= 36'sb11000100000100101000001100110001101;
        end
        2276: begin
            cosine_reg0 <= 36'sb10100100100001010010101111011111011;
            sine_reg0   <= 36'sb11000100001000101010101011111011100;
        end
        2277: begin
            cosine_reg0 <= 36'sb10100100011100011110100110101000110;
            sine_reg0   <= 36'sb11000100001100101101000011100001100;
        end
        2278: begin
            cosine_reg0 <= 36'sb10100100010111101010010111011100010;
            sine_reg0   <= 36'sb11000100010000101111010011100011011;
        end
        2279: begin
            cosine_reg0 <= 36'sb10100100010010110110000001111010010;
            sine_reg0   <= 36'sb11000100010100110001011100000001000;
        end
        2280: begin
            cosine_reg0 <= 36'sb10100100001110000001100110000011000;
            sine_reg0   <= 36'sb11000100011000110011011100111010001;
        end
        2281: begin
            cosine_reg0 <= 36'sb10100100001001001101000011110110011;
            sine_reg0   <= 36'sb11000100011100110101010110001110110;
        end
        2282: begin
            cosine_reg0 <= 36'sb10100100000100011000011011010100111;
            sine_reg0   <= 36'sb11000100100000110111000111111110110;
        end
        2283: begin
            cosine_reg0 <= 36'sb10100011111111100011101100011110011;
            sine_reg0   <= 36'sb11000100100100111000110010001001110;
        end
        2284: begin
            cosine_reg0 <= 36'sb10100011111010101110110111010011011;
            sine_reg0   <= 36'sb11000100101000111010010100101111110;
        end
        2285: begin
            cosine_reg0 <= 36'sb10100011110101111001111011110100000;
            sine_reg0   <= 36'sb11000100101100111011101111110000101;
        end
        2286: begin
            cosine_reg0 <= 36'sb10100011110001000100111010000000010;
            sine_reg0   <= 36'sb11000100110000111101000011001100000;
        end
        2287: begin
            cosine_reg0 <= 36'sb10100011101100001111110001111000011;
            sine_reg0   <= 36'sb11000100110100111110001111000010000;
        end
        2288: begin
            cosine_reg0 <= 36'sb10100011100111011010100011011100101;
            sine_reg0   <= 36'sb11000100111000111111010011010010011;
        end
        2289: begin
            cosine_reg0 <= 36'sb10100011100010100101001110101101010;
            sine_reg0   <= 36'sb11000100111101000000001111111100111;
        end
        2290: begin
            cosine_reg0 <= 36'sb10100011011101101111110011101010011;
            sine_reg0   <= 36'sb11000101000001000001000101000001011;
        end
        2291: begin
            cosine_reg0 <= 36'sb10100011011000111010010010010100001;
            sine_reg0   <= 36'sb11000101000101000001110010011111111;
        end
        2292: begin
            cosine_reg0 <= 36'sb10100011010100000100101010101010101;
            sine_reg0   <= 36'sb11000101001001000010011000011000000;
        end
        2293: begin
            cosine_reg0 <= 36'sb10100011001111001110111100101110010;
            sine_reg0   <= 36'sb11000101001101000010110110101001110;
        end
        2294: begin
            cosine_reg0 <= 36'sb10100011001010011001001000011111001;
            sine_reg0   <= 36'sb11000101010001000011001101010100111;
        end
        2295: begin
            cosine_reg0 <= 36'sb10100011000101100011001101111101011;
            sine_reg0   <= 36'sb11000101010101000011011100011001011;
        end
        2296: begin
            cosine_reg0 <= 36'sb10100011000000101101001101001001010;
            sine_reg0   <= 36'sb11000101011001000011100011110110111;
        end
        2297: begin
            cosine_reg0 <= 36'sb10100010111011110111000110000010111;
            sine_reg0   <= 36'sb11000101011101000011100011101101011;
        end
        2298: begin
            cosine_reg0 <= 36'sb10100010110111000000111000101010100;
            sine_reg0   <= 36'sb11000101100001000011011011111100101;
        end
        2299: begin
            cosine_reg0 <= 36'sb10100010110010001010100101000000011;
            sine_reg0   <= 36'sb11000101100101000011001100100100100;
        end
        2300: begin
            cosine_reg0 <= 36'sb10100010101101010100001011000100100;
            sine_reg0   <= 36'sb11000101101001000010110101100101000;
        end
        2301: begin
            cosine_reg0 <= 36'sb10100010101000011101101010110111001;
            sine_reg0   <= 36'sb11000101101101000010010110111101110;
        end
        2302: begin
            cosine_reg0 <= 36'sb10100010100011100111000100011000100;
            sine_reg0   <= 36'sb11000101110001000001110000101110110;
        end
        2303: begin
            cosine_reg0 <= 36'sb10100010011110110000010111101000111;
            sine_reg0   <= 36'sb11000101110101000001000010110111110;
        end
        2304: begin
            cosine_reg0 <= 36'sb10100010011001111001100100101000010;
            sine_reg0   <= 36'sb11000101111001000000001101011000100;
        end
        2305: begin
            cosine_reg0 <= 36'sb10100010010101000010101011010110111;
            sine_reg0   <= 36'sb11000101111100111111010000010001001;
        end
        2306: begin
            cosine_reg0 <= 36'sb10100010010000001011101011110101000;
            sine_reg0   <= 36'sb11000110000000111110001011100001010;
        end
        2307: begin
            cosine_reg0 <= 36'sb10100010001011010100100110000010111;
            sine_reg0   <= 36'sb11000110000100111100111111001000111;
        end
        2308: begin
            cosine_reg0 <= 36'sb10100010000110011101011010000000100;
            sine_reg0   <= 36'sb11000110001000111011101011000111110;
        end
        2309: begin
            cosine_reg0 <= 36'sb10100010000001100110000111101110001;
            sine_reg0   <= 36'sb11000110001100111010001111011101101;
        end
        2310: begin
            cosine_reg0 <= 36'sb10100001111100101110101111001100000;
            sine_reg0   <= 36'sb11000110010000111000101100001010101;
        end
        2311: begin
            cosine_reg0 <= 36'sb10100001110111110111010000011010011;
            sine_reg0   <= 36'sb11000110010100110111000001001110010;
        end
        2312: begin
            cosine_reg0 <= 36'sb10100001110010111111101011011001010;
            sine_reg0   <= 36'sb11000110011000110101001110101000101;
        end
        2313: begin
            cosine_reg0 <= 36'sb10100001101110001000000000001000111;
            sine_reg0   <= 36'sb11000110011100110011010100011001100;
        end
        2314: begin
            cosine_reg0 <= 36'sb10100001101001010000001110101001101;
            sine_reg0   <= 36'sb11000110100000110001010010100000110;
        end
        2315: begin
            cosine_reg0 <= 36'sb10100001100100011000010110111011011;
            sine_reg0   <= 36'sb11000110100100101111001000111110001;
        end
        2316: begin
            cosine_reg0 <= 36'sb10100001011111100000011000111110100;
            sine_reg0   <= 36'sb11000110101000101100110111110001100;
        end
        2317: begin
            cosine_reg0 <= 36'sb10100001011010101000010100110011010;
            sine_reg0   <= 36'sb11000110101100101010011110111010111;
        end
        2318: begin
            cosine_reg0 <= 36'sb10100001010101110000001010011001101;
            sine_reg0   <= 36'sb11000110110000100111111110011001111;
        end
        2319: begin
            cosine_reg0 <= 36'sb10100001010000110111111001110010000;
            sine_reg0   <= 36'sb11000110110100100101010110001110100;
        end
        2320: begin
            cosine_reg0 <= 36'sb10100001001011111111100010111100011;
            sine_reg0   <= 36'sb11000110111000100010100110011000101;
        end
        2321: begin
            cosine_reg0 <= 36'sb10100001000111000111000101111001001;
            sine_reg0   <= 36'sb11000110111100011111101110111000000;
        end
        2322: begin
            cosine_reg0 <= 36'sb10100001000010001110100010101000010;
            sine_reg0   <= 36'sb11000111000000011100101111101100011;
        end
        2323: begin
            cosine_reg0 <= 36'sb10100000111101010101111001001010001;
            sine_reg0   <= 36'sb11000111000100011001101000110101111;
        end
        2324: begin
            cosine_reg0 <= 36'sb10100000111000011101001001011110110;
            sine_reg0   <= 36'sb11000111001000010110011010010100001;
        end
        2325: begin
            cosine_reg0 <= 36'sb10100000110011100100010011100110100;
            sine_reg0   <= 36'sb11000111001100010011000100000111000;
        end
        2326: begin
            cosine_reg0 <= 36'sb10100000101110101011010111100001100;
            sine_reg0   <= 36'sb11000111010000001111100110001110011;
        end
        2327: begin
            cosine_reg0 <= 36'sb10100000101001110010010101001111111;
            sine_reg0   <= 36'sb11000111010100001100000000101010001;
        end
        2328: begin
            cosine_reg0 <= 36'sb10100000100100111001001100110001111;
            sine_reg0   <= 36'sb11000111011000001000010011011010001;
        end
        2329: begin
            cosine_reg0 <= 36'sb10100000011111111111111110000111101;
            sine_reg0   <= 36'sb11000111011100000100011110011110010;
        end
        2330: begin
            cosine_reg0 <= 36'sb10100000011011000110101001010001011;
            sine_reg0   <= 36'sb11000111100000000000100001110110001;
        end
        2331: begin
            cosine_reg0 <= 36'sb10100000010110001101001110001111010;
            sine_reg0   <= 36'sb11000111100011111100011101100001111;
        end
        2332: begin
            cosine_reg0 <= 36'sb10100000010001010011101101000001101;
            sine_reg0   <= 36'sb11000111100111111000010001100001001;
        end
        2333: begin
            cosine_reg0 <= 36'sb10100000001100011010000101101000011;
            sine_reg0   <= 36'sb11000111101011110011111101110011111;
        end
        2334: begin
            cosine_reg0 <= 36'sb10100000000111100000011000000100000;
            sine_reg0   <= 36'sb11000111101111101111100010011010000;
        end
        2335: begin
            cosine_reg0 <= 36'sb10100000000010100110100100010100100;
            sine_reg0   <= 36'sb11000111110011101010111111010011010;
        end
        2336: begin
            cosine_reg0 <= 36'sb10011111111101101100101010011010001;
            sine_reg0   <= 36'sb11000111110111100110010100011111011;
        end
        2337: begin
            cosine_reg0 <= 36'sb10011111111000110010101010010101000;
            sine_reg0   <= 36'sb11000111111011100001100001111110011;
        end
        2338: begin
            cosine_reg0 <= 36'sb10011111110011111000100100000101011;
            sine_reg0   <= 36'sb11000111111111011100100111110000001;
        end
        2339: begin
            cosine_reg0 <= 36'sb10011111101110111110010111101011100;
            sine_reg0   <= 36'sb11001000000011010111100101110100011;
        end
        2340: begin
            cosine_reg0 <= 36'sb10011111101010000100000101000111100;
            sine_reg0   <= 36'sb11001000000111010010011100001011001;
        end
        2341: begin
            cosine_reg0 <= 36'sb10011111100101001001101100011001100;
            sine_reg0   <= 36'sb11001000001011001101001010110100000;
        end
        2342: begin
            cosine_reg0 <= 36'sb10011111100000001111001101100001110;
            sine_reg0   <= 36'sb11001000001111000111110001101111000;
        end
        2343: begin
            cosine_reg0 <= 36'sb10011111011011010100101000100000100;
            sine_reg0   <= 36'sb11001000010011000010010000111011111;
        end
        2344: begin
            cosine_reg0 <= 36'sb10011111010110011001111101010101111;
            sine_reg0   <= 36'sb11001000010110111100101000011010101;
        end
        2345: begin
            cosine_reg0 <= 36'sb10011111010001011111001100000010000;
            sine_reg0   <= 36'sb11001000011010110110111000001011000;
        end
        2346: begin
            cosine_reg0 <= 36'sb10011111001100100100010100100101010;
            sine_reg0   <= 36'sb11001000011110110001000000001100111;
        end
        2347: begin
            cosine_reg0 <= 36'sb10011111000111101001010110111111101;
            sine_reg0   <= 36'sb11001000100010101011000000100000000;
        end
        2348: begin
            cosine_reg0 <= 36'sb10011111000010101110010011010001011;
            sine_reg0   <= 36'sb11001000100110100100111001000100011;
        end
        2349: begin
            cosine_reg0 <= 36'sb10011110111101110011001001011010110;
            sine_reg0   <= 36'sb11001000101010011110101001111001110;
        end
        2350: begin
            cosine_reg0 <= 36'sb10011110111000110111111001011011110;
            sine_reg0   <= 36'sb11001000101110011000010011000000000;
        end
        2351: begin
            cosine_reg0 <= 36'sb10011110110011111100100011010100111;
            sine_reg0   <= 36'sb11001000110010010001110100010111000;
        end
        2352: begin
            cosine_reg0 <= 36'sb10011110101111000001000111000110001;
            sine_reg0   <= 36'sb11001000110110001011001101111110100;
        end
        2353: begin
            cosine_reg0 <= 36'sb10011110101010000101100100101111101;
            sine_reg0   <= 36'sb11001000111010000100011111110110100;
        end
        2354: begin
            cosine_reg0 <= 36'sb10011110100101001001111100010001110;
            sine_reg0   <= 36'sb11001000111101111101101001111110111;
        end
        2355: begin
            cosine_reg0 <= 36'sb10011110100000001110001101101100100;
            sine_reg0   <= 36'sb11001001000001110110101100010111010;
        end
        2356: begin
            cosine_reg0 <= 36'sb10011110011011010010011001000000010;
            sine_reg0   <= 36'sb11001001000101101111100110111111101;
        end
        2357: begin
            cosine_reg0 <= 36'sb10011110010110010110011110001101000;
            sine_reg0   <= 36'sb11001001001001101000011001110111111;
        end
        2358: begin
            cosine_reg0 <= 36'sb10011110010001011010011101010011001;
            sine_reg0   <= 36'sb11001001001101100001000100111111110;
        end
        2359: begin
            cosine_reg0 <= 36'sb10011110001100011110010110010010110;
            sine_reg0   <= 36'sb11001001010001011001101000010111010;
        end
        2360: begin
            cosine_reg0 <= 36'sb10011110000111100010001001001100000;
            sine_reg0   <= 36'sb11001001010101010010000011111110001;
        end
        2361: begin
            cosine_reg0 <= 36'sb10011110000010100101110101111111001;
            sine_reg0   <= 36'sb11001001011001001010010111110100001;
        end
        2362: begin
            cosine_reg0 <= 36'sb10011101111101101001011100101100010;
            sine_reg0   <= 36'sb11001001011101000010100011111001010;
        end
        2363: begin
            cosine_reg0 <= 36'sb10011101111000101100111101010011101;
            sine_reg0   <= 36'sb11001001100000111010101000001101011;
        end
        2364: begin
            cosine_reg0 <= 36'sb10011101110011110000010111110101100;
            sine_reg0   <= 36'sb11001001100100110010100100110000010;
        end
        2365: begin
            cosine_reg0 <= 36'sb10011101101110110011101100010001111;
            sine_reg0   <= 36'sb11001001101000101010011001100001110;
        end
        2366: begin
            cosine_reg0 <= 36'sb10011101101001110110111010101001010;
            sine_reg0   <= 36'sb11001001101100100010000110100001101;
        end
        2367: begin
            cosine_reg0 <= 36'sb10011101100100111010000010111011100;
            sine_reg0   <= 36'sb11001001110000011001101011110000000;
        end
        2368: begin
            cosine_reg0 <= 36'sb10011101011111111101000101001000111;
            sine_reg0   <= 36'sb11001001110100010001001001001100100;
        end
        2369: begin
            cosine_reg0 <= 36'sb10011101011011000000000001010001110;
            sine_reg0   <= 36'sb11001001111000001000011110110111000;
        end
        2370: begin
            cosine_reg0 <= 36'sb10011101010110000010110111010110010;
            sine_reg0   <= 36'sb11001001111011111111101100101111011;
        end
        2371: begin
            cosine_reg0 <= 36'sb10011101010001000101100111010110011;
            sine_reg0   <= 36'sb11001001111111110110110010110101101;
        end
        2372: begin
            cosine_reg0 <= 36'sb10011101001100001000010001010010101;
            sine_reg0   <= 36'sb11001010000011101101110001001001011;
        end
        2373: begin
            cosine_reg0 <= 36'sb10011101000111001010110101001010111;
            sine_reg0   <= 36'sb11001010000111100100100111101010100;
        end
        2374: begin
            cosine_reg0 <= 36'sb10011101000010001101010010111111100;
            sine_reg0   <= 36'sb11001010001011011011010110011001000;
        end
        2375: begin
            cosine_reg0 <= 36'sb10011100111101001111101010110000110;
            sine_reg0   <= 36'sb11001010001111010001111101010100101;
        end
        2376: begin
            cosine_reg0 <= 36'sb10011100111000010001111100011110101;
            sine_reg0   <= 36'sb11001010010011001000011100011101010;
        end
        2377: begin
            cosine_reg0 <= 36'sb10011100110011010100001000001001100;
            sine_reg0   <= 36'sb11001010010110111110110011110010110;
        end
        2378: begin
            cosine_reg0 <= 36'sb10011100101110010110001101110001011;
            sine_reg0   <= 36'sb11001010011010110101000011010100111;
        end
        2379: begin
            cosine_reg0 <= 36'sb10011100101001011000001101010110101;
            sine_reg0   <= 36'sb11001010011110101011001011000011101;
        end
        2380: begin
            cosine_reg0 <= 36'sb10011100100100011010000110111001011;
            sine_reg0   <= 36'sb11001010100010100001001010111110110;
        end
        2381: begin
            cosine_reg0 <= 36'sb10011100011111011011111010011001110;
            sine_reg0   <= 36'sb11001010100110010111000011000110001;
        end
        2382: begin
            cosine_reg0 <= 36'sb10011100011010011101100111111000000;
            sine_reg0   <= 36'sb11001010101010001100110011011001101;
        end
        2383: begin
            cosine_reg0 <= 36'sb10011100010101011111001111010100011;
            sine_reg0   <= 36'sb11001010101110000010011011111001001;
        end
        2384: begin
            cosine_reg0 <= 36'sb10011100010000100000110000101110111;
            sine_reg0   <= 36'sb11001010110001110111111100100100011;
        end
        2385: begin
            cosine_reg0 <= 36'sb10011100001011100010001100001000000;
            sine_reg0   <= 36'sb11001010110101101101010101011011010;
        end
        2386: begin
            cosine_reg0 <= 36'sb10011100000110100011100001011111101;
            sine_reg0   <= 36'sb11001010111001100010100110011101110;
        end
        2387: begin
            cosine_reg0 <= 36'sb10011100000001100100110000110110001;
            sine_reg0   <= 36'sb11001010111101010111101111101011100;
        end
        2388: begin
            cosine_reg0 <= 36'sb10011011111100100101111010001011110;
            sine_reg0   <= 36'sb11001011000001001100110001000100100;
        end
        2389: begin
            cosine_reg0 <= 36'sb10011011110111100110111101100000100;
            sine_reg0   <= 36'sb11001011000101000001101010101000101;
        end
        2390: begin
            cosine_reg0 <= 36'sb10011011110010100111111010110100101;
            sine_reg0   <= 36'sb11001011001000110110011100010111101;
        end
        2391: begin
            cosine_reg0 <= 36'sb10011011101101101000110010001000011;
            sine_reg0   <= 36'sb11001011001100101011000110010001011;
        end
        2392: begin
            cosine_reg0 <= 36'sb10011011101000101001100011011100000;
            sine_reg0   <= 36'sb11001011010000011111101000010101111;
        end
        2393: begin
            cosine_reg0 <= 36'sb10011011100011101010001110101111100;
            sine_reg0   <= 36'sb11001011010100010100000010100100110;
        end
        2394: begin
            cosine_reg0 <= 36'sb10011011011110101010110100000011010;
            sine_reg0   <= 36'sb11001011011000001000010100111110000;
        end
        2395: begin
            cosine_reg0 <= 36'sb10011011011001101011010011010111011;
            sine_reg0   <= 36'sb11001011011011111100011111100001011;
        end
        2396: begin
            cosine_reg0 <= 36'sb10011011010100101011101100101100000;
            sine_reg0   <= 36'sb11001011011111110000100010001110111;
        end
        2397: begin
            cosine_reg0 <= 36'sb10011011001111101100000000000001011;
            sine_reg0   <= 36'sb11001011100011100100011101000110010;
        end
        2398: begin
            cosine_reg0 <= 36'sb10011011001010101100001101010111110;
            sine_reg0   <= 36'sb11001011100111011000010000000111010;
        end
        2399: begin
            cosine_reg0 <= 36'sb10011011000101101100010100101111010;
            sine_reg0   <= 36'sb11001011101011001011111011010010000;
        end
        2400: begin
            cosine_reg0 <= 36'sb10011011000000101100010110001000001;
            sine_reg0   <= 36'sb11001011101110111111011110100110001;
        end
        2401: begin
            cosine_reg0 <= 36'sb10011010111011101100010001100010100;
            sine_reg0   <= 36'sb11001011110010110010111010000011101;
        end
        2402: begin
            cosine_reg0 <= 36'sb10011010110110101100000110111110101;
            sine_reg0   <= 36'sb11001011110110100110001101101010010;
        end
        2403: begin
            cosine_reg0 <= 36'sb10011010110001101011110110011100101;
            sine_reg0   <= 36'sb11001011111010011001011001011001111;
        end
        2404: begin
            cosine_reg0 <= 36'sb10011010101100101011011111111100101;
            sine_reg0   <= 36'sb11001011111110001100011101010010011;
        end
        2405: begin
            cosine_reg0 <= 36'sb10011010100111101011000011011111000;
            sine_reg0   <= 36'sb11001100000001111111011001010011101;
        end
        2406: begin
            cosine_reg0 <= 36'sb10011010100010101010100001000100000;
            sine_reg0   <= 36'sb11001100000101110010001101011101011;
        end
        2407: begin
            cosine_reg0 <= 36'sb10011010011101101001111000101011100;
            sine_reg0   <= 36'sb11001100001001100100111001101111101;
        end
        2408: begin
            cosine_reg0 <= 36'sb10011010011000101001001010010110000;
            sine_reg0   <= 36'sb11001100001101010111011110001010001;
        end
        2409: begin
            cosine_reg0 <= 36'sb10011010010011101000010110000011100;
            sine_reg0   <= 36'sb11001100010001001001111010101100110;
        end
        2410: begin
            cosine_reg0 <= 36'sb10011010001110100111011011110100010;
            sine_reg0   <= 36'sb11001100010100111100001111010111011;
        end
        2411: begin
            cosine_reg0 <= 36'sb10011010001001100110011011101000100;
            sine_reg0   <= 36'sb11001100011000101110011100001001110;
        end
        2412: begin
            cosine_reg0 <= 36'sb10011010000100100101010101100000011;
            sine_reg0   <= 36'sb11001100011100100000100001000100000;
        end
        2413: begin
            cosine_reg0 <= 36'sb10011001111111100100001001011100001;
            sine_reg0   <= 36'sb11001100100000010010011110000101101;
        end
        2414: begin
            cosine_reg0 <= 36'sb10011001111010100010110111011011111;
            sine_reg0   <= 36'sb11001100100100000100010011001110110;
        end
        2415: begin
            cosine_reg0 <= 36'sb10011001110101100001011111011111111;
            sine_reg0   <= 36'sb11001100100111110110000000011111001;
        end
        2416: begin
            cosine_reg0 <= 36'sb10011001110000100000000001101000011;
            sine_reg0   <= 36'sb11001100101011100111100101110110101;
        end
        2417: begin
            cosine_reg0 <= 36'sb10011001101011011110011101110101011;
            sine_reg0   <= 36'sb11001100101111011001000011010101001;
        end
        2418: begin
            cosine_reg0 <= 36'sb10011001100110011100110100000111010;
            sine_reg0   <= 36'sb11001100110011001010011000111010011;
        end
        2419: begin
            cosine_reg0 <= 36'sb10011001100001011011000100011110001;
            sine_reg0   <= 36'sb11001100110110111011100110100110011;
        end
        2420: begin
            cosine_reg0 <= 36'sb10011001011100011001001110111010001;
            sine_reg0   <= 36'sb11001100111010101100101100011000111;
        end
        2421: begin
            cosine_reg0 <= 36'sb10011001010111010111010011011011101;
            sine_reg0   <= 36'sb11001100111110011101101010010001110;
        end
        2422: begin
            cosine_reg0 <= 36'sb10011001010010010101010010000010101;
            sine_reg0   <= 36'sb11001101000010001110100000010000111;
        end
        2423: begin
            cosine_reg0 <= 36'sb10011001001101010011001010101111011;
            sine_reg0   <= 36'sb11001101000101111111001110010110001;
        end
        2424: begin
            cosine_reg0 <= 36'sb10011001001000010000111101100010010;
            sine_reg0   <= 36'sb11001101001001101111110100100001010;
        end
        2425: begin
            cosine_reg0 <= 36'sb10011001000011001110101010011011010;
            sine_reg0   <= 36'sb11001101001101100000010010110010010;
        end
        2426: begin
            cosine_reg0 <= 36'sb10011000111110001100010001011010100;
            sine_reg0   <= 36'sb11001101010001010000101001001000111;
        end
        2427: begin
            cosine_reg0 <= 36'sb10011000111001001001110010100000011;
            sine_reg0   <= 36'sb11001101010101000000110111100101000;
        end
        2428: begin
            cosine_reg0 <= 36'sb10011000110100000111001101101101000;
            sine_reg0   <= 36'sb11001101011000110000111110000110100;
        end
        2429: begin
            cosine_reg0 <= 36'sb10011000101111000100100011000000101;
            sine_reg0   <= 36'sb11001101011100100000111100101101010;
        end
        2430: begin
            cosine_reg0 <= 36'sb10011000101010000001110010011011011;
            sine_reg0   <= 36'sb11001101100000010000110011011001001;
        end
        2431: begin
            cosine_reg0 <= 36'sb10011000100100111110111011111101011;
            sine_reg0   <= 36'sb11001101100100000000100010001001111;
        end
        2432: begin
            cosine_reg0 <= 36'sb10011000011111111011111111100111000;
            sine_reg0   <= 36'sb11001101100111110000001000111111100;
        end
        2433: begin
            cosine_reg0 <= 36'sb10011000011010111000111101011000010;
            sine_reg0   <= 36'sb11001101101011011111100111111001110;
        end
        2434: begin
            cosine_reg0 <= 36'sb10011000010101110101110101010001100;
            sine_reg0   <= 36'sb11001101101111001110111110111000100;
        end
        2435: begin
            cosine_reg0 <= 36'sb10011000010000110010100111010010111;
            sine_reg0   <= 36'sb11001101110010111110001101111011100;
        end
        2436: begin
            cosine_reg0 <= 36'sb10011000001011101111010011011100100;
            sine_reg0   <= 36'sb11001101110110101101010101000010111;
        end
        2437: begin
            cosine_reg0 <= 36'sb10011000000110101011111001101110101;
            sine_reg0   <= 36'sb11001101111010011100010100001110010;
        end
        2438: begin
            cosine_reg0 <= 36'sb10011000000001101000011010001001100;
            sine_reg0   <= 36'sb11001101111110001011001011011101101;
        end
        2439: begin
            cosine_reg0 <= 36'sb10010111111100100100110100101101010;
            sine_reg0   <= 36'sb11001110000001111001111010110000101;
        end
        2440: begin
            cosine_reg0 <= 36'sb10010111110111100001001001011010000;
            sine_reg0   <= 36'sb11001110000101101000100010000111011;
        end
        2441: begin
            cosine_reg0 <= 36'sb10010111110010011101011000010000001;
            sine_reg0   <= 36'sb11001110001001010111000001100001101;
        end
        2442: begin
            cosine_reg0 <= 36'sb10010111101101011001100001001111110;
            sine_reg0   <= 36'sb11001110001101000101011000111111010;
        end
        2443: begin
            cosine_reg0 <= 36'sb10010111101000010101100100011001000;
            sine_reg0   <= 36'sb11001110010000110011101000100000000;
        end
        2444: begin
            cosine_reg0 <= 36'sb10010111100011010001100001101100001;
            sine_reg0   <= 36'sb11001110010100100001110000000011111;
        end
        2445: begin
            cosine_reg0 <= 36'sb10010111011110001101011001001001011;
            sine_reg0   <= 36'sb11001110011000001111101111101010110;
        end
        2446: begin
            cosine_reg0 <= 36'sb10010111011001001001001010110000110;
            sine_reg0   <= 36'sb11001110011011111101100111010100010;
        end
        2447: begin
            cosine_reg0 <= 36'sb10010111010100000100110110100010101;
            sine_reg0   <= 36'sb11001110011111101011010111000000100;
        end
        2448: begin
            cosine_reg0 <= 36'sb10010111001111000000011100011111010;
            sine_reg0   <= 36'sb11001110100011011000111110101111010;
        end
        2449: begin
            cosine_reg0 <= 36'sb10010111001001111011111100100110101;
            sine_reg0   <= 36'sb11001110100111000110011110100000010;
        end
        2450: begin
            cosine_reg0 <= 36'sb10010111000100110111010110111001000;
            sine_reg0   <= 36'sb11001110101010110011110110010011100;
        end
        2451: begin
            cosine_reg0 <= 36'sb10010110111111110010101011010110110;
            sine_reg0   <= 36'sb11001110101110100001000110001000111;
        end
        2452: begin
            cosine_reg0 <= 36'sb10010110111010101101111001111111110;
            sine_reg0   <= 36'sb11001110110010001110001110000000001;
        end
        2453: begin
            cosine_reg0 <= 36'sb10010110110101101001000010110100100;
            sine_reg0   <= 36'sb11001110110101111011001101111001001;
        end
        2454: begin
            cosine_reg0 <= 36'sb10010110110000100100000101110101000;
            sine_reg0   <= 36'sb11001110111001101000000101110011111;
        end
        2455: begin
            cosine_reg0 <= 36'sb10010110101011011111000011000001101;
            sine_reg0   <= 36'sb11001110111101010100110101110000000;
        end
        2456: begin
            cosine_reg0 <= 36'sb10010110100110011001111010011010011;
            sine_reg0   <= 36'sb11001111000001000001011101101101100;
        end
        2457: begin
            cosine_reg0 <= 36'sb10010110100001010100101011111111101;
            sine_reg0   <= 36'sb11001111000100101101111101101100010;
        end
        2458: begin
            cosine_reg0 <= 36'sb10010110011100001111010111110001011;
            sine_reg0   <= 36'sb11001111001000011010010101101100000;
        end
        2459: begin
            cosine_reg0 <= 36'sb10010110010111001001111101110000000;
            sine_reg0   <= 36'sb11001111001100000110100101101100110;
        end
        2460: begin
            cosine_reg0 <= 36'sb10010110010010000100011101111011100;
            sine_reg0   <= 36'sb11001111001111110010101101101110010;
        end
        2461: begin
            cosine_reg0 <= 36'sb10010110001100111110111000010100010;
            sine_reg0   <= 36'sb11001111010011011110101101110000011;
        end
        2462: begin
            cosine_reg0 <= 36'sb10010110000111111001001100111010100;
            sine_reg0   <= 36'sb11001111010111001010100101110011000;
        end
        2463: begin
            cosine_reg0 <= 36'sb10010110000010110011011011101110010;
            sine_reg0   <= 36'sb11001111011010110110010101110110000;
        end
        2464: begin
            cosine_reg0 <= 36'sb10010101111101101101100100101111110;
            sine_reg0   <= 36'sb11001111011110100001111101111001010;
        end
        2465: begin
            cosine_reg0 <= 36'sb10010101111000100111100111111111010;
            sine_reg0   <= 36'sb11001111100010001101011101111100100;
        end
        2466: begin
            cosine_reg0 <= 36'sb10010101110011100001100101011101000;
            sine_reg0   <= 36'sb11001111100101111000110101111111101;
        end
        2467: begin
            cosine_reg0 <= 36'sb10010101101110011011011101001001000;
            sine_reg0   <= 36'sb11001111101001100100000110000010101;
        end
        2468: begin
            cosine_reg0 <= 36'sb10010101101001010101001111000011101;
            sine_reg0   <= 36'sb11001111101101001111001110000101010;
        end
        2469: begin
            cosine_reg0 <= 36'sb10010101100100001110111011001101000;
            sine_reg0   <= 36'sb11001111110000111010001110000111011;
        end
        2470: begin
            cosine_reg0 <= 36'sb10010101011111001000100001100101011;
            sine_reg0   <= 36'sb11001111110100100101000110001000111;
        end
        2471: begin
            cosine_reg0 <= 36'sb10010101011010000010000010001100111;
            sine_reg0   <= 36'sb11001111111000001111110110001001101;
        end
        2472: begin
            cosine_reg0 <= 36'sb10010101010100111011011101000011110;
            sine_reg0   <= 36'sb11001111111011111010011110001001100;
        end
        2473: begin
            cosine_reg0 <= 36'sb10010101001111110100110010001010001;
            sine_reg0   <= 36'sb11001111111111100100111110001000001;
        end
        2474: begin
            cosine_reg0 <= 36'sb10010101001010101110000001100000011;
            sine_reg0   <= 36'sb11010000000011001111010110000101110;
        end
        2475: begin
            cosine_reg0 <= 36'sb10010101000101100111001011000110100;
            sine_reg0   <= 36'sb11010000000110111001100110000001111;
        end
        2476: begin
            cosine_reg0 <= 36'sb10010101000000100000001110111100101;
            sine_reg0   <= 36'sb11010000001010100011101101111100101;
        end
        2477: begin
            cosine_reg0 <= 36'sb10010100111011011001001101000011010;
            sine_reg0   <= 36'sb11010000001110001101101101110101101;
        end
        2478: begin
            cosine_reg0 <= 36'sb10010100110110010010000101011010011;
            sine_reg0   <= 36'sb11010000010001110111100101101101000;
        end
        2479: begin
            cosine_reg0 <= 36'sb10010100110001001010111000000010010;
            sine_reg0   <= 36'sb11010000010101100001010101100010011;
        end
        2480: begin
            cosine_reg0 <= 36'sb10010100101100000011100100111011000;
            sine_reg0   <= 36'sb11010000011001001010111101010101110;
        end
        2481: begin
            cosine_reg0 <= 36'sb10010100100110111100001100000100111;
            sine_reg0   <= 36'sb11010000011100110100011101000110111;
        end
        2482: begin
            cosine_reg0 <= 36'sb10010100100001110100101101100000001;
            sine_reg0   <= 36'sb11010000100000011101110100110101110;
        end
        2483: begin
            cosine_reg0 <= 36'sb10010100011100101101001001001100111;
            sine_reg0   <= 36'sb11010000100100000111000100100010001;
        end
        2484: begin
            cosine_reg0 <= 36'sb10010100010111100101011111001011011;
            sine_reg0   <= 36'sb11010000100111110000001100001011111;
        end
        2485: begin
            cosine_reg0 <= 36'sb10010100010010011101101111011011110;
            sine_reg0   <= 36'sb11010000101011011001001011110010111;
        end
        2486: begin
            cosine_reg0 <= 36'sb10010100001101010101111001111110010;
            sine_reg0   <= 36'sb11010000101111000010000011010111000;
        end
        2487: begin
            cosine_reg0 <= 36'sb10010100001000001101111110110011000;
            sine_reg0   <= 36'sb11010000110010101010110010111000000;
        end
        2488: begin
            cosine_reg0 <= 36'sb10010100000011000101111101111010011;
            sine_reg0   <= 36'sb11010000110110010011011010010101111;
        end
        2489: begin
            cosine_reg0 <= 36'sb10010011111101111101110111010100011;
            sine_reg0   <= 36'sb11010000111001111011111001110000100;
        end
        2490: begin
            cosine_reg0 <= 36'sb10010011111000110101101011000001010;
            sine_reg0   <= 36'sb11010000111101100100010001000111101;
        end
        2491: begin
            cosine_reg0 <= 36'sb10010011110011101101011001000001010;
            sine_reg0   <= 36'sb11010001000001001100100000011011001;
        end
        2492: begin
            cosine_reg0 <= 36'sb10010011101110100101000001010100101;
            sine_reg0   <= 36'sb11010001000100110100100111101011000;
        end
        2493: begin
            cosine_reg0 <= 36'sb10010011101001011100100011111011011;
            sine_reg0   <= 36'sb11010001001000011100100110110110111;
        end
        2494: begin
            cosine_reg0 <= 36'sb10010011100100010100000000110110000;
            sine_reg0   <= 36'sb11010001001100000100011101111110111;
        end
        2495: begin
            cosine_reg0 <= 36'sb10010011011111001011011000000100011;
            sine_reg0   <= 36'sb11010001001111101100001101000010101;
        end
        2496: begin
            cosine_reg0 <= 36'sb10010011011010000010101001100110111;
            sine_reg0   <= 36'sb11010001010011010011110100000010001;
        end
        2497: begin
            cosine_reg0 <= 36'sb10010011010100111001110101011101101;
            sine_reg0   <= 36'sb11010001010110111011010010111101001;
        end
        2498: begin
            cosine_reg0 <= 36'sb10010011001111110000111011101000111;
            sine_reg0   <= 36'sb11010001011010100010101001110011101;
        end
        2499: begin
            cosine_reg0 <= 36'sb10010011001010100111111100001000111;
            sine_reg0   <= 36'sb11010001011110001001111000100101011;
        end
        2500: begin
            cosine_reg0 <= 36'sb10010011000101011110110110111101101;
            sine_reg0   <= 36'sb11010001100001110000111111010010010;
        end
        2501: begin
            cosine_reg0 <= 36'sb10010011000000010101101100000111101;
            sine_reg0   <= 36'sb11010001100101010111111101111010010;
        end
        2502: begin
            cosine_reg0 <= 36'sb10010010111011001100011011100110110;
            sine_reg0   <= 36'sb11010001101000111110110100011101000;
        end
        2503: begin
            cosine_reg0 <= 36'sb10010010110110000011000101011011100;
            sine_reg0   <= 36'sb11010001101100100101100010111010100;
        end
        2504: begin
            cosine_reg0 <= 36'sb10010010110000111001101001100101110;
            sine_reg0   <= 36'sb11010001110000001100001001010010101;
        end
        2505: begin
            cosine_reg0 <= 36'sb10010010101011110000001000000110000;
            sine_reg0   <= 36'sb11010001110011110010100111100101010;
        end
        2506: begin
            cosine_reg0 <= 36'sb10010010100110100110100000111100010;
            sine_reg0   <= 36'sb11010001110111011000111101110010001;
        end
        2507: begin
            cosine_reg0 <= 36'sb10010010100001011100110100001000111;
            sine_reg0   <= 36'sb11010001111010111111001011111001010;
        end
        2508: begin
            cosine_reg0 <= 36'sb10010010011100010011000001101011111;
            sine_reg0   <= 36'sb11010001111110100101010001111010011;
        end
        2509: begin
            cosine_reg0 <= 36'sb10010010010111001001001001100101101;
            sine_reg0   <= 36'sb11010010000010001011001111110101011;
        end
        2510: begin
            cosine_reg0 <= 36'sb10010010010001111111001011110110001;
            sine_reg0   <= 36'sb11010010000101110001000101101010001;
        end
        2511: begin
            cosine_reg0 <= 36'sb10010010001100110101001000011101110;
            sine_reg0   <= 36'sb11010010001001010110110011011000100;
        end
        2512: begin
            cosine_reg0 <= 36'sb10010010000111101010111111011100110;
            sine_reg0   <= 36'sb11010010001100111100011001000000100;
        end
        2513: begin
            cosine_reg0 <= 36'sb10010010000010100000110000110011001;
            sine_reg0   <= 36'sb11010010010000100001110110100001101;
        end
        2514: begin
            cosine_reg0 <= 36'sb10010001111101010110011100100001001;
            sine_reg0   <= 36'sb11010010010100000111001011111100001;
        end
        2515: begin
            cosine_reg0 <= 36'sb10010001111000001100000010100111000;
            sine_reg0   <= 36'sb11010010010111101100011001001111101;
        end
        2516: begin
            cosine_reg0 <= 36'sb10010001110011000001100011000100111;
            sine_reg0   <= 36'sb11010010011011010001011110011100001;
        end
        2517: begin
            cosine_reg0 <= 36'sb10010001101101110110111101111011001;
            sine_reg0   <= 36'sb11010010011110110110011011100001011;
        end
        2518: begin
            cosine_reg0 <= 36'sb10010001101000101100010011001001110;
            sine_reg0   <= 36'sb11010010100010011011010000011111010;
        end
        2519: begin
            cosine_reg0 <= 36'sb10010001100011100001100010110001001;
            sine_reg0   <= 36'sb11010010100101111111111101010101101;
        end
        2520: begin
            cosine_reg0 <= 36'sb10010001011110010110101100110001010;
            sine_reg0   <= 36'sb11010010101001100100100010000100011;
        end
        2521: begin
            cosine_reg0 <= 36'sb10010001011001001011110001001010100;
            sine_reg0   <= 36'sb11010010101101001000111110101011100;
        end
        2522: begin
            cosine_reg0 <= 36'sb10010001010100000000101111111101000;
            sine_reg0   <= 36'sb11010010110000101101010011001010101;
        end
        2523: begin
            cosine_reg0 <= 36'sb10010001001110110101101001001001000;
            sine_reg0   <= 36'sb11010010110100010001011111100001110;
        end
        2524: begin
            cosine_reg0 <= 36'sb10010001001001101010011100101110101;
            sine_reg0   <= 36'sb11010010110111110101100011110000101;
        end
        2525: begin
            cosine_reg0 <= 36'sb10010001000100011111001010101110000;
            sine_reg0   <= 36'sb11010010111011011001011111110111010;
        end
        2526: begin
            cosine_reg0 <= 36'sb10010000111111010011110011000111101;
            sine_reg0   <= 36'sb11010010111110111101010011110101100;
        end
        2527: begin
            cosine_reg0 <= 36'sb10010000111010001000010101111011011;
            sine_reg0   <= 36'sb11010011000010100000111111101011001;
        end
        2528: begin
            cosine_reg0 <= 36'sb10010000110100111100110011001001100;
            sine_reg0   <= 36'sb11010011000110000100100011011000000;
        end
        2529: begin
            cosine_reg0 <= 36'sb10010000101111110001001010110010011;
            sine_reg0   <= 36'sb11010011001001100111111110111100000;
        end
        2530: begin
            cosine_reg0 <= 36'sb10010000101010100101011100110110001;
            sine_reg0   <= 36'sb11010011001101001011010010010111001;
        end
        2531: begin
            cosine_reg0 <= 36'sb10010000100101011001101001010100111;
            sine_reg0   <= 36'sb11010011010000101110011101101001000;
        end
        2532: begin
            cosine_reg0 <= 36'sb10010000100000001101110000001111000;
            sine_reg0   <= 36'sb11010011010100010001100000110001101;
        end
        2533: begin
            cosine_reg0 <= 36'sb10010000011011000001110001100100100;
            sine_reg0   <= 36'sb11010011010111110100011011110000111;
        end
        2534: begin
            cosine_reg0 <= 36'sb10010000010101110101101101010101101;
            sine_reg0   <= 36'sb11010011011011010111001110100110101;
        end
        2535: begin
            cosine_reg0 <= 36'sb10010000010000101001100011100010100;
            sine_reg0   <= 36'sb11010011011110111001111001010010101;
        end
        2536: begin
            cosine_reg0 <= 36'sb10010000001011011101010100001011101;
            sine_reg0   <= 36'sb11010011100010011100011011110100111;
        end
        2537: begin
            cosine_reg0 <= 36'sb10010000000110010000111111010000111;
            sine_reg0   <= 36'sb11010011100101111110110110001101001;
        end
        2538: begin
            cosine_reg0 <= 36'sb10010000000001000100100100110010101;
            sine_reg0   <= 36'sb11010011101001100001001000011011010;
        end
        2539: begin
            cosine_reg0 <= 36'sb10001111111011111000000100110001000;
            sine_reg0   <= 36'sb11010011101101000011010010011111010;
        end
        2540: begin
            cosine_reg0 <= 36'sb10001111110110101011011111001100010;
            sine_reg0   <= 36'sb11010011110000100101010100011000110;
        end
        2541: begin
            cosine_reg0 <= 36'sb10001111110001011110110100000100101;
            sine_reg0   <= 36'sb11010011110100000111001110000111111;
        end
        2542: begin
            cosine_reg0 <= 36'sb10001111101100010010000011011010001;
            sine_reg0   <= 36'sb11010011110111101000111111101100011;
        end
        2543: begin
            cosine_reg0 <= 36'sb10001111100111000101001101001101001;
            sine_reg0   <= 36'sb11010011111011001010101001000110001;
        end
        2544: begin
            cosine_reg0 <= 36'sb10001111100001111000010001011101111;
            sine_reg0   <= 36'sb11010011111110101100001010010100111;
        end
        2545: begin
            cosine_reg0 <= 36'sb10001111011100101011010000001100011;
            sine_reg0   <= 36'sb11010100000010001101100011011000101;
        end
        2546: begin
            cosine_reg0 <= 36'sb10001111010111011110001001011000111;
            sine_reg0   <= 36'sb11010100000101101110110100010001010;
        end
        2547: begin
            cosine_reg0 <= 36'sb10001111010010010000111101000011110;
            sine_reg0   <= 36'sb11010100001001001111111100111110100;
        end
        2548: begin
            cosine_reg0 <= 36'sb10001111001101000011101011001101000;
            sine_reg0   <= 36'sb11010100001100110000111101100000011;
        end
        2549: begin
            cosine_reg0 <= 36'sb10001111000111110110010011110101000;
            sine_reg0   <= 36'sb11010100010000010001110101110110101;
        end
        2550: begin
            cosine_reg0 <= 36'sb10001111000010101000110110111011111;
            sine_reg0   <= 36'sb11010100010011110010100110000001001;
        end
        2551: begin
            cosine_reg0 <= 36'sb10001110111101011011010100100001101;
            sine_reg0   <= 36'sb11010100010111010011001101111111111;
        end
        2552: begin
            cosine_reg0 <= 36'sb10001110111000001101101100100110111;
            sine_reg0   <= 36'sb11010100011010110011101101110010100;
        end
        2553: begin
            cosine_reg0 <= 36'sb10001110110010111111111111001011011;
            sine_reg0   <= 36'sb11010100011110010100000101011001001;
        end
        2554: begin
            cosine_reg0 <= 36'sb10001110101101110010001100001111101;
            sine_reg0   <= 36'sb11010100100001110100010100110011011;
        end
        2555: begin
            cosine_reg0 <= 36'sb10001110101000100100010011110011110;
            sine_reg0   <= 36'sb11010100100101010100011100000001011;
        end
        2556: begin
            cosine_reg0 <= 36'sb10001110100011010110010101111000000;
            sine_reg0   <= 36'sb11010100101000110100011011000010110;
        end
        2557: begin
            cosine_reg0 <= 36'sb10001110011110001000010010011100011;
            sine_reg0   <= 36'sb11010100101100010100010001110111100;
        end
        2558: begin
            cosine_reg0 <= 36'sb10001110011000111010001001100001011;
            sine_reg0   <= 36'sb11010100101111110100000000011111011;
        end
        2559: begin
            cosine_reg0 <= 36'sb10001110010011101011111011000110111;
            sine_reg0   <= 36'sb11010100110011010011100110111010011;
        end
        2560: begin
            cosine_reg0 <= 36'sb10001110001110011101100111001101011;
            sine_reg0   <= 36'sb11010100110110110011000101001000011;
        end
        2561: begin
            cosine_reg0 <= 36'sb10001110001001001111001101110100111;
            sine_reg0   <= 36'sb11010100111010010010011011001001001;
        end
        2562: begin
            cosine_reg0 <= 36'sb10001110000100000000101110111101110;
            sine_reg0   <= 36'sb11010100111101110001101000111100100;
        end
        2563: begin
            cosine_reg0 <= 36'sb10001101111110110010001010101000000;
            sine_reg0   <= 36'sb11010101000001010000101110100010011;
        end
        2564: begin
            cosine_reg0 <= 36'sb10001101111001100011100000110100000;
            sine_reg0   <= 36'sb11010101000100101111101011111010110;
        end
        2565: begin
            cosine_reg0 <= 36'sb10001101110100010100110001100001110;
            sine_reg0   <= 36'sb11010101001000001110100001000101011;
        end
        2566: begin
            cosine_reg0 <= 36'sb10001101101111000101111100110001101;
            sine_reg0   <= 36'sb11010101001011101101001110000010000;
        end
        2567: begin
            cosine_reg0 <= 36'sb10001101101001110111000010100011111;
            sine_reg0   <= 36'sb11010101001111001011110010110000110;
        end
        2568: begin
            cosine_reg0 <= 36'sb10001101100100101000000010111000100;
            sine_reg0   <= 36'sb11010101010010101010001111010001010;
        end
        2569: begin
            cosine_reg0 <= 36'sb10001101011111011000111101101111111;
            sine_reg0   <= 36'sb11010101010110001000100011100011101;
        end
        2570: begin
            cosine_reg0 <= 36'sb10001101011010001001110011001010001;
            sine_reg0   <= 36'sb11010101011001100110101111100111100;
        end
        2571: begin
            cosine_reg0 <= 36'sb10001101010100111010100011000111100;
            sine_reg0   <= 36'sb11010101011101000100110011011100110;
        end
        2572: begin
            cosine_reg0 <= 36'sb10001101001111101011001101101000001;
            sine_reg0   <= 36'sb11010101100000100010101111000011100;
        end
        2573: begin
            cosine_reg0 <= 36'sb10001101001010011011110010101100010;
            sine_reg0   <= 36'sb11010101100100000000100010011011010;
        end
        2574: begin
            cosine_reg0 <= 36'sb10001101000101001100010010010100000;
            sine_reg0   <= 36'sb11010101100111011110001101100100001;
        end
        2575: begin
            cosine_reg0 <= 36'sb10001100111111111100101100011111110;
            sine_reg0   <= 36'sb11010101101010111011110000011110000;
        end
        2576: begin
            cosine_reg0 <= 36'sb10001100111010101101000001001111100;
            sine_reg0   <= 36'sb11010101101110011001001011001000101;
        end
        2577: begin
            cosine_reg0 <= 36'sb10001100110101011101010000100011101;
            sine_reg0   <= 36'sb11010101110001110110011101100011111;
        end
        2578: begin
            cosine_reg0 <= 36'sb10001100110000001101011010011100010;
            sine_reg0   <= 36'sb11010101110101010011100111101111101;
        end
        2579: begin
            cosine_reg0 <= 36'sb10001100101010111101011110111001100;
            sine_reg0   <= 36'sb11010101111000110000101001101011111;
        end
        2580: begin
            cosine_reg0 <= 36'sb10001100100101101101011101111011110;
            sine_reg0   <= 36'sb11010101111100001101100011011000010;
        end
        2581: begin
            cosine_reg0 <= 36'sb10001100100000011101010111100011001;
            sine_reg0   <= 36'sb11010101111111101010010100110100110;
        end
        2582: begin
            cosine_reg0 <= 36'sb10001100011011001101001011101111110;
            sine_reg0   <= 36'sb11010110000011000110111110000001011;
        end
        2583: begin
            cosine_reg0 <= 36'sb10001100010101111100111010100001111;
            sine_reg0   <= 36'sb11010110000110100011011110111101110;
        end
        2584: begin
            cosine_reg0 <= 36'sb10001100010000101100100011111001110;
            sine_reg0   <= 36'sb11010110001001111111110111101001111;
        end
        2585: begin
            cosine_reg0 <= 36'sb10001100001011011100000111110111100;
            sine_reg0   <= 36'sb11010110001101011100001000000101101;
        end
        2586: begin
            cosine_reg0 <= 36'sb10001100000110001011100110011011100;
            sine_reg0   <= 36'sb11010110010000111000010000010000110;
        end
        2587: begin
            cosine_reg0 <= 36'sb10001100000000111010111111100101110;
            sine_reg0   <= 36'sb11010110010100010100010000001011010;
        end
        2588: begin
            cosine_reg0 <= 36'sb10001011111011101010010011010110100;
            sine_reg0   <= 36'sb11010110010111110000000111110100111;
        end
        2589: begin
            cosine_reg0 <= 36'sb10001011110110011001100001101110000;
            sine_reg0   <= 36'sb11010110011011001011110111001101101;
        end
        2590: begin
            cosine_reg0 <= 36'sb10001011110001001000101010101100011;
            sine_reg0   <= 36'sb11010110011110100111011110010101011;
        end
        2591: begin
            cosine_reg0 <= 36'sb10001011101011110111101110010010000;
            sine_reg0   <= 36'sb11010110100010000010111101001011111;
        end
        2592: begin
            cosine_reg0 <= 36'sb10001011100110100110101100011110111;
            sine_reg0   <= 36'sb11010110100101011110010011110001000;
        end
        2593: begin
            cosine_reg0 <= 36'sb10001011100001010101100101010011011;
            sine_reg0   <= 36'sb11010110101000111001100010000100101;
        end
        2594: begin
            cosine_reg0 <= 36'sb10001011011100000100011000101111100;
            sine_reg0   <= 36'sb11010110101100010100101000000110101;
        end
        2595: begin
            cosine_reg0 <= 36'sb10001011010110110011000110110011110;
            sine_reg0   <= 36'sb11010110101111101111100101110111000;
        end
        2596: begin
            cosine_reg0 <= 36'sb10001011010001100001101111100000000;
            sine_reg0   <= 36'sb11010110110011001010011011010101100;
        end
        2597: begin
            cosine_reg0 <= 36'sb10001011001100010000010010110100101;
            sine_reg0   <= 36'sb11010110110110100101001000100010000;
        end
        2598: begin
            cosine_reg0 <= 36'sb10001011000110111110110000110001111;
            sine_reg0   <= 36'sb11010110111001111111101101011100010;
        end
        2599: begin
            cosine_reg0 <= 36'sb10001011000001101101001001010111111;
            sine_reg0   <= 36'sb11010110111101011010001010000100011;
        end
        2600: begin
            cosine_reg0 <= 36'sb10001010111100011011011100100110110;
            sine_reg0   <= 36'sb11010111000000110100011110011010001;
        end
        2601: begin
            cosine_reg0 <= 36'sb10001010110111001001101010011110111;
            sine_reg0   <= 36'sb11010111000100001110101010011101010;
        end
        2602: begin
            cosine_reg0 <= 36'sb10001010110001110111110011000000011;
            sine_reg0   <= 36'sb11010111000111101000101110001101110;
        end
        2603: begin
            cosine_reg0 <= 36'sb10001010101100100101110110001011100;
            sine_reg0   <= 36'sb11010111001011000010101001101011100;
        end
        2604: begin
            cosine_reg0 <= 36'sb10001010100111010011110100000000010;
            sine_reg0   <= 36'sb11010111001110011100011100110110010;
        end
        2605: begin
            cosine_reg0 <= 36'sb10001010100010000001101100011111001;
            sine_reg0   <= 36'sb11010111010001110110000111101110001;
        end
        2606: begin
            cosine_reg0 <= 36'sb10001010011100101111011111101000001;
            sine_reg0   <= 36'sb11010111010101001111101010010010101;
        end
        2607: begin
            cosine_reg0 <= 36'sb10001010010111011101001101011011100;
            sine_reg0   <= 36'sb11010111011000101001000100100100000;
        end
        2608: begin
            cosine_reg0 <= 36'sb10001010010010001010110101111001100;
            sine_reg0   <= 36'sb11010111011100000010010110100001110;
        end
        2609: begin
            cosine_reg0 <= 36'sb10001010001100111000011001000010011;
            sine_reg0   <= 36'sb11010111011111011011100000001100000;
        end
        2610: begin
            cosine_reg0 <= 36'sb10001010000111100101110110110110001;
            sine_reg0   <= 36'sb11010111100010110100100001100010101;
        end
        2611: begin
            cosine_reg0 <= 36'sb10001010000010010011001111010101001;
            sine_reg0   <= 36'sb11010111100110001101011010100101011;
        end
        2612: begin
            cosine_reg0 <= 36'sb10001001111101000000100010011111100;
            sine_reg0   <= 36'sb11010111101001100110001011010100001;
        end
        2613: begin
            cosine_reg0 <= 36'sb10001001110111101101110000010101101;
            sine_reg0   <= 36'sb11010111101100111110110011101110110;
        end
        2614: begin
            cosine_reg0 <= 36'sb10001001110010011010111000110111011;
            sine_reg0   <= 36'sb11010111110000010111010011110101010;
        end
        2615: begin
            cosine_reg0 <= 36'sb10001001101101000111111100000101010;
            sine_reg0   <= 36'sb11010111110011101111101011100111010;
        end
        2616: begin
            cosine_reg0 <= 36'sb10001001100111110100111001111111011;
            sine_reg0   <= 36'sb11010111110111000111111011000100111;
        end
        2617: begin
            cosine_reg0 <= 36'sb10001001100010100001110010100101111;
            sine_reg0   <= 36'sb11010111111010100000000010001101111;
        end
        2618: begin
            cosine_reg0 <= 36'sb10001001011101001110100101111001000;
            sine_reg0   <= 36'sb11010111111101111000000001000010001;
        end
        2619: begin
            cosine_reg0 <= 36'sb10001001010111111011010011111001000;
            sine_reg0   <= 36'sb11011000000001001111110111100001100;
        end
        2620: begin
            cosine_reg0 <= 36'sb10001001010010100111111100100110001;
            sine_reg0   <= 36'sb11011000000100100111100101101011110;
        end
        2621: begin
            cosine_reg0 <= 36'sb10001001001101010100100000000000011;
            sine_reg0   <= 36'sb11011000000111111111001011100001000;
        end
        2622: begin
            cosine_reg0 <= 36'sb10001001001000000000111110001000001;
            sine_reg0   <= 36'sb11011000001011010110101001000001000;
        end
        2623: begin
            cosine_reg0 <= 36'sb10001001000010101101010110111101100;
            sine_reg0   <= 36'sb11011000001110101101111110001011100;
        end
        2624: begin
            cosine_reg0 <= 36'sb10001000111101011001101010100000110;
            sine_reg0   <= 36'sb11011000010010000101001011000000100;
        end
        2625: begin
            cosine_reg0 <= 36'sb10001000111000000101111000110010001;
            sine_reg0   <= 36'sb11011000010101011100001111011111111;
        end
        2626: begin
            cosine_reg0 <= 36'sb10001000110010110010000001110001110;
            sine_reg0   <= 36'sb11011000011000110011001011101001100;
        end
        2627: begin
            cosine_reg0 <= 36'sb10001000101101011110000101011111110;
            sine_reg0   <= 36'sb11011000011100001001111111011101001;
        end
        2628: begin
            cosine_reg0 <= 36'sb10001000101000001010000011111100100;
            sine_reg0   <= 36'sb11011000011111100000101010111010110;
        end
        2629: begin
            cosine_reg0 <= 36'sb10001000100010110101111101001000001;
            sine_reg0   <= 36'sb11011000100010110111001110000010010;
        end
        2630: begin
            cosine_reg0 <= 36'sb10001000011101100001110001000010111;
            sine_reg0   <= 36'sb11011000100110001101101000110011011;
        end
        2631: begin
            cosine_reg0 <= 36'sb10001000011000001101011111101100111;
            sine_reg0   <= 36'sb11011000101001100011111011001110001;
        end
        2632: begin
            cosine_reg0 <= 36'sb10001000010010111001001001000110100;
            sine_reg0   <= 36'sb11011000101100111010000101010010010;
        end
        2633: begin
            cosine_reg0 <= 36'sb10001000001101100100101101001111101;
            sine_reg0   <= 36'sb11011000110000010000000110111111110;
        end
        2634: begin
            cosine_reg0 <= 36'sb10001000001000010000001100001000111;
            sine_reg0   <= 36'sb11011000110011100110000000010110011;
        end
        2635: begin
            cosine_reg0 <= 36'sb10001000000010111011100101110010001;
            sine_reg0   <= 36'sb11011000110110111011110001010110001;
        end
        2636: begin
            cosine_reg0 <= 36'sb10000111111101100110111010001011101;
            sine_reg0   <= 36'sb11011000111010010001011001111110110;
        end
        2637: begin
            cosine_reg0 <= 36'sb10000111111000010010001001010101110;
            sine_reg0   <= 36'sb11011000111101100110111010010000001;
        end
        2638: begin
            cosine_reg0 <= 36'sb10000111110010111101010011010000101;
            sine_reg0   <= 36'sb11011001000000111100010010001010010;
        end
        2639: begin
            cosine_reg0 <= 36'sb10000111101101101000010111111100011;
            sine_reg0   <= 36'sb11011001000100010001100001101100111;
        end
        2640: begin
            cosine_reg0 <= 36'sb10000111101000010011010111011001010;
            sine_reg0   <= 36'sb11011001000111100110101000110111111;
        end
        2641: begin
            cosine_reg0 <= 36'sb10000111100010111110010001100111100;
            sine_reg0   <= 36'sb11011001001010111011100111101011010;
        end
        2642: begin
            cosine_reg0 <= 36'sb10000111011101101001000110100111011;
            sine_reg0   <= 36'sb11011001001110010000011110000110101;
        end
        2643: begin
            cosine_reg0 <= 36'sb10000111011000010011110110011000111;
            sine_reg0   <= 36'sb11011001010001100101001100001010001;
        end
        2644: begin
            cosine_reg0 <= 36'sb10000111010010111110100000111100011;
            sine_reg0   <= 36'sb11011001010100111001110001110101100;
        end
        2645: begin
            cosine_reg0 <= 36'sb10000111001101101001000110010010001;
            sine_reg0   <= 36'sb11011001011000001110001111001000110;
        end
        2646: begin
            cosine_reg0 <= 36'sb10000111001000010011100110011010010;
            sine_reg0   <= 36'sb11011001011011100010100100000011100;
        end
        2647: begin
            cosine_reg0 <= 36'sb10000111000010111110000001010100111;
            sine_reg0   <= 36'sb11011001011110110110110000100101110;
        end
        2648: begin
            cosine_reg0 <= 36'sb10000110111101101000010111000010010;
            sine_reg0   <= 36'sb11011001100010001010110100101111100;
        end
        2649: begin
            cosine_reg0 <= 36'sb10000110111000010010100111100010110;
            sine_reg0   <= 36'sb11011001100101011110110000100000100;
        end
        2650: begin
            cosine_reg0 <= 36'sb10000110110010111100110010110110011;
            sine_reg0   <= 36'sb11011001101000110010100011111000100;
        end
        2651: begin
            cosine_reg0 <= 36'sb10000110101101100110111000111101011;
            sine_reg0   <= 36'sb11011001101100000110001110110111101;
        end
        2652: begin
            cosine_reg0 <= 36'sb10000110101000010000111001111000000;
            sine_reg0   <= 36'sb11011001101111011001110001011101100;
        end
        2653: begin
            cosine_reg0 <= 36'sb10000110100010111010110101100110100;
            sine_reg0   <= 36'sb11011001110010101101001011101010010;
        end
        2654: begin
            cosine_reg0 <= 36'sb10000110011101100100101100001001000;
            sine_reg0   <= 36'sb11011001110110000000011101011101101;
        end
        2655: begin
            cosine_reg0 <= 36'sb10000110011000001110011101011111110;
            sine_reg0   <= 36'sb11011001111001010011100110110111011;
        end
        2656: begin
            cosine_reg0 <= 36'sb10000110010010111000001001101010111;
            sine_reg0   <= 36'sb11011001111100100110100111110111100;
        end
        2657: begin
            cosine_reg0 <= 36'sb10000110001101100001110000101010101;
            sine_reg0   <= 36'sb11011001111111111001100000011110000;
        end
        2658: begin
            cosine_reg0 <= 36'sb10000110001000001011010010011111010;
            sine_reg0   <= 36'sb11011010000011001100010000101010100;
        end
        2659: begin
            cosine_reg0 <= 36'sb10000110000010110100101111001001000;
            sine_reg0   <= 36'sb11011010000110011110111000011101000;
        end
        2660: begin
            cosine_reg0 <= 36'sb10000101111101011110000110100111111;
            sine_reg0   <= 36'sb11011010001001110001010111110101011;
        end
        2661: begin
            cosine_reg0 <= 36'sb10000101111000000111011000111100011;
            sine_reg0   <= 36'sb11011010001101000011101110110011100;
        end
        2662: begin
            cosine_reg0 <= 36'sb10000101110010110000100110000110011;
            sine_reg0   <= 36'sb11011010010000010101111101010111001;
        end
        2663: begin
            cosine_reg0 <= 36'sb10000101101101011001101110000110011;
            sine_reg0   <= 36'sb11011010010011101000000011100000011;
        end
        2664: begin
            cosine_reg0 <= 36'sb10000101101000000010110000111100011;
            sine_reg0   <= 36'sb11011010010110111010000001001110111;
        end
        2665: begin
            cosine_reg0 <= 36'sb10000101100010101011101110101000110;
            sine_reg0   <= 36'sb11011010011010001011110110100010101;
        end
        2666: begin
            cosine_reg0 <= 36'sb10000101011101010100100111001011101;
            sine_reg0   <= 36'sb11011010011101011101100011011011011;
        end
        2667: begin
            cosine_reg0 <= 36'sb10000101010111111101011010100101001;
            sine_reg0   <= 36'sb11011010100000101111000111111001010;
        end
        2668: begin
            cosine_reg0 <= 36'sb10000101010010100110001000110101101;
            sine_reg0   <= 36'sb11011010100100000000100011111011111;
        end
        2669: begin
            cosine_reg0 <= 36'sb10000101001101001110110001111101001;
            sine_reg0   <= 36'sb11011010100111010001110111100011010;
        end
        2670: begin
            cosine_reg0 <= 36'sb10000101000111110111010101111100001;
            sine_reg0   <= 36'sb11011010101010100011000010101111010;
        end
        2671: begin
            cosine_reg0 <= 36'sb10000101000010011111110100110010100;
            sine_reg0   <= 36'sb11011010101101110100000101011111101;
        end
        2672: begin
            cosine_reg0 <= 36'sb10000100111101001000001110100000101;
            sine_reg0   <= 36'sb11011010110001000100111111110100100;
        end
        2673: begin
            cosine_reg0 <= 36'sb10000100110111110000100011000110110;
            sine_reg0   <= 36'sb11011010110100010101110001101101100;
        end
        2674: begin
            cosine_reg0 <= 36'sb10000100110010011000110010100101001;
            sine_reg0   <= 36'sb11011010110111100110011011001010100;
        end
        2675: begin
            cosine_reg0 <= 36'sb10000100101101000000111100111011110;
            sine_reg0   <= 36'sb11011010111010110110111100001011101;
        end
        2676: begin
            cosine_reg0 <= 36'sb10000100100111101001000010001010111;
            sine_reg0   <= 36'sb11011010111110000111010100110000100;
        end
        2677: begin
            cosine_reg0 <= 36'sb10000100100010010001000010010010111;
            sine_reg0   <= 36'sb11011011000001010111100100111001000;
        end
        2678: begin
            cosine_reg0 <= 36'sb10000100011100111000111101010011111;
            sine_reg0   <= 36'sb11011011000100100111101100100101010;
        end
        2679: begin
            cosine_reg0 <= 36'sb10000100010111100000110011001110000;
            sine_reg0   <= 36'sb11011011000111110111101011110100111;
        end
        2680: begin
            cosine_reg0 <= 36'sb10000100010010001000100100000001100;
            sine_reg0   <= 36'sb11011011001011000111100010100111111;
        end
        2681: begin
            cosine_reg0 <= 36'sb10000100001100110000001111101110101;
            sine_reg0   <= 36'sb11011011001110010111010000111110000;
        end
        2682: begin
            cosine_reg0 <= 36'sb10000100000111010111110110010101101;
            sine_reg0   <= 36'sb11011011010001100110110110110111010;
        end
        2683: begin
            cosine_reg0 <= 36'sb10000100000001111111010111110110101;
            sine_reg0   <= 36'sb11011011010100110110010100010011100;
        end
        2684: begin
            cosine_reg0 <= 36'sb10000011111100100110110100010001110;
            sine_reg0   <= 36'sb11011011011000000101101001010010101;
        end
        2685: begin
            cosine_reg0 <= 36'sb10000011110111001110001011100111100;
            sine_reg0   <= 36'sb11011011011011010100110101110100011;
        end
        2686: begin
            cosine_reg0 <= 36'sb10000011110001110101011101110111110;
            sine_reg0   <= 36'sb11011011011110100011111001111000110;
        end
        2687: begin
            cosine_reg0 <= 36'sb10000011101100011100101011000010111;
            sine_reg0   <= 36'sb11011011100001110010110101011111100;
        end
        2688: begin
            cosine_reg0 <= 36'sb10000011100111000011110011001001000;
            sine_reg0   <= 36'sb11011011100101000001101000101000101;
        end
        2689: begin
            cosine_reg0 <= 36'sb10000011100001101010110110001010100;
            sine_reg0   <= 36'sb11011011101000010000010011010100000;
        end
        2690: begin
            cosine_reg0 <= 36'sb10000011011100010001110100000111011;
            sine_reg0   <= 36'sb11011011101011011110110101100001100;
        end
        2691: begin
            cosine_reg0 <= 36'sb10000011010110111000101101000000000;
            sine_reg0   <= 36'sb11011011101110101101001111010000111;
        end
        2692: begin
            cosine_reg0 <= 36'sb10000011010001011111100000110100100;
            sine_reg0   <= 36'sb11011011110001111011100000100010010;
        end
        2693: begin
            cosine_reg0 <= 36'sb10000011001100000110001111100101001;
            sine_reg0   <= 36'sb11011011110101001001101001010101001;
        end
        2694: begin
            cosine_reg0 <= 36'sb10000011000110101100111001010010000;
            sine_reg0   <= 36'sb11011011111000010111101001101001110;
        end
        2695: begin
            cosine_reg0 <= 36'sb10000011000001010011011101111011011;
            sine_reg0   <= 36'sb11011011111011100101100001011111110;
        end
        2696: begin
            cosine_reg0 <= 36'sb10000010111011111001111101100001100;
            sine_reg0   <= 36'sb11011011111110110011010000110111001;
        end
        2697: begin
            cosine_reg0 <= 36'sb10000010110110100000011000000100100;
            sine_reg0   <= 36'sb11011100000010000000110111101111110;
        end
        2698: begin
            cosine_reg0 <= 36'sb10000010110001000110101101100100110;
            sine_reg0   <= 36'sb11011100000101001110010110001001011;
        end
        2699: begin
            cosine_reg0 <= 36'sb10000010101011101100111110000010010;
            sine_reg0   <= 36'sb11011100001000011011101100000100000;
        end
        2700: begin
            cosine_reg0 <= 36'sb10000010100110010011001001011101011;
            sine_reg0   <= 36'sb11011100001011101000111001011111100;
        end
        2701: begin
            cosine_reg0 <= 36'sb10000010100000111001001111110110010;
            sine_reg0   <= 36'sb11011100001110110101111110011011110;
        end
        2702: begin
            cosine_reg0 <= 36'sb10000010011011011111010001001101000;
            sine_reg0   <= 36'sb11011100010010000010111010111000101;
        end
        2703: begin
            cosine_reg0 <= 36'sb10000010010110000101001101100010000;
            sine_reg0   <= 36'sb11011100010101001111101110110101111;
        end
        2704: begin
            cosine_reg0 <= 36'sb10000010010000101011000100110101011;
            sine_reg0   <= 36'sb11011100011000011100011010010011100;
        end
        2705: begin
            cosine_reg0 <= 36'sb10000010001011010000110111000111011;
            sine_reg0   <= 36'sb11011100011011101000111101010001011;
        end
        2706: begin
            cosine_reg0 <= 36'sb10000010000101110110100100011000001;
            sine_reg0   <= 36'sb11011100011110110101010111101111011;
        end
        2707: begin
            cosine_reg0 <= 36'sb10000010000000011100001100100111111;
            sine_reg0   <= 36'sb11011100100010000001101001101101011;
        end
        2708: begin
            cosine_reg0 <= 36'sb10000001111011000001101111110110111;
            sine_reg0   <= 36'sb11011100100101001101110011001011010;
        end
        2709: begin
            cosine_reg0 <= 36'sb10000001110101100111001110000101011;
            sine_reg0   <= 36'sb11011100101000011001110100001000110;
        end
        2710: begin
            cosine_reg0 <= 36'sb10000001110000001100100111010011100;
            sine_reg0   <= 36'sb11011100101011100101101100100110000;
        end
        2711: begin
            cosine_reg0 <= 36'sb10000001101010110001111011100001011;
            sine_reg0   <= 36'sb11011100101110110001011100100010101;
        end
        2712: begin
            cosine_reg0 <= 36'sb10000001100101010111001010101111011;
            sine_reg0   <= 36'sb11011100110001111101000011111110101;
        end
        2713: begin
            cosine_reg0 <= 36'sb10000001011111111100010100111101101;
            sine_reg0   <= 36'sb11011100110101001000100010111010000;
        end
        2714: begin
            cosine_reg0 <= 36'sb10000001011010100001011010001100011;
            sine_reg0   <= 36'sb11011100111000010011111001010100011;
        end
        2715: begin
            cosine_reg0 <= 36'sb10000001010101000110011010011011110;
            sine_reg0   <= 36'sb11011100111011011111000111001101110;
        end
        2716: begin
            cosine_reg0 <= 36'sb10000001001111101011010101101100000;
            sine_reg0   <= 36'sb11011100111110101010001100100110001;
        end
        2717: begin
            cosine_reg0 <= 36'sb10000001001010010000001011111101011;
            sine_reg0   <= 36'sb11011101000001110101001001011101001;
        end
        2718: begin
            cosine_reg0 <= 36'sb10000001000100110100111101010000001;
            sine_reg0   <= 36'sb11011101000100111111111101110010110;
        end
        2719: begin
            cosine_reg0 <= 36'sb10000000111111011001101001100100011;
            sine_reg0   <= 36'sb11011101001000001010101001100111000;
        end
        2720: begin
            cosine_reg0 <= 36'sb10000000111001111110010000111010011;
            sine_reg0   <= 36'sb11011101001011010101001100111001101;
        end
        2721: begin
            cosine_reg0 <= 36'sb10000000110100100010110011010010010;
            sine_reg0   <= 36'sb11011101001110011111100111101010011;
        end
        2722: begin
            cosine_reg0 <= 36'sb10000000101111000111010000101100010;
            sine_reg0   <= 36'sb11011101010001101001111001111001011;
        end
        2723: begin
            cosine_reg0 <= 36'sb10000000101001101011101001001000101;
            sine_reg0   <= 36'sb11011101010100110100000011100110011;
        end
        2724: begin
            cosine_reg0 <= 36'sb10000000100100001111111100100111101;
            sine_reg0   <= 36'sb11011101010111111110000100110001011;
        end
        2725: begin
            cosine_reg0 <= 36'sb10000000011110110100001011001001011;
            sine_reg0   <= 36'sb11011101011011000111111101011010000;
        end
        2726: begin
            cosine_reg0 <= 36'sb10000000011001011000010100101110001;
            sine_reg0   <= 36'sb11011101011110010001101101100000011;
        end
        2727: begin
            cosine_reg0 <= 36'sb10000000010011111100011001010110000;
            sine_reg0   <= 36'sb11011101100001011011010101000100010;
        end
        2728: begin
            cosine_reg0 <= 36'sb10000000001110100000011001000001010;
            sine_reg0   <= 36'sb11011101100100100100110100000101101;
        end
        2729: begin
            cosine_reg0 <= 36'sb10000000001001000100010011110000010;
            sine_reg0   <= 36'sb11011101100111101110001010100100010;
        end
        2730: begin
            cosine_reg0 <= 36'sb10000000000011101000001001100011000;
            sine_reg0   <= 36'sb11011101101010110111011000100000000;
        end
        2731: begin
            cosine_reg0 <= 36'sb1111111111110001011111010011001110;
            sine_reg0   <= 36'sb11011101101110000000011101111000111;
        end
        2732: begin
            cosine_reg0 <= 36'sb1111111111000101111100110010100110;
            sine_reg0   <= 36'sb11011101110001001001011010101110101;
        end
        2733: begin
            cosine_reg0 <= 36'sb1111111110011010011001101010100010;
            sine_reg0   <= 36'sb11011101110100010010001111000001001;
        end
        2734: begin
            cosine_reg0 <= 36'sb1111111101101110110101111011000011;
            sine_reg0   <= 36'sb11011101110111011010111010110000011;
        end
        2735: begin
            cosine_reg0 <= 36'sb1111111101000011010001100100001100;
            sine_reg0   <= 36'sb11011101111010100011011101111100010;
        end
        2736: begin
            cosine_reg0 <= 36'sb1111111100010111101100100101111100;
            sine_reg0   <= 36'sb11011101111101101011111000100100100;
        end
        2737: begin
            cosine_reg0 <= 36'sb1111111011101100000111000000011000;
            sine_reg0   <= 36'sb11011110000000110100001010101001001;
        end
        2738: begin
            cosine_reg0 <= 36'sb1111111011000000100000110011011111;
            sine_reg0   <= 36'sb11011110000011111100010100001001111;
        end
        2739: begin
            cosine_reg0 <= 36'sb1111111010010100111001111111010100;
            sine_reg0   <= 36'sb11011110000111000100010101000110110;
        end
        2740: begin
            cosine_reg0 <= 36'sb1111111001101001010010100011111000;
            sine_reg0   <= 36'sb11011110001010001100001101011111101;
        end
        2741: begin
            cosine_reg0 <= 36'sb1111111000111101101010100001001101;
            sine_reg0   <= 36'sb11011110001101010011111101010100011;
        end
        2742: begin
            cosine_reg0 <= 36'sb1111111000010010000001110111010101;
            sine_reg0   <= 36'sb11011110010000011011100100100100110;
        end
        2743: begin
            cosine_reg0 <= 36'sb1111110111100110011000100110010010;
            sine_reg0   <= 36'sb11011110010011100011000011010000110;
        end
        2744: begin
            cosine_reg0 <= 36'sb1111110110111010101110101110000100;
            sine_reg0   <= 36'sb11011110010110101010011001011000010;
        end
        2745: begin
            cosine_reg0 <= 36'sb1111110110001111000100001110101110;
            sine_reg0   <= 36'sb11011110011001110001100110111011001;
        end
        2746: begin
            cosine_reg0 <= 36'sb1111110101100011011001001000010010;
            sine_reg0   <= 36'sb11011110011100111000101011111001010;
        end
        2747: begin
            cosine_reg0 <= 36'sb1111110100110111101101011010110001;
            sine_reg0   <= 36'sb11011110011111111111101000010010100;
        end
        2748: begin
            cosine_reg0 <= 36'sb1111110100001100000001000110001101;
            sine_reg0   <= 36'sb11011110100011000110011100000110110;
        end
        2749: begin
            cosine_reg0 <= 36'sb1111110011100000010100001010100111;
            sine_reg0   <= 36'sb11011110100110001101000111010101111;
        end
        2750: begin
            cosine_reg0 <= 36'sb1111110010110100100110101000000010;
            sine_reg0   <= 36'sb11011110101001010011101001111111110;
        end
        2751: begin
            cosine_reg0 <= 36'sb1111110010001000111000011110011111;
            sine_reg0   <= 36'sb11011110101100011010000100000100011;
        end
        2752: begin
            cosine_reg0 <= 36'sb1111110001011101001001101101111111;
            sine_reg0   <= 36'sb11011110101111100000010101100011011;
        end
        2753: begin
            cosine_reg0 <= 36'sb1111110000110001011010010110100100;
            sine_reg0   <= 36'sb11011110110010100110011110011100111;
        end
        2754: begin
            cosine_reg0 <= 36'sb1111110000000101101010011000010000;
            sine_reg0   <= 36'sb11011110110101101100011110110000101;
        end
        2755: begin
            cosine_reg0 <= 36'sb1111101111011001111001110011000101;
            sine_reg0   <= 36'sb11011110111000110010010110011110100;
        end
        2756: begin
            cosine_reg0 <= 36'sb1111101110101110001000100111000100;
            sine_reg0   <= 36'sb11011110111011111000000101100110100;
        end
        2757: begin
            cosine_reg0 <= 36'sb1111101110000010010110110100010000;
            sine_reg0   <= 36'sb11011110111110111101101100001000011;
        end
        2758: begin
            cosine_reg0 <= 36'sb1111101101010110100100011010101001;
            sine_reg0   <= 36'sb11011111000010000011001010000100001;
        end
        2759: begin
            cosine_reg0 <= 36'sb1111101100101010110001011010010001;
            sine_reg0   <= 36'sb11011111000101001000011111011001100;
        end
        2760: begin
            cosine_reg0 <= 36'sb1111101011111110111101110011001010;
            sine_reg0   <= 36'sb11011111001000001101101100001000011;
        end
        2761: begin
            cosine_reg0 <= 36'sb1111101011010011001001100101010111;
            sine_reg0   <= 36'sb11011111001011010010110000010000111;
        end
        2762: begin
            cosine_reg0 <= 36'sb1111101010100111010100110000110111;
            sine_reg0   <= 36'sb11011111001110010111101011110010101;
        end
        2763: begin
            cosine_reg0 <= 36'sb1111101001111011011111010101101110;
            sine_reg0   <= 36'sb11011111010001011100011110101101101;
        end
        2764: begin
            cosine_reg0 <= 36'sb1111101001001111101001010011111101;
            sine_reg0   <= 36'sb11011111010100100001001001000001101;
        end
        2765: begin
            cosine_reg0 <= 36'sb1111101000100011110010101011100101;
            sine_reg0   <= 36'sb11011111010111100101101010101110101;
        end
        2766: begin
            cosine_reg0 <= 36'sb1111100111110111111011011100101000;
            sine_reg0   <= 36'sb11011111011010101010000011110100101;
        end
        2767: begin
            cosine_reg0 <= 36'sb1111100111001100000011100111001001;
            sine_reg0   <= 36'sb11011111011101101110010100010011010;
        end
        2768: begin
            cosine_reg0 <= 36'sb1111100110100000001011001011000111;
            sine_reg0   <= 36'sb11011111100000110010011100001010100;
        end
        2769: begin
            cosine_reg0 <= 36'sb1111100101110100010010001000100111;
            sine_reg0   <= 36'sb11011111100011110110011011011010010;
        end
        2770: begin
            cosine_reg0 <= 36'sb1111100101001000011000011111101000;
            sine_reg0   <= 36'sb11011111100110111010010010000010011;
        end
        2771: begin
            cosine_reg0 <= 36'sb1111100100011100011110010000001101;
            sine_reg0   <= 36'sb11011111101001111110000000000010111;
        end
        2772: begin
            cosine_reg0 <= 36'sb1111100011110000100011011010010111;
            sine_reg0   <= 36'sb11011111101101000001100101011011100;
        end
        2773: begin
            cosine_reg0 <= 36'sb1111100011000100100111111110001000;
            sine_reg0   <= 36'sb11011111110000000101000010001100001;
        end
        2774: begin
            cosine_reg0 <= 36'sb1111100010011000101011111011100010;
            sine_reg0   <= 36'sb11011111110011001000010110010100101;
        end
        2775: begin
            cosine_reg0 <= 36'sb1111100001101100101111010010100111;
            sine_reg0   <= 36'sb11011111110110001011100001110100111;
        end
        2776: begin
            cosine_reg0 <= 36'sb1111100001000000110010000011011000;
            sine_reg0   <= 36'sb11011111111001001110100100101101000;
        end
        2777: begin
            cosine_reg0 <= 36'sb1111100000010100110100001101110110;
            sine_reg0   <= 36'sb11011111111100010001011110111100100;
        end
        2778: begin
            cosine_reg0 <= 36'sb1111011111101000110101110010000100;
            sine_reg0   <= 36'sb11011111111111010100010000100011100;
        end
        2779: begin
            cosine_reg0 <= 36'sb1111011110111100110110110000000011;
            sine_reg0   <= 36'sb11100000000010010110111001100001111;
        end
        2780: begin
            cosine_reg0 <= 36'sb1111011110010000110111000111110101;
            sine_reg0   <= 36'sb11100000000101011001011001110111100;
        end
        2781: begin
            cosine_reg0 <= 36'sb1111011101100100110110111001011100;
            sine_reg0   <= 36'sb11100000001000011011110001100100001;
        end
        2782: begin
            cosine_reg0 <= 36'sb1111011100111000110110000100111001;
            sine_reg0   <= 36'sb11100000001011011110000000100111110;
        end
        2783: begin
            cosine_reg0 <= 36'sb1111011100001100110100101010001111;
            sine_reg0   <= 36'sb11100000001110100000000111000010010;
        end
        2784: begin
            cosine_reg0 <= 36'sb1111011011100000110010101001011101;
            sine_reg0   <= 36'sb11100000010001100010000100110011100;
        end
        2785: begin
            cosine_reg0 <= 36'sb1111011010110100110000000010101000;
            sine_reg0   <= 36'sb11100000010100100011111001111011011;
        end
        2786: begin
            cosine_reg0 <= 36'sb1111011010001000101100110101101111;
            sine_reg0   <= 36'sb11100000010111100101100110011001110;
        end
        2787: begin
            cosine_reg0 <= 36'sb1111011001011100101001000010110101;
            sine_reg0   <= 36'sb11100000011010100111001010001110100;
        end
        2788: begin
            cosine_reg0 <= 36'sb1111011000110000100100101001111100;
            sine_reg0   <= 36'sb11100000011101101000100101011001100;
        end
        2789: begin
            cosine_reg0 <= 36'sb1111011000000100011111101011000101;
            sine_reg0   <= 36'sb11100000100000101001110111111010110;
        end
        2790: begin
            cosine_reg0 <= 36'sb1111010111011000011010000110010010;
            sine_reg0   <= 36'sb11100000100011101011000001110010000;
        end
        2791: begin
            cosine_reg0 <= 36'sb1111010110101100010011111011100100;
            sine_reg0   <= 36'sb11100000100110101100000010111111001;
        end
        2792: begin
            cosine_reg0 <= 36'sb1111010110000000001101001010111110;
            sine_reg0   <= 36'sb11100000101001101100111011100010001;
        end
        2793: begin
            cosine_reg0 <= 36'sb1111010101010100000101110100100001;
            sine_reg0   <= 36'sb11100000101100101101101011011010110;
        end
        2794: begin
            cosine_reg0 <= 36'sb1111010100100111111101111000001110;
            sine_reg0   <= 36'sb11100000101111101110010010101001000;
        end
        2795: begin
            cosine_reg0 <= 36'sb1111010011111011110101010110001000;
            sine_reg0   <= 36'sb11100000110010101110110001001100110;
        end
        2796: begin
            cosine_reg0 <= 36'sb1111010011001111101100001110010000;
            sine_reg0   <= 36'sb11100000110101101111000111000101110;
        end
        2797: begin
            cosine_reg0 <= 36'sb1111010010100011100010100000100111;
            sine_reg0   <= 36'sb11100000111000101111010100010100001;
        end
        2798: begin
            cosine_reg0 <= 36'sb1111010001110111011000001101010001;
            sine_reg0   <= 36'sb11100000111011101111011000110111100;
        end
        2799: begin
            cosine_reg0 <= 36'sb1111010001001011001101010100001101;
            sine_reg0   <= 36'sb11100000111110101111010100101111111;
        end
        2800: begin
            cosine_reg0 <= 36'sb1111010000011111000001110101011111;
            sine_reg0   <= 36'sb11100001000001101111000111111101001;
        end
        2801: begin
            cosine_reg0 <= 36'sb1111001111110010110101110001000111;
            sine_reg0   <= 36'sb11100001000100101110110010011111010;
        end
        2802: begin
            cosine_reg0 <= 36'sb1111001111000110101001000111000111;
            sine_reg0   <= 36'sb11100001000111101110010100010110000;
        end
        2803: begin
            cosine_reg0 <= 36'sb1111001110011010011011110111100001;
            sine_reg0   <= 36'sb11100001001010101101101101100001010;
        end
        2804: begin
            cosine_reg0 <= 36'sb1111001101101110001110000010010111;
            sine_reg0   <= 36'sb11100001001101101100111110000000111;
        end
        2805: begin
            cosine_reg0 <= 36'sb1111001101000001111111100111101011;
            sine_reg0   <= 36'sb11100001010000101100000101110100111;
        end
        2806: begin
            cosine_reg0 <= 36'sb1111001100010101110000100111011110;
            sine_reg0   <= 36'sb11100001010011101011000100111101000;
        end
        2807: begin
            cosine_reg0 <= 36'sb1111001011101001100001000001110001;
            sine_reg0   <= 36'sb11100001010110101001111011011001010;
        end
        2808: begin
            cosine_reg0 <= 36'sb1111001010111101010000110110100111;
            sine_reg0   <= 36'sb11100001011001101000101001001001100;
        end
        2809: begin
            cosine_reg0 <= 36'sb1111001010010001000000000110000001;
            sine_reg0   <= 36'sb11100001011100100111001110001101100;
        end
        2810: begin
            cosine_reg0 <= 36'sb1111001001100100101110110000000010;
            sine_reg0   <= 36'sb11100001011111100101101010100101010;
        end
        2811: begin
            cosine_reg0 <= 36'sb1111001000111000011100110100101010;
            sine_reg0   <= 36'sb11100001100010100011111110010000101;
        end
        2812: begin
            cosine_reg0 <= 36'sb1111001000001100001010010011111011;
            sine_reg0   <= 36'sb11100001100101100010001001001111101;
        end
        2813: begin
            cosine_reg0 <= 36'sb1111000111011111110111001101110111;
            sine_reg0   <= 36'sb11100001101000100000001011100001111;
        end
        2814: begin
            cosine_reg0 <= 36'sb1111000110110011100011100010100001;
            sine_reg0   <= 36'sb11100001101011011110000101000111011;
        end
        2815: begin
            cosine_reg0 <= 36'sb1111000110000111001111010001111000;
            sine_reg0   <= 36'sb11100001101110011011110110000000001;
        end
        2816: begin
            cosine_reg0 <= 36'sb1111000101011010111010011100000000;
            sine_reg0   <= 36'sb11100001110001011001011110001011111;
        end
        2817: begin
            cosine_reg0 <= 36'sb1111000100101110100101000000111010;
            sine_reg0   <= 36'sb11100001110100010110111101101010101;
        end
        2818: begin
            cosine_reg0 <= 36'sb1111000100000010001111000000101000;
            sine_reg0   <= 36'sb11100001110111010100010100011100001;
        end
        2819: begin
            cosine_reg0 <= 36'sb1111000011010101111000011011001011;
            sine_reg0   <= 36'sb11100001111010010001100010100000011;
        end
        2820: begin
            cosine_reg0 <= 36'sb1111000010101001100001010000100100;
            sine_reg0   <= 36'sb11100001111101001110100111110111001;
        end
        2821: begin
            cosine_reg0 <= 36'sb1111000001111101001001100000110111;
            sine_reg0   <= 36'sb11100010000000001011100100100000011;
        end
        2822: begin
            cosine_reg0 <= 36'sb1111000001010000110001001100000100;
            sine_reg0   <= 36'sb11100010000011001000011000011100000;
        end
        2823: begin
            cosine_reg0 <= 36'sb1111000000100100011000010010001110;
            sine_reg0   <= 36'sb11100010000110000101000011101001111;
        end
        2824: begin
            cosine_reg0 <= 36'sb1110111111110111111110110011010101;
            sine_reg0   <= 36'sb11100010001001000001100110001010000;
        end
        2825: begin
            cosine_reg0 <= 36'sb1110111111001011100100101111011011;
            sine_reg0   <= 36'sb11100010001011111101111111111100000;
        end
        2826: begin
            cosine_reg0 <= 36'sb1110111110011111001010000110100100;
            sine_reg0   <= 36'sb11100010001110111010010000111111111;
        end
        2827: begin
            cosine_reg0 <= 36'sb1110111101110010101110111000101111;
            sine_reg0   <= 36'sb11100010010001110110011001010101101;
        end
        2828: begin
            cosine_reg0 <= 36'sb1110111101000110010011000101111111;
            sine_reg0   <= 36'sb11100010010100110010011000111101001;
        end
        2829: begin
            cosine_reg0 <= 36'sb1110111100011001110110101110010101;
            sine_reg0   <= 36'sb11100010010111101110001111110110000;
        end
        2830: begin
            cosine_reg0 <= 36'sb1110111011101101011001110001110011;
            sine_reg0   <= 36'sb11100010011010101001111110000000100;
        end
        2831: begin
            cosine_reg0 <= 36'sb1110111011000000111100010000011100;
            sine_reg0   <= 36'sb11100010011101100101100011011100010;
        end
        2832: begin
            cosine_reg0 <= 36'sb1110111010010100011110001010010000;
            sine_reg0   <= 36'sb11100010100000100001000000001001010;
        end
        2833: begin
            cosine_reg0 <= 36'sb1110111001100111111111011111010001;
            sine_reg0   <= 36'sb11100010100011011100010100000111011;
        end
        2834: begin
            cosine_reg0 <= 36'sb1110111000111011100000001111100001;
            sine_reg0   <= 36'sb11100010100110010111011111010110100;
        end
        2835: begin
            cosine_reg0 <= 36'sb1110111000001111000000011011000010;
            sine_reg0   <= 36'sb11100010101001010010100001110110100;
        end
        2836: begin
            cosine_reg0 <= 36'sb1110110111100010100000000001110110;
            sine_reg0   <= 36'sb11100010101100001101011011100111010;
        end
        2837: begin
            cosine_reg0 <= 36'sb1110110110110101111111000011111110;
            sine_reg0   <= 36'sb11100010101111001000001100101000101;
        end
        2838: begin
            cosine_reg0 <= 36'sb1110110110001001011101100001011011;
            sine_reg0   <= 36'sb11100010110010000010110100111010101;
        end
        2839: begin
            cosine_reg0 <= 36'sb1110110101011100111011011010010000;
            sine_reg0   <= 36'sb11100010110100111101010100011101001;
        end
        2840: begin
            cosine_reg0 <= 36'sb1110110100110000011000101110011111;
            sine_reg0   <= 36'sb11100010110111110111101011001111111;
        end
        2841: begin
            cosine_reg0 <= 36'sb1110110100000011110101011110001000;
            sine_reg0   <= 36'sb11100010111010110001111001010010111;
        end
        2842: begin
            cosine_reg0 <= 36'sb1110110011010111010001101001001111;
            sine_reg0   <= 36'sb11100010111101101011111110100101111;
        end
        2843: begin
            cosine_reg0 <= 36'sb1110110010101010101101001111110011;
            sine_reg0   <= 36'sb11100011000000100101111011001001000;
        end
        2844: begin
            cosine_reg0 <= 36'sb1110110001111110001000010001111000;
            sine_reg0   <= 36'sb11100011000011011111101110111011111;
        end
        2845: begin
            cosine_reg0 <= 36'sb1110110001010001100010101111011111;
            sine_reg0   <= 36'sb11100011000110011001011001111110101;
        end
        2846: begin
            cosine_reg0 <= 36'sb1110110000100100111100101000101010;
            sine_reg0   <= 36'sb11100011001001010010111100010000111;
        end
        2847: begin
            cosine_reg0 <= 36'sb1110101111111000010101111101011001;
            sine_reg0   <= 36'sb11100011001100001100010101110010111;
        end
        2848: begin
            cosine_reg0 <= 36'sb1110101111001011101110101101110000;
            sine_reg0   <= 36'sb11100011001111000101100110100100001;
        end
        2849: begin
            cosine_reg0 <= 36'sb1110101110011111000110111001110000;
            sine_reg0   <= 36'sb11100011010001111110101110100100110;
        end
        2850: begin
            cosine_reg0 <= 36'sb1110101101110010011110100001011010;
            sine_reg0   <= 36'sb11100011010100110111101101110100101;
        end
        2851: begin
            cosine_reg0 <= 36'sb1110101101000101110101100100110001;
            sine_reg0   <= 36'sb11100011010111110000100100010011101;
        end
        2852: begin
            cosine_reg0 <= 36'sb1110101100011001001100000011110101;
            sine_reg0   <= 36'sb11100011011010101001010010000001100;
        end
        2853: begin
            cosine_reg0 <= 36'sb1110101011101100100001111110101001;
            sine_reg0   <= 36'sb11100011011101100001110110111110011;
        end
        2854: begin
            cosine_reg0 <= 36'sb1110101010111111110111010101001111;
            sine_reg0   <= 36'sb11100011100000011010010011001001111;
        end
        2855: begin
            cosine_reg0 <= 36'sb1110101010010011001100000111100111;
            sine_reg0   <= 36'sb11100011100011010010100110100100001;
        end
        2856: begin
            cosine_reg0 <= 36'sb1110101001100110100000010101110101;
            sine_reg0   <= 36'sb11100011100110001010110001001100111;
        end
        2857: begin
            cosine_reg0 <= 36'sb1110101000111001110011111111111001;
            sine_reg0   <= 36'sb11100011101001000010110011000100000;
        end
        2858: begin
            cosine_reg0 <= 36'sb1110101000001101000111000101110101;
            sine_reg0   <= 36'sb11100011101011111010101100001001100;
        end
        2859: begin
            cosine_reg0 <= 36'sb1110100111100000011001100111101011;
            sine_reg0   <= 36'sb11100011101110110010011100011101010;
        end
        2860: begin
            cosine_reg0 <= 36'sb1110100110110011101011100101011101;
            sine_reg0   <= 36'sb11100011110001101010000011111111000;
        end
        2861: begin
            cosine_reg0 <= 36'sb1110100110000110111100111111001100;
            sine_reg0   <= 36'sb11100011110100100001100010101110111;
        end
        2862: begin
            cosine_reg0 <= 36'sb1110100101011010001101110100111011;
            sine_reg0   <= 36'sb11100011110111011000111000101100100;
        end
        2863: begin
            cosine_reg0 <= 36'sb1110100100101101011110000110101011;
            sine_reg0   <= 36'sb11100011111010010000000101110111111;
        end
        2864: begin
            cosine_reg0 <= 36'sb1110100100000000101101110100011101;
            sine_reg0   <= 36'sb11100011111101000111001010010001000;
        end
        2865: begin
            cosine_reg0 <= 36'sb1110100011010011111100111110010011;
            sine_reg0   <= 36'sb11100011111111111110000101110111101;
        end
        2866: begin
            cosine_reg0 <= 36'sb1110100010100111001011100100010000;
            sine_reg0   <= 36'sb11100100000010110100111000101011101;
        end
        2867: begin
            cosine_reg0 <= 36'sb1110100001111010011001100110010100;
            sine_reg0   <= 36'sb11100100000101101011100010101101000;
        end
        2868: begin
            cosine_reg0 <= 36'sb1110100001001101100111000100100010;
            sine_reg0   <= 36'sb11100100001000100010000011111011101;
        end
        2869: begin
            cosine_reg0 <= 36'sb1110100000100000110011111110111011;
            sine_reg0   <= 36'sb11100100001011011000011100010111011;
        end
        2870: begin
            cosine_reg0 <= 36'sb1110011111110100000000010101100010;
            sine_reg0   <= 36'sb11100100001110001110101100000000000;
        end
        2871: begin
            cosine_reg0 <= 36'sb1110011111000111001100001000010110;
            sine_reg0   <= 36'sb11100100010001000100110010110101101;
        end
        2872: begin
            cosine_reg0 <= 36'sb1110011110011010010111010111011100;
            sine_reg0   <= 36'sb11100100010011111010110000111000000;
        end
        2873: begin
            cosine_reg0 <= 36'sb1110011101101101100010000010110011;
            sine_reg0   <= 36'sb11100100010110110000100110000111000;
        end
        2874: begin
            cosine_reg0 <= 36'sb1110011101000000101100001010011111;
            sine_reg0   <= 36'sb11100100011001100110010010100010100;
        end
        2875: begin
            cosine_reg0 <= 36'sb1110011100010011110101101110100000;
            sine_reg0   <= 36'sb11100100011100011011110110001010101;
        end
        2876: begin
            cosine_reg0 <= 36'sb1110011011100110111110101110111000;
            sine_reg0   <= 36'sb11100100011111010001010000111110111;
        end
        2877: begin
            cosine_reg0 <= 36'sb1110011010111010000111001011101010;
            sine_reg0   <= 36'sb11100100100010000110100010111111100;
        end
        2878: begin
            cosine_reg0 <= 36'sb1110011010001101001111000100110110;
            sine_reg0   <= 36'sb11100100100100111011101100001100010;
        end
        2879: begin
            cosine_reg0 <= 36'sb1110011001100000010110011010011111;
            sine_reg0   <= 36'sb11100100100111110000101100100100111;
        end
        2880: begin
            cosine_reg0 <= 36'sb1110011000110011011101001100100110;
            sine_reg0   <= 36'sb11100100101010100101100100001001100;
        end
        2881: begin
            cosine_reg0 <= 36'sb1110011000000110100011011011001101;
            sine_reg0   <= 36'sb11100100101101011010010010111001111;
        end
        2882: begin
            cosine_reg0 <= 36'sb1110010111011001101001000110010110;
            sine_reg0   <= 36'sb11100100110000001110111000110110000;
        end
        2883: begin
            cosine_reg0 <= 36'sb1110010110101100101110001110000010;
            sine_reg0   <= 36'sb11100100110011000011010101111101101;
        end
        2884: begin
            cosine_reg0 <= 36'sb1110010101111111110010110010010100;
            sine_reg0   <= 36'sb11100100110101110111101010010000110;
        end
        2885: begin
            cosine_reg0 <= 36'sb1110010101010010110110110011001100;
            sine_reg0   <= 36'sb11100100111000101011110101101111010;
        end
        2886: begin
            cosine_reg0 <= 36'sb1110010100100101111010010000101101;
            sine_reg0   <= 36'sb11100100111011011111111000011001000;
        end
        2887: begin
            cosine_reg0 <= 36'sb1110010011111000111101001010111001;
            sine_reg0   <= 36'sb11100100111110010011110010001101110;
        end
        2888: begin
            cosine_reg0 <= 36'sb1110010011001011111111100001110000;
            sine_reg0   <= 36'sb11100101000001000111100011001101110;
        end
        2889: begin
            cosine_reg0 <= 36'sb1110010010011111000001010101010110;
            sine_reg0   <= 36'sb11100101000011111011001011011000100;
        end
        2890: begin
            cosine_reg0 <= 36'sb1110010001110010000010100101101011;
            sine_reg0   <= 36'sb11100101000110101110101010101110001;
        end
        2891: begin
            cosine_reg0 <= 36'sb1110010001000101000011010010110001;
            sine_reg0   <= 36'sb11100101001001100010000001001110100;
        end
        2892: begin
            cosine_reg0 <= 36'sb1110010000011000000011011100101011;
            sine_reg0   <= 36'sb11100101001100010101001110111001011;
        end
        2893: begin
            cosine_reg0 <= 36'sb1110001111101011000011000011011001;
            sine_reg0   <= 36'sb11100101001111001000010011101110110;
        end
        2894: begin
            cosine_reg0 <= 36'sb1110001110111110000010000110111110;
            sine_reg0   <= 36'sb11100101010001111011001111101110101;
        end
        2895: begin
            cosine_reg0 <= 36'sb1110001110010001000000100111011011;
            sine_reg0   <= 36'sb11100101010100101110000010111000101;
        end
        2896: begin
            cosine_reg0 <= 36'sb1110001101100011111110100100110010;
            sine_reg0   <= 36'sb11100101010111100000101101001100111;
        end
        2897: begin
            cosine_reg0 <= 36'sb1110001100110110111011111111000101;
            sine_reg0   <= 36'sb11100101011010010011001110101011010;
        end
        2898: begin
            cosine_reg0 <= 36'sb1110001100001001111000110110010110;
            sine_reg0   <= 36'sb11100101011101000101100111010011100;
        end
        2899: begin
            cosine_reg0 <= 36'sb1110001011011100110101001010100101;
            sine_reg0   <= 36'sb11100101011111110111110111000101100;
        end
        2900: begin
            cosine_reg0 <= 36'sb1110001010101111110000111011110110;
            sine_reg0   <= 36'sb11100101100010101001111110000001011;
        end
        2901: begin
            cosine_reg0 <= 36'sb1110001010000010101100001010001001;
            sine_reg0   <= 36'sb11100101100101011011111100000110111;
        end
        2902: begin
            cosine_reg0 <= 36'sb1110001001010101100110110101100001;
            sine_reg0   <= 36'sb11100101101000001101110001010101111;
        end
        2903: begin
            cosine_reg0 <= 36'sb1110001000101000100000111101111111;
            sine_reg0   <= 36'sb11100101101010111111011101101110010;
        end
        2904: begin
            cosine_reg0 <= 36'sb1110000111111011011010100011100100;
            sine_reg0   <= 36'sb11100101101101110001000001001111111;
        end
        2905: begin
            cosine_reg0 <= 36'sb1110000111001110010011100110010100;
            sine_reg0   <= 36'sb11100101110000100010011011111010111;
        end
        2906: begin
            cosine_reg0 <= 36'sb1110000110100001001100000110001111;
            sine_reg0   <= 36'sb11100101110011010011101101101110111;
        end
        2907: begin
            cosine_reg0 <= 36'sb1110000101110100000100000011010110;
            sine_reg0   <= 36'sb11100101110110000100110110101011110;
        end
        2908: begin
            cosine_reg0 <= 36'sb1110000101000110111011011101101101;
            sine_reg0   <= 36'sb11100101111000110101110110110001101;
        end
        2909: begin
            cosine_reg0 <= 36'sb1110000100011001110010010101010101;
            sine_reg0   <= 36'sb11100101111011100110101110000000010;
        end
        2910: begin
            cosine_reg0 <= 36'sb1110000011101100101000101010001110;
            sine_reg0   <= 36'sb11100101111110010111011100010111101;
        end
        2911: begin
            cosine_reg0 <= 36'sb1110000010111111011110011100011100;
            sine_reg0   <= 36'sb11100110000001001000000001110111100;
        end
        2912: begin
            cosine_reg0 <= 36'sb1110000010010010010011101100000000;
            sine_reg0   <= 36'sb11100110000011111000011110011111110;
        end
        2913: begin
            cosine_reg0 <= 36'sb1110000001100101001000011000111011;
            sine_reg0   <= 36'sb11100110000110101000110010010000100;
        end
        2914: begin
            cosine_reg0 <= 36'sb1110000000110111111100100011001111;
            sine_reg0   <= 36'sb11100110001001011000111101001001011;
        end
        2915: begin
            cosine_reg0 <= 36'sb1110000000001010110000001010111111;
            sine_reg0   <= 36'sb11100110001100001000111111001010011;
        end
        2916: begin
            cosine_reg0 <= 36'sb1101111111011101100011010000001011;
            sine_reg0   <= 36'sb11100110001110111000111000010011100;
        end
        2917: begin
            cosine_reg0 <= 36'sb1101111110110000010101110010110110;
            sine_reg0   <= 36'sb11100110010001101000101000100100100;
        end
        2918: begin
            cosine_reg0 <= 36'sb1101111110000011000111110011000001;
            sine_reg0   <= 36'sb11100110010100011000001111111101010;
        end
        2919: begin
            cosine_reg0 <= 36'sb1101111101010101111001010000101111;
            sine_reg0   <= 36'sb11100110010111000111101110011101111;
        end
        2920: begin
            cosine_reg0 <= 36'sb1101111100101000101010001100000000;
            sine_reg0   <= 36'sb11100110011001110111000100000110000;
        end
        2921: begin
            cosine_reg0 <= 36'sb1101111011111011011010100100110110;
            sine_reg0   <= 36'sb11100110011100100110010000110101101;
        end
        2922: begin
            cosine_reg0 <= 36'sb1101111011001110001010011011010100;
            sine_reg0   <= 36'sb11100110011111010101010100101100101;
        end
        2923: begin
            cosine_reg0 <= 36'sb1101111010100000111001101111011010;
            sine_reg0   <= 36'sb11100110100010000100001111101011000;
        end
        2924: begin
            cosine_reg0 <= 36'sb1101111001110011101000100001001100;
            sine_reg0   <= 36'sb11100110100100110011000001110000100;
        end
        2925: begin
            cosine_reg0 <= 36'sb1101111001000110010110110000101010;
            sine_reg0   <= 36'sb11100110100111100001101010111101000;
        end
        2926: begin
            cosine_reg0 <= 36'sb1101111000011001000100011101110110;
            sine_reg0   <= 36'sb11100110101010010000001011010000101;
        end
        2927: begin
            cosine_reg0 <= 36'sb1101110111101011110001101000110010;
            sine_reg0   <= 36'sb11100110101100111110100010101011000;
        end
        2928: begin
            cosine_reg0 <= 36'sb1101110110111110011110010001100000;
            sine_reg0   <= 36'sb11100110101111101100110001001100010;
        end
        2929: begin
            cosine_reg0 <= 36'sb1101110110010001001010011000000010;
            sine_reg0   <= 36'sb11100110110010011010110110110100001;
        end
        2930: begin
            cosine_reg0 <= 36'sb1101110101100011110101111100011000;
            sine_reg0   <= 36'sb11100110110101001000110011100010100;
        end
        2931: begin
            cosine_reg0 <= 36'sb1101110100110110100000111110100110;
            sine_reg0   <= 36'sb11100110110111110110100111010111011;
        end
        2932: begin
            cosine_reg0 <= 36'sb1101110100001001001011011110101100;
            sine_reg0   <= 36'sb11100110111010100100010010010010100;
        end
        2933: begin
            cosine_reg0 <= 36'sb1101110011011011110101011100101101;
            sine_reg0   <= 36'sb11100110111101010001110100010100000;
        end
        2934: begin
            cosine_reg0 <= 36'sb1101110010101110011110111000101010;
            sine_reg0   <= 36'sb11100110111111111111001101011011100;
        end
        2935: begin
            cosine_reg0 <= 36'sb1101110010000001000111110010100101;
            sine_reg0   <= 36'sb11100111000010101100011101101001001;
        end
        2936: begin
            cosine_reg0 <= 36'sb1101110001010011110000001010011111;
            sine_reg0   <= 36'sb11100111000101011001100100111100110;
        end
        2937: begin
            cosine_reg0 <= 36'sb1101110000100110011000000000011011;
            sine_reg0   <= 36'sb11100111001000000110100011010110000;
        end
        2938: begin
            cosine_reg0 <= 36'sb1101101111111000111111010100011011;
            sine_reg0   <= 36'sb11100111001010110011011000110101001;
        end
        2939: begin
            cosine_reg0 <= 36'sb1101101111001011100110000110011111;
            sine_reg0   <= 36'sb11100111001101100000000101011001110;
        end
        2940: begin
            cosine_reg0 <= 36'sb1101101110011110001100010110101010;
            sine_reg0   <= 36'sb11100111010000001100101001000100000;
        end
        2941: begin
            cosine_reg0 <= 36'sb1101101101110000110010000100111101;
            sine_reg0   <= 36'sb11100111010010111001000011110011101;
        end
        2942: begin
            cosine_reg0 <= 36'sb1101101101000011010111010001011011;
            sine_reg0   <= 36'sb11100111010101100101010101101000100;
        end
        2943: begin
            cosine_reg0 <= 36'sb1101101100010101111011111100000100;
            sine_reg0   <= 36'sb11100111011000010001011110100010101;
        end
        2944: begin
            cosine_reg0 <= 36'sb1101101011101000100000000100111100;
            sine_reg0   <= 36'sb11100111011010111101011110100001110;
        end
        2945: begin
            cosine_reg0 <= 36'sb1101101010111011000011101100000011;
            sine_reg0   <= 36'sb11100111011101101001010101100110000;
        end
        2946: begin
            cosine_reg0 <= 36'sb1101101010001101100110110001011010;
            sine_reg0   <= 36'sb11100111100000010101000011101111000;
        end
        2947: begin
            cosine_reg0 <= 36'sb1101101001100000001001010101000101;
            sine_reg0   <= 36'sb11100111100011000000101000111100111;
        end
        2948: begin
            cosine_reg0 <= 36'sb1101101000110010101011010111000101;
            sine_reg0   <= 36'sb11100111100101101100000101001111100;
        end
        2949: begin
            cosine_reg0 <= 36'sb1101101000000101001100110111011011;
            sine_reg0   <= 36'sb11100111101000010111011000100110100;
        end
        2950: begin
            cosine_reg0 <= 36'sb1101100111010111101101110110001010;
            sine_reg0   <= 36'sb11100111101011000010100011000010001;
        end
        2951: begin
            cosine_reg0 <= 36'sb1101100110101010001110010011010010;
            sine_reg0   <= 36'sb11100111101101101101100100100010001;
        end
        2952: begin
            cosine_reg0 <= 36'sb1101100101111100101110001110110110;
            sine_reg0   <= 36'sb11100111110000011000011101000110011;
        end
        2953: begin
            cosine_reg0 <= 36'sb1101100101001111001101101000111000;
            sine_reg0   <= 36'sb11100111110011000011001100101110110;
        end
        2954: begin
            cosine_reg0 <= 36'sb1101100100100001101100100001011000;
            sine_reg0   <= 36'sb11100111110101101101110011011011001;
        end
        2955: begin
            cosine_reg0 <= 36'sb1101100011110100001010111000011010;
            sine_reg0   <= 36'sb11100111111000011000010001001011101;
        end
        2956: begin
            cosine_reg0 <= 36'sb1101100011000110101000101101111111;
            sine_reg0   <= 36'sb11100111111011000010100101111111111;
        end
        2957: begin
            cosine_reg0 <= 36'sb1101100010011001000110000010001000;
            sine_reg0   <= 36'sb11100111111101101100110001110111111;
        end
        2958: begin
            cosine_reg0 <= 36'sb1101100001101011100010110100110111;
            sine_reg0   <= 36'sb11101000000000010110110100110011101;
        end
        2959: begin
            cosine_reg0 <= 36'sb1101100000111101111111000110001110;
            sine_reg0   <= 36'sb11101000000011000000101110110010110;
        end
        2960: begin
            cosine_reg0 <= 36'sb1101100000010000011010110110001111;
            sine_reg0   <= 36'sb11101000000101101010011111110101100;
        end
        2961: begin
            cosine_reg0 <= 36'sb1101011111100010110110000100111100;
            sine_reg0   <= 36'sb11101000001000010100000111111011100;
        end
        2962: begin
            cosine_reg0 <= 36'sb1101011110110101010000110010010110;
            sine_reg0   <= 36'sb11101000001010111101100111000100110;
        end
        2963: begin
            cosine_reg0 <= 36'sb1101011110000111101010111110011111;
            sine_reg0   <= 36'sb11101000001101100110111101010001001;
        end
        2964: begin
            cosine_reg0 <= 36'sb1101011101011010000100101001011001;
            sine_reg0   <= 36'sb11101000010000010000001010100000101;
        end
        2965: begin
            cosine_reg0 <= 36'sb1101011100101100011101110011000101;
            sine_reg0   <= 36'sb11101000010010111001001110110011000;
        end
        2966: begin
            cosine_reg0 <= 36'sb1101011011111110110110011011100110;
            sine_reg0   <= 36'sb11101000010101100010001010001000001;
        end
        2967: begin
            cosine_reg0 <= 36'sb1101011011010001001110100010111101;
            sine_reg0   <= 36'sb11101000011000001010111100100000001;
        end
        2968: begin
            cosine_reg0 <= 36'sb1101011010100011100110001001001011;
            sine_reg0   <= 36'sb11101000011010110011100101111010110;
        end
        2969: begin
            cosine_reg0 <= 36'sb1101011001110101111101001110010011;
            sine_reg0   <= 36'sb11101000011101011100000110010111110;
        end
        2970: begin
            cosine_reg0 <= 36'sb1101011001001000010011110010010111;
            sine_reg0   <= 36'sb11101000100000000100011101110111011;
        end
        2971: begin
            cosine_reg0 <= 36'sb1101011000011010101001110101011000;
            sine_reg0   <= 36'sb11101000100010101100101100011001001;
        end
        2972: begin
            cosine_reg0 <= 36'sb1101010111101100111111010111010111;
            sine_reg0   <= 36'sb11101000100101010100110001111101010;
        end
        2973: begin
            cosine_reg0 <= 36'sb1101010110111111010100011000010111;
            sine_reg0   <= 36'sb11101000100111111100101110100011100;
        end
        2974: begin
            cosine_reg0 <= 36'sb1101010110010001101000111000011010;
            sine_reg0   <= 36'sb11101000101010100100100010001011110;
        end
        2975: begin
            cosine_reg0 <= 36'sb1101010101100011111100110111100001;
            sine_reg0   <= 36'sb11101000101101001100001100110101111;
        end
        2976: begin
            cosine_reg0 <= 36'sb1101010100110110010000010101101101;
            sine_reg0   <= 36'sb11101000101111110011101110100001111;
        end
        2977: begin
            cosine_reg0 <= 36'sb1101010100001000100011010011000010;
            sine_reg0   <= 36'sb11101000110010011011000111001111100;
        end
        2978: begin
            cosine_reg0 <= 36'sb1101010011011010110101101111011111;
            sine_reg0   <= 36'sb11101000110101000010010110111110111;
        end
        2979: begin
            cosine_reg0 <= 36'sb1101010010101101000111101011001000;
            sine_reg0   <= 36'sb11101000110111101001011101101111101;
        end
        2980: begin
            cosine_reg0 <= 36'sb1101010001111111011001000101111110;
            sine_reg0   <= 36'sb11101000111010010000011011100001111;
        end
        2981: begin
            cosine_reg0 <= 36'sb1101010001010001101010000000000011;
            sine_reg0   <= 36'sb11101000111100110111010000010101100;
        end
        2982: begin
            cosine_reg0 <= 36'sb1101010000100011111010011001011000;
            sine_reg0   <= 36'sb11101000111111011101111100001010010;
        end
        2983: begin
            cosine_reg0 <= 36'sb1101001111110110001010010010000000;
            sine_reg0   <= 36'sb11101001000010000100011111000000001;
        end
        2984: begin
            cosine_reg0 <= 36'sb1101001111001000011001101001111011;
            sine_reg0   <= 36'sb11101001000100101010111000110111001;
        end
        2985: begin
            cosine_reg0 <= 36'sb1101001110011010101000100001001100;
            sine_reg0   <= 36'sb11101001000111010001001001101110111;
        end
        2986: begin
            cosine_reg0 <= 36'sb1101001101101100110110110111110101;
            sine_reg0   <= 36'sb11101001001001110111010001100111100;
        end
        2987: begin
            cosine_reg0 <= 36'sb1101001100111111000100101101110111;
            sine_reg0   <= 36'sb11101001001100011101010000100000111;
        end
        2988: begin
            cosine_reg0 <= 36'sb1101001100010001010010000011010100;
            sine_reg0   <= 36'sb11101001001111000011000110011010111;
        end
        2989: begin
            cosine_reg0 <= 36'sb1101001011100011011110111000001111;
            sine_reg0   <= 36'sb11101001010001101000110011010101011;
        end
        2990: begin
            cosine_reg0 <= 36'sb1101001010110101101011001100100111;
            sine_reg0   <= 36'sb11101001010100001110010111010000010;
        end
        2991: begin
            cosine_reg0 <= 36'sb1101001010000111110111000000100000;
            sine_reg0   <= 36'sb11101001010110110011110010001011100;
        end
        2992: begin
            cosine_reg0 <= 36'sb1101001001011010000010010011111011;
            sine_reg0   <= 36'sb11101001011001011001000100000110111;
        end
        2993: begin
            cosine_reg0 <= 36'sb1101001000101100001101000110111011;
            sine_reg0   <= 36'sb11101001011011111110001101000010100;
        end
        2994: begin
            cosine_reg0 <= 36'sb1101000111111110010111011001011111;
            sine_reg0   <= 36'sb11101001011110100011001100111110000;
        end
        2995: begin
            cosine_reg0 <= 36'sb1101000111010000100001001011101100;
            sine_reg0   <= 36'sb11101001100001001000000011111001100;
        end
        2996: begin
            cosine_reg0 <= 36'sb1101000110100010101010011101100001;
            sine_reg0   <= 36'sb11101001100011101100110001110100111;
        end
        2997: begin
            cosine_reg0 <= 36'sb1101000101110100110011001111000001;
            sine_reg0   <= 36'sb11101001100110010001010110101111111;
        end
        2998: begin
            cosine_reg0 <= 36'sb1101000101000110111011100000001111;
            sine_reg0   <= 36'sb11101001101000110101110010101010100;
        end
        2999: begin
            cosine_reg0 <= 36'sb1101000100011001000011010001001010;
            sine_reg0   <= 36'sb11101001101011011010000101100100101;
        end
        3000: begin
            cosine_reg0 <= 36'sb1101000011101011001010100001110110;
            sine_reg0   <= 36'sb11101001101101111110001111011110010;
        end
        3001: begin
            cosine_reg0 <= 36'sb1101000010111101010001010010010100;
            sine_reg0   <= 36'sb11101001110000100010010000010111001;
        end
        3002: begin
            cosine_reg0 <= 36'sb1101000010001111010111100010100110;
            sine_reg0   <= 36'sb11101001110011000110001000001111010;
        end
        3003: begin
            cosine_reg0 <= 36'sb1101000001100001011101010010101110;
            sine_reg0   <= 36'sb11101001110101101001110111000110101;
        end
        3004: begin
            cosine_reg0 <= 36'sb1101000000110011100010100010101100;
            sine_reg0   <= 36'sb11101001111000001101011100111100111;
        end
        3005: begin
            cosine_reg0 <= 36'sb1101000000000101100111010010100100;
            sine_reg0   <= 36'sb11101001111010110000111001110010001;
        end
        3006: begin
            cosine_reg0 <= 36'sb1100111111010111101011100010010111;
            sine_reg0   <= 36'sb11101001111101010100001101100110001;
        end
        3007: begin
            cosine_reg0 <= 36'sb1100111110101001101111010010000111;
            sine_reg0   <= 36'sb11101001111111110111011000011000111;
        end
        3008: begin
            cosine_reg0 <= 36'sb1100111101111011110010100001110101;
            sine_reg0   <= 36'sb11101010000010011010011010001010011;
        end
        3009: begin
            cosine_reg0 <= 36'sb1100111101001101110101010001100011;
            sine_reg0   <= 36'sb11101010000100111101010010111010010;
        end
        3010: begin
            cosine_reg0 <= 36'sb1100111100011111110111100001010011;
            sine_reg0   <= 36'sb11101010000111100000000010101000101;
        end
        3011: begin
            cosine_reg0 <= 36'sb1100111011110001111001010001000111;
            sine_reg0   <= 36'sb11101010001010000010101001010101011;
        end
        3012: begin
            cosine_reg0 <= 36'sb1100111011000011111010100001000001;
            sine_reg0   <= 36'sb11101010001100100101000111000000011;
        end
        3013: begin
            cosine_reg0 <= 36'sb1100111010010101111011010001000001;
            sine_reg0   <= 36'sb11101010001111000111011011101001100;
        end
        3014: begin
            cosine_reg0 <= 36'sb1100111001100111111011100001001011;
            sine_reg0   <= 36'sb11101010010001101001100111010000101;
        end
        3015: begin
            cosine_reg0 <= 36'sb1100111000111001111011010001100000;
            sine_reg0   <= 36'sb11101010010100001011101001110101110;
        end
        3016: begin
            cosine_reg0 <= 36'sb1100111000001011111010100010000001;
            sine_reg0   <= 36'sb11101010010110101101100011011000101;
        end
        3017: begin
            cosine_reg0 <= 36'sb1100110111011101111001010010110001;
            sine_reg0   <= 36'sb11101010011001001111010011111001011;
        end
        3018: begin
            cosine_reg0 <= 36'sb1100110110101111110111100011110001;
            sine_reg0   <= 36'sb11101010011011110000111011010111110;
        end
        3019: begin
            cosine_reg0 <= 36'sb1100110110000001110101010101000011;
            sine_reg0   <= 36'sb11101010011110010010011001110011101;
        end
        3020: begin
            cosine_reg0 <= 36'sb1100110101010011110010100110101001;
            sine_reg0   <= 36'sb11101010100000110011101111001101000;
        end
        3021: begin
            cosine_reg0 <= 36'sb1100110100100101101111011000100100;
            sine_reg0   <= 36'sb11101010100011010100111011100011110;
        end
        3022: begin
            cosine_reg0 <= 36'sb1100110011110111101011101010110110;
            sine_reg0   <= 36'sb11101010100101110101111110110111110;
        end
        3023: begin
            cosine_reg0 <= 36'sb1100110011001001100111011101100010;
            sine_reg0   <= 36'sb11101010101000010110111001001000111;
        end
        3024: begin
            cosine_reg0 <= 36'sb1100110010011011100010110000101000;
            sine_reg0   <= 36'sb11101010101010110111101010010111001;
        end
        3025: begin
            cosine_reg0 <= 36'sb1100110001101101011101100100001011;
            sine_reg0   <= 36'sb11101010101101011000010010100010011;
        end
        3026: begin
            cosine_reg0 <= 36'sb1100110000111111010111111000001100;
            sine_reg0   <= 36'sb11101010101111111000110001101010100;
        end
        3027: begin
            cosine_reg0 <= 36'sb1100110000010001010001101100101101;
            sine_reg0   <= 36'sb11101010110010011001000111101111011;
        end
        3028: begin
            cosine_reg0 <= 36'sb1100101111100011001011000001110001;
            sine_reg0   <= 36'sb11101010110100111001010100110001000;
        end
        3029: begin
            cosine_reg0 <= 36'sb1100101110110101000011110111011000;
            sine_reg0   <= 36'sb11101010110111011001011000101111001;
        end
        3030: begin
            cosine_reg0 <= 36'sb1100101110000110111100001101100100;
            sine_reg0   <= 36'sb11101010111001111001010011101001110;
        end
        3031: begin
            cosine_reg0 <= 36'sb1100101101011000110100000100011000;
            sine_reg0   <= 36'sb11101010111100011001000101100000110;
        end
        3032: begin
            cosine_reg0 <= 36'sb1100101100101010101011011011110101;
            sine_reg0   <= 36'sb11101010111110111000101110010100001;
        end
        3033: begin
            cosine_reg0 <= 36'sb1100101011111100100010010011111101;
            sine_reg0   <= 36'sb11101011000001011000001110000011110;
        end
        3034: begin
            cosine_reg0 <= 36'sb1100101011001110011000101100110001;
            sine_reg0   <= 36'sb11101011000011110111100100101111011;
        end
        3035: begin
            cosine_reg0 <= 36'sb1100101010100000001110100110010100;
            sine_reg0   <= 36'sb11101011000110010110110010010111000;
        end
        3036: begin
            cosine_reg0 <= 36'sb1100101001110010000100000000100111;
            sine_reg0   <= 36'sb11101011001000110101110110111010101;
        end
        3037: begin
            cosine_reg0 <= 36'sb1100101001000011111000111011101011;
            sine_reg0   <= 36'sb11101011001011010100110010011010000;
        end
        3038: begin
            cosine_reg0 <= 36'sb1100101000010101101101010111100100;
            sine_reg0   <= 36'sb11101011001101110011100100110101001;
        end
        3039: begin
            cosine_reg0 <= 36'sb1100100111100111100001010100010010;
            sine_reg0   <= 36'sb11101011010000010010001110001011111;
        end
        3040: begin
            cosine_reg0 <= 36'sb1100100110111001010100110001110111;
            sine_reg0   <= 36'sb11101011010010110000101110011110010;
        end
        3041: begin
            cosine_reg0 <= 36'sb1100100110001011000111110000010110;
            sine_reg0   <= 36'sb11101011010101001111000101101011111;
        end
        3042: begin
            cosine_reg0 <= 36'sb1100100101011100111010001111101111;
            sine_reg0   <= 36'sb11101011010111101101010011110101000;
        end
        3043: begin
            cosine_reg0 <= 36'sb1100100100101110101100010000000101;
            sine_reg0   <= 36'sb11101011011010001011011000111001010;
        end
        3044: begin
            cosine_reg0 <= 36'sb1100100100000000011101110001011001;
            sine_reg0   <= 36'sb11101011011100101001010100111000110;
        end
        3045: begin
            cosine_reg0 <= 36'sb1100100011010010001110110011101101;
            sine_reg0   <= 36'sb11101011011111000111000111110011010;
        end
        3046: begin
            cosine_reg0 <= 36'sb1100100010100011111111010111000100;
            sine_reg0   <= 36'sb11101011100001100100110001101000110;
        end
        3047: begin
            cosine_reg0 <= 36'sb1100100001110101101111011011011110;
            sine_reg0   <= 36'sb11101011100100000010010010011001001;
        end
        3048: begin
            cosine_reg0 <= 36'sb1100100001000111011111000000111110;
            sine_reg0   <= 36'sb11101011100110011111101010000100010;
        end
        3049: begin
            cosine_reg0 <= 36'sb1100100000011001001110000111100101;
            sine_reg0   <= 36'sb11101011101000111100111000101010000;
        end
        3050: begin
            cosine_reg0 <= 36'sb1100011111101010111100101111010101;
            sine_reg0   <= 36'sb11101011101011011001111110001010100;
        end
        3051: begin
            cosine_reg0 <= 36'sb1100011110111100101010111000010000;
            sine_reg0   <= 36'sb11101011101101110110111010100101011;
        end
        3052: begin
            cosine_reg0 <= 36'sb1100011110001110011000100010010111;
            sine_reg0   <= 36'sb11101011110000010011101101111010101;
        end
        3053: begin
            cosine_reg0 <= 36'sb1100011101100000000101101101101110;
            sine_reg0   <= 36'sb11101011110010110000011000001010001;
        end
        3054: begin
            cosine_reg0 <= 36'sb1100011100110001110010011010010100;
            sine_reg0   <= 36'sb11101011110101001100111001010011111;
        end
        3055: begin
            cosine_reg0 <= 36'sb1100011100000011011110101000001100;
            sine_reg0   <= 36'sb11101011110111101001010001010111110;
        end
        3056: begin
            cosine_reg0 <= 36'sb1100011011010101001010010111011001;
            sine_reg0   <= 36'sb11101011111010000101100000010101101;
        end
        3057: begin
            cosine_reg0 <= 36'sb1100011010100110110101100111111011;
            sine_reg0   <= 36'sb11101011111100100001100110001101100;
        end
        3058: begin
            cosine_reg0 <= 36'sb1100011001111000100000011001110100;
            sine_reg0   <= 36'sb11101011111110111101100010111111001;
        end
        3059: begin
            cosine_reg0 <= 36'sb1100011001001010001010101101000110;
            sine_reg0   <= 36'sb11101100000001011001010110101010100;
        end
        3060: begin
            cosine_reg0 <= 36'sb1100011000011011110100100001110100;
            sine_reg0   <= 36'sb11101100000011110101000001001111100;
        end
        3061: begin
            cosine_reg0 <= 36'sb1100010111101101011101110111111110;
            sine_reg0   <= 36'sb11101100000110010000100010101110000;
        end
        3062: begin
            cosine_reg0 <= 36'sb1100010110111111000110101111100110;
            sine_reg0   <= 36'sb11101100001000101011111011000110000;
        end
        3063: begin
            cosine_reg0 <= 36'sb1100010110010000101111001000101111;
            sine_reg0   <= 36'sb11101100001011000111001010010111011;
        end
        3064: begin
            cosine_reg0 <= 36'sb1100010101100010010111000011011010;
            sine_reg0   <= 36'sb11101100001101100010010000100010000;
        end
        3065: begin
            cosine_reg0 <= 36'sb1100010100110011111110011111101001;
            sine_reg0   <= 36'sb11101100001111111101001101100101111;
        end
        3066: begin
            cosine_reg0 <= 36'sb1100010100000101100101011101011110;
            sine_reg0   <= 36'sb11101100010010011000000001100010110;
        end
        3067: begin
            cosine_reg0 <= 36'sb1100010011010111001011111100111010;
            sine_reg0   <= 36'sb11101100010100110010101100011000101;
        end
        3068: begin
            cosine_reg0 <= 36'sb1100010010101000110001111101111111;
            sine_reg0   <= 36'sb11101100010111001101001110000111011;
        end
        3069: begin
            cosine_reg0 <= 36'sb1100010001111010010111100000110000;
            sine_reg0   <= 36'sb11101100011001100111100110101110111;
        end
        3070: begin
            cosine_reg0 <= 36'sb1100010001001011111100100101001101;
            sine_reg0   <= 36'sb11101100011100000001110110001111010;
        end
        3071: begin
            cosine_reg0 <= 36'sb1100010000011101100001001011011001;
            sine_reg0   <= 36'sb11101100011110011011111100101000001;
        end
        3072: begin
            cosine_reg0 <= 36'sb1100001111101111000101010011010101;
            sine_reg0   <= 36'sb11101100100000110101111001111001100;
        end
        3073: begin
            cosine_reg0 <= 36'sb1100001111000000101000111101000100;
            sine_reg0   <= 36'sb11101100100011001111101110000011010;
        end
        3074: begin
            cosine_reg0 <= 36'sb1100001110010010001100001000100111;
            sine_reg0   <= 36'sb11101100100101101001011001000101100;
        end
        3075: begin
            cosine_reg0 <= 36'sb1100001101100011101110110101111111;
            sine_reg0   <= 36'sb11101100101000000010111010111111111;
        end
        3076: begin
            cosine_reg0 <= 36'sb1100001100110101010001000101001111;
            sine_reg0   <= 36'sb11101100101010011100010011110010011;
        end
        3077: begin
            cosine_reg0 <= 36'sb1100001100000110110010110110011000;
            sine_reg0   <= 36'sb11101100101100110101100011011101000;
        end
        3078: begin
            cosine_reg0 <= 36'sb1100001011011000010100001001011101;
            sine_reg0   <= 36'sb11101100101111001110101001111111101;
        end
        3079: begin
            cosine_reg0 <= 36'sb1100001010101001110100111110011110;
            sine_reg0   <= 36'sb11101100110001100111100111011010000;
        end
        3080: begin
            cosine_reg0 <= 36'sb1100001001111011010101010101011110;
            sine_reg0   <= 36'sb11101100110100000000011011101100010;
        end
        3081: begin
            cosine_reg0 <= 36'sb1100001001001100110101001110011111;
            sine_reg0   <= 36'sb11101100110110011001000110110110001;
        end
        3082: begin
            cosine_reg0 <= 36'sb1100001000011110010100101001100010;
            sine_reg0   <= 36'sb11101100111000110001101000110111101;
        end
        3083: begin
            cosine_reg0 <= 36'sb1100000111101111110011100110101001;
            sine_reg0   <= 36'sb11101100111011001010000001110000101;
        end
        3084: begin
            cosine_reg0 <= 36'sb1100000111000001010010000101110110;
            sine_reg0   <= 36'sb11101100111101100010010001100001001;
        end
        3085: begin
            cosine_reg0 <= 36'sb1100000110010010110000000111001011;
            sine_reg0   <= 36'sb11101100111111111010011000001000111;
        end
        3086: begin
            cosine_reg0 <= 36'sb1100000101100100001101101010101001;
            sine_reg0   <= 36'sb11101101000010010010010101100111111;
        end
        3087: begin
            cosine_reg0 <= 36'sb1100000100110101101010110000010011;
            sine_reg0   <= 36'sb11101101000100101010001001111101111;
        end
        3088: begin
            cosine_reg0 <= 36'sb1100000100000111000111011000001001;
            sine_reg0   <= 36'sb11101101000111000001110101001011001;
        end
        3089: begin
            cosine_reg0 <= 36'sb1100000011011000100011100010001111;
            sine_reg0   <= 36'sb11101101001001011001010111001111010;
        end
        3090: begin
            cosine_reg0 <= 36'sb1100000010101001111111001110100101;
            sine_reg0   <= 36'sb11101101001011110000110000001010001;
        end
        3091: begin
            cosine_reg0 <= 36'sb1100000001111011011010011101001110;
            sine_reg0   <= 36'sb11101101001110000111111111111011111;
        end
        3092: begin
            cosine_reg0 <= 36'sb1100000001001100110101001110001011;
            sine_reg0   <= 36'sb11101101010000011111000110100100011;
        end
        3093: begin
            cosine_reg0 <= 36'sb1100000000011110001111100001011110;
            sine_reg0   <= 36'sb11101101010010110110000100000011011;
        end
        3094: begin
            cosine_reg0 <= 36'sb1011111111101111101001010111001001;
            sine_reg0   <= 36'sb11101101010101001100111000011000111;
        end
        3095: begin
            cosine_reg0 <= 36'sb1011111111000001000010101111001110;
            sine_reg0   <= 36'sb11101101010111100011100011100100111;
        end
        3096: begin
            cosine_reg0 <= 36'sb1011111110010010011011101001101110;
            sine_reg0   <= 36'sb11101101011001111010000101100111001;
        end
        3097: begin
            cosine_reg0 <= 36'sb1011111101100011110100000110101011;
            sine_reg0   <= 36'sb11101101011100010000011110011111101;
        end
        3098: begin
            cosine_reg0 <= 36'sb1011111100110101001100000110001000;
            sine_reg0   <= 36'sb11101101011110100110101110001110001;
        end
        3099: begin
            cosine_reg0 <= 36'sb1011111100000110100011101000000101;
            sine_reg0   <= 36'sb11101101100000111100110100110010111;
        end
        3100: begin
            cosine_reg0 <= 36'sb1011111011010111111010101100100101;
            sine_reg0   <= 36'sb11101101100011010010110010001101100;
        end
        3101: begin
            cosine_reg0 <= 36'sb1011111010101001010001010011101001;
            sine_reg0   <= 36'sb11101101100101101000100110011101111;
        end
        3102: begin
            cosine_reg0 <= 36'sb1011111001111010100111011101010100;
            sine_reg0   <= 36'sb11101101100111111110010001100100001;
        end
        3103: begin
            cosine_reg0 <= 36'sb1011111001001011111101001001100111;
            sine_reg0   <= 36'sb11101101101010010011110011100000001;
        end
        3104: begin
            cosine_reg0 <= 36'sb1011111000011101010010011000100011;
            sine_reg0   <= 36'sb11101101101100101001001100010001101;
        end
        3105: begin
            cosine_reg0 <= 36'sb1011110111101110100111001010001100;
            sine_reg0   <= 36'sb11101101101110111110011011111000110;
        end
        3106: begin
            cosine_reg0 <= 36'sb1011110110111111111011011110100001;
            sine_reg0   <= 36'sb11101101110001010011100010010101001;
        end
        3107: begin
            cosine_reg0 <= 36'sb1011110110010001001111010101100110;
            sine_reg0   <= 36'sb11101101110011101000011111100110111;
        end
        3108: begin
            cosine_reg0 <= 36'sb1011110101100010100010101111011100;
            sine_reg0   <= 36'sb11101101110101111101010011101110000;
        end
        3109: begin
            cosine_reg0 <= 36'sb1011110100110011110101101100000101;
            sine_reg0   <= 36'sb11101101111000010001111110101010001;
        end
        3110: begin
            cosine_reg0 <= 36'sb1011110100000101001000001011100010;
            sine_reg0   <= 36'sb11101101111010100110100000011011011;
        end
        3111: begin
            cosine_reg0 <= 36'sb1011110011010110011010001101110110;
            sine_reg0   <= 36'sb11101101111100111010111001000001100;
        end
        3112: begin
            cosine_reg0 <= 36'sb1011110010100111101011110011000010;
            sine_reg0   <= 36'sb11101101111111001111001000011100100;
        end
        3113: begin
            cosine_reg0 <= 36'sb1011110001111000111100111011001000;
            sine_reg0   <= 36'sb11101110000001100011001110101100011;
        end
        3114: begin
            cosine_reg0 <= 36'sb1011110001001010001101100110001010;
            sine_reg0   <= 36'sb11101110000011110111001011110001000;
        end
        3115: begin
            cosine_reg0 <= 36'sb1011110000011011011101110100001010;
            sine_reg0   <= 36'sb11101110000110001010111111101010001;
        end
        3116: begin
            cosine_reg0 <= 36'sb1011101111101100101101100101001001;
            sine_reg0   <= 36'sb11101110001000011110101010010111110;
        end
        3117: begin
            cosine_reg0 <= 36'sb1011101110111101111100111001001001;
            sine_reg0   <= 36'sb11101110001010110010001011111001111;
        end
        3118: begin
            cosine_reg0 <= 36'sb1011101110001111001011110000001101;
            sine_reg0   <= 36'sb11101110001101000101100100010000011;
        end
        3119: begin
            cosine_reg0 <= 36'sb1011101101100000011010001010010101;
            sine_reg0   <= 36'sb11101110001111011000110011011011000;
        end
        3120: begin
            cosine_reg0 <= 36'sb1011101100110001101000000111100100;
            sine_reg0   <= 36'sb11101110010001101011111001011001111;
        end
        3121: begin
            cosine_reg0 <= 36'sb1011101100000010110101100111111100;
            sine_reg0   <= 36'sb11101110010011111110110110001100111;
        end
        3122: begin
            cosine_reg0 <= 36'sb1011101011010100000010101011011101;
            sine_reg0   <= 36'sb11101110010110010001101001110011110;
        end
        3123: begin
            cosine_reg0 <= 36'sb1011101010100101001111010010001011;
            sine_reg0   <= 36'sb11101110011000100100010100001110101;
        end
        3124: begin
            cosine_reg0 <= 36'sb1011101001110110011011011100000111;
            sine_reg0   <= 36'sb11101110011010110110110101011101010;
        end
        3125: begin
            cosine_reg0 <= 36'sb1011101001000111100111001001010010;
            sine_reg0   <= 36'sb11101110011101001001001101011111101;
        end
        3126: begin
            cosine_reg0 <= 36'sb1011101000011000110010011001101111;
            sine_reg0   <= 36'sb11101110011111011011011100010101101;
        end
        3127: begin
            cosine_reg0 <= 36'sb1011100111101001111101001101011111;
            sine_reg0   <= 36'sb11101110100001101101100001111111010;
        end
        3128: begin
            cosine_reg0 <= 36'sb1011100110111011000111100100100100;
            sine_reg0   <= 36'sb11101110100011111111011110011100010;
        end
        3129: begin
            cosine_reg0 <= 36'sb1011100110001100010001011111000001;
            sine_reg0   <= 36'sb11101110100110010001010001101100101;
        end
        3130: begin
            cosine_reg0 <= 36'sb1011100101011101011010111100110101;
            sine_reg0   <= 36'sb11101110101000100010111011110000010;
        end
        3131: begin
            cosine_reg0 <= 36'sb1011100100101110100011111110000101;
            sine_reg0   <= 36'sb11101110101010110100011100100111001;
        end
        3132: begin
            cosine_reg0 <= 36'sb1011100011111111101100100010110001;
            sine_reg0   <= 36'sb11101110101101000101110100010001001;
        end
        3133: begin
            cosine_reg0 <= 36'sb1011100011010000110100101010111010;
            sine_reg0   <= 36'sb11101110101111010111000010101110001;
        end
        3134: begin
            cosine_reg0 <= 36'sb1011100010100001111100010110100100;
            sine_reg0   <= 36'sb11101110110001101000000111111110000;
        end
        3135: begin
            cosine_reg0 <= 36'sb1011100001110011000011100101110000;
            sine_reg0   <= 36'sb11101110110011111001000100000000110;
        end
        3136: begin
            cosine_reg0 <= 36'sb1011100001000100001010011000011111;
            sine_reg0   <= 36'sb11101110110110001001110110110110010;
        end
        3137: begin
            cosine_reg0 <= 36'sb1011100000010101010000101110110011;
            sine_reg0   <= 36'sb11101110111000011010100000011110100;
        end
        3138: begin
            cosine_reg0 <= 36'sb1011011111100110010110101000101111;
            sine_reg0   <= 36'sb11101110111010101011000000111001010;
        end
        3139: begin
            cosine_reg0 <= 36'sb1011011110110111011100000110010100;
            sine_reg0   <= 36'sb11101110111100111011011000000110100;
        end
        3140: begin
            cosine_reg0 <= 36'sb1011011110001000100001000111100011;
            sine_reg0   <= 36'sb11101110111111001011100110000110010;
        end
        3141: begin
            cosine_reg0 <= 36'sb1011011101011001100101101100011111;
            sine_reg0   <= 36'sb11101111000001011011101010111000010;
        end
        3142: begin
            cosine_reg0 <= 36'sb1011011100101010101001110101001010;
            sine_reg0   <= 36'sb11101111000011101011100110011100100;
        end
        3143: begin
            cosine_reg0 <= 36'sb1011011011111011101101100001100100;
            sine_reg0   <= 36'sb11101111000101111011011000110010111;
        end
        3144: begin
            cosine_reg0 <= 36'sb1011011011001100110000110001110001;
            sine_reg0   <= 36'sb11101111001000001011000001111011010;
        end
        3145: begin
            cosine_reg0 <= 36'sb1011011010011101110011100101110001;
            sine_reg0   <= 36'sb11101111001010011010100001110101110;
        end
        3146: begin
            cosine_reg0 <= 36'sb1011011001101110110101111101101000;
            sine_reg0   <= 36'sb11101111001100101001111000100010000;
        end
        3147: begin
            cosine_reg0 <= 36'sb1011011000111111110111111001010101;
            sine_reg0   <= 36'sb11101111001110111001000110000000001;
        end
        3148: begin
            cosine_reg0 <= 36'sb1011011000010000111001011000111100;
            sine_reg0   <= 36'sb11101111010001001000001010010000000;
        end
        3149: begin
            cosine_reg0 <= 36'sb1011010111100001111010011100011110;
            sine_reg0   <= 36'sb11101111010011010111000101010001100;
        end
        3150: begin
            cosine_reg0 <= 36'sb1011010110110010111011000011111101;
            sine_reg0   <= 36'sb11101111010101100101110111000100100;
        end
        3151: begin
            cosine_reg0 <= 36'sb1011010110000011111011001111011010;
            sine_reg0   <= 36'sb11101111010111110100011111101001000;
        end
        3152: begin
            cosine_reg0 <= 36'sb1011010101010100111010111110111001;
            sine_reg0   <= 36'sb11101111011010000010111110111110111;
        end
        3153: begin
            cosine_reg0 <= 36'sb1011010100100101111010010010011001;
            sine_reg0   <= 36'sb11101111011100010001010101000110000;
        end
        3154: begin
            cosine_reg0 <= 36'sb1011010011110110111001001001111110;
            sine_reg0   <= 36'sb11101111011110011111100001111110010;
        end
        3155: begin
            cosine_reg0 <= 36'sb1011010011000111110111100101101000;
            sine_reg0   <= 36'sb11101111100000101101100101100111110;
        end
        3156: begin
            cosine_reg0 <= 36'sb1011010010011000110101100101011010;
            sine_reg0   <= 36'sb11101111100010111011100000000010010;
        end
        3157: begin
            cosine_reg0 <= 36'sb1011010001101001110011001001010110;
            sine_reg0   <= 36'sb11101111100101001001010001001101101;
        end
        3158: begin
            cosine_reg0 <= 36'sb1011010000111010110000010001011101;
            sine_reg0   <= 36'sb11101111100111010110111001001010000;
        end
        3159: begin
            cosine_reg0 <= 36'sb1011010000001011101100111101110010;
            sine_reg0   <= 36'sb11101111101001100100010111110111000;
        end
        3160: begin
            cosine_reg0 <= 36'sb1011001111011100101001001110010101;
            sine_reg0   <= 36'sb11101111101011110001101101010100110;
        end
        3161: begin
            cosine_reg0 <= 36'sb1011001110101101100101000011001010;
            sine_reg0   <= 36'sb11101111101101111110111001100011001;
        end
        3162: begin
            cosine_reg0 <= 36'sb1011001101111110100000011100010001;
            sine_reg0   <= 36'sb11101111110000001011111100100010000;
        end
        3163: begin
            cosine_reg0 <= 36'sb1011001101001111011011011001101100;
            sine_reg0   <= 36'sb11101111110010011000110110010001010;
        end
        3164: begin
            cosine_reg0 <= 36'sb1011001100100000010101111011011110;
            sine_reg0   <= 36'sb11101111110100100101100110110000111;
        end
        3165: begin
            cosine_reg0 <= 36'sb1011001011110001010000000001100111;
            sine_reg0   <= 36'sb11101111110110110010001110000000111;
        end
        3166: begin
            cosine_reg0 <= 36'sb1011001011000010001001101100001011;
            sine_reg0   <= 36'sb11101111111000111110101100000000111;
        end
        3167: begin
            cosine_reg0 <= 36'sb1011001010010011000010111011001011;
            sine_reg0   <= 36'sb11101111111011001011000000110001001;
        end
        3168: begin
            cosine_reg0 <= 36'sb1011001001100011111011101110101000;
            sine_reg0   <= 36'sb11101111111101010111001100010001010;
        end
        3169: begin
            cosine_reg0 <= 36'sb1011001000110100110100000110100100;
            sine_reg0   <= 36'sb11101111111111100011001110100001011;
        end
        3170: begin
            cosine_reg0 <= 36'sb1011001000000101101100000011000001;
            sine_reg0   <= 36'sb11110000000001101111000111100001011;
        end
        3171: begin
            cosine_reg0 <= 36'sb1011000111010110100011100100000010;
            sine_reg0   <= 36'sb11110000000011111010110111010001001;
        end
        3172: begin
            cosine_reg0 <= 36'sb1011000110100111011010101001100111;
            sine_reg0   <= 36'sb11110000000110000110011101110000100;
        end
        3173: begin
            cosine_reg0 <= 36'sb1011000101111000010001010011110011;
            sine_reg0   <= 36'sb11110000001000010001111010111111100;
        end
        3174: begin
            cosine_reg0 <= 36'sb1011000101001001000111100010100111;
            sine_reg0   <= 36'sb11110000001010011101001110111110000;
        end
        3175: begin
            cosine_reg0 <= 36'sb1011000100011001111101010110000110;
            sine_reg0   <= 36'sb11110000001100101000011001101011111;
        end
        3176: begin
            cosine_reg0 <= 36'sb1011000011101010110010101110010001;
            sine_reg0   <= 36'sb11110000001110110011011011001001001;
        end
        3177: begin
            cosine_reg0 <= 36'sb1011000010111011100111101011001001;
            sine_reg0   <= 36'sb11110000010000111110010011010101101;
        end
        3178: begin
            cosine_reg0 <= 36'sb1011000010001100011100001100110010;
            sine_reg0   <= 36'sb11110000010011001001000010010001010;
        end
        3179: begin
            cosine_reg0 <= 36'sb1011000001011101010000010011001100;
            sine_reg0   <= 36'sb11110000010101010011100111111100000;
        end
        3180: begin
            cosine_reg0 <= 36'sb1011000000101110000011111110011001;
            sine_reg0   <= 36'sb11110000010111011110000100010101110;
        end
        3181: begin
            cosine_reg0 <= 36'sb1010111111111110110111001110011011;
            sine_reg0   <= 36'sb11110000011001101000010111011110100;
        end
        3182: begin
            cosine_reg0 <= 36'sb1010111111001111101010000011010100;
            sine_reg0   <= 36'sb11110000011011110010100001010110000;
        end
        3183: begin
            cosine_reg0 <= 36'sb1010111110100000011100011101000111;
            sine_reg0   <= 36'sb11110000011101111100100001111100010;
        end
        3184: begin
            cosine_reg0 <= 36'sb1010111101110001001110011011110011;
            sine_reg0   <= 36'sb11110000100000000110011001010001001;
        end
        3185: begin
            cosine_reg0 <= 36'sb1010111101000001111111111111011101;
            sine_reg0   <= 36'sb11110000100010010000000111010100110;
        end
        3186: begin
            cosine_reg0 <= 36'sb1010111100010010110001001000000100;
            sine_reg0   <= 36'sb11110000100100011001101100000110110;
        end
        3187: begin
            cosine_reg0 <= 36'sb1010111011100011100001110101101100;
            sine_reg0   <= 36'sb11110000100110100011000111100111001;
        end
        3188: begin
            cosine_reg0 <= 36'sb1010111010110100010010001000010110;
            sine_reg0   <= 36'sb11110000101000101100011001110101111;
        end
        3189: begin
            cosine_reg0 <= 36'sb1010111010000101000010000000000011;
            sine_reg0   <= 36'sb11110000101010110101100010110011000;
        end
        3190: begin
            cosine_reg0 <= 36'sb1010111001010101110001011100110110;
            sine_reg0   <= 36'sb11110000101100111110100010011110001;
        end
        3191: begin
            cosine_reg0 <= 36'sb1010111000100110100000011110110000;
            sine_reg0   <= 36'sb11110000101111000111011000110111100;
        end
        3192: begin
            cosine_reg0 <= 36'sb1010110111110111001111000101110011;
            sine_reg0   <= 36'sb11110000110001010000000101111110110;
        end
        3193: begin
            cosine_reg0 <= 36'sb1010110111000111111101010010000010;
            sine_reg0   <= 36'sb11110000110011011000101001110100000;
        end
        3194: begin
            cosine_reg0 <= 36'sb1010110110011000101011000011011101;
            sine_reg0   <= 36'sb11110000110101100001000100010111001;
        end
        3195: begin
            cosine_reg0 <= 36'sb1010110101101001011000011010000111;
            sine_reg0   <= 36'sb11110000110111101001010101100111111;
        end
        3196: begin
            cosine_reg0 <= 36'sb1010110100111010000101010110000010;
            sine_reg0   <= 36'sb11110000111001110001011101100110011;
        end
        3197: begin
            cosine_reg0 <= 36'sb1010110100001010110001110111001110;
            sine_reg0   <= 36'sb11110000111011111001011100010010100;
        end
        3198: begin
            cosine_reg0 <= 36'sb1010110011011011011101111101101111;
            sine_reg0   <= 36'sb11110000111110000001010001101100001;
        end
        3199: begin
            cosine_reg0 <= 36'sb1010110010101100001001101001100110;
            sine_reg0   <= 36'sb11110001000000001000111101110011001;
        end
        3200: begin
            cosine_reg0 <= 36'sb1010110001111100110100111010110101;
            sine_reg0   <= 36'sb11110001000010010000100000100111101;
        end
        3201: begin
            cosine_reg0 <= 36'sb1010110001001101011111110001011101;
            sine_reg0   <= 36'sb11110001000100010111111010001001010;
        end
        3202: begin
            cosine_reg0 <= 36'sb1010110000011110001010001101100001;
            sine_reg0   <= 36'sb11110001000110011111001010011000001;
        end
        3203: begin
            cosine_reg0 <= 36'sb1010101111101110110100001111000010;
            sine_reg0   <= 36'sb11110001001000100110010001010100001;
        end
        3204: begin
            cosine_reg0 <= 36'sb1010101110111111011101110110000010;
            sine_reg0   <= 36'sb11110001001010101101001110111101001;
        end
        3205: begin
            cosine_reg0 <= 36'sb1010101110010000000111000010100011;
            sine_reg0   <= 36'sb11110001001100110100000011010011000;
        end
        3206: begin
            cosine_reg0 <= 36'sb1010101101100000101111110100100111;
            sine_reg0   <= 36'sb11110001001110111010101110010101110;
        end
        3207: begin
            cosine_reg0 <= 36'sb1010101100110001011000001100001111;
            sine_reg0   <= 36'sb11110001010001000001010000000101011;
        end
        3208: begin
            cosine_reg0 <= 36'sb1010101100000010000000001001011110;
            sine_reg0   <= 36'sb11110001010011000111101000100001101;
        end
        3209: begin
            cosine_reg0 <= 36'sb1010101011010010100111101100010101;
            sine_reg0   <= 36'sb11110001010101001101110111101010101;
        end
        3210: begin
            cosine_reg0 <= 36'sb1010101010100011001110110100110110;
            sine_reg0   <= 36'sb11110001010111010011111101100000000;
        end
        3211: begin
            cosine_reg0 <= 36'sb1010101001110011110101100011000011;
            sine_reg0   <= 36'sb11110001011001011001111010000001111;
        end
        3212: begin
            cosine_reg0 <= 36'sb1010101001000100011011110110111110;
            sine_reg0   <= 36'sb11110001011011011111101101010000001;
        end
        3213: begin
            cosine_reg0 <= 36'sb1010101000010101000001110000101000;
            sine_reg0   <= 36'sb11110001011101100101010111001010110;
        end
        3214: begin
            cosine_reg0 <= 36'sb1010100111100101100111010000000011;
            sine_reg0   <= 36'sb11110001011111101010110111110001100;
        end
        3215: begin
            cosine_reg0 <= 36'sb1010100110110110001100010101010010;
            sine_reg0   <= 36'sb11110001100001110000001111000100011;
        end
        3216: begin
            cosine_reg0 <= 36'sb1010100110000110110001000000010110;
            sine_reg0   <= 36'sb11110001100011110101011101000011011;
        end
        3217: begin
            cosine_reg0 <= 36'sb1010100101010111010101010001010000;
            sine_reg0   <= 36'sb11110001100101111010100001101110011;
        end
        3218: begin
            cosine_reg0 <= 36'sb1010100100100111111001001000000011;
            sine_reg0   <= 36'sb11110001100111111111011101000101010;
        end
        3219: begin
            cosine_reg0 <= 36'sb1010100011111000011100100100110001;
            sine_reg0   <= 36'sb11110001101010000100001111000111111;
        end
        3220: begin
            cosine_reg0 <= 36'sb1010100011001000111111100111011011;
            sine_reg0   <= 36'sb11110001101100001000110111110110010;
        end
        3221: begin
            cosine_reg0 <= 36'sb1010100010011001100010010000000011;
            sine_reg0   <= 36'sb11110001101110001101010111010000010;
        end
        3222: begin
            cosine_reg0 <= 36'sb1010100001101010000100011110101011;
            sine_reg0   <= 36'sb11110001110000010001101101010101111;
        end
        3223: begin
            cosine_reg0 <= 36'sb1010100000111010100110010011010101;
            sine_reg0   <= 36'sb11110001110010010101111010000111000;
        end
        3224: begin
            cosine_reg0 <= 36'sb1010100000001011000111101110000011;
            sine_reg0   <= 36'sb11110001110100011001111101100011101;
        end
        3225: begin
            cosine_reg0 <= 36'sb1010011111011011101000101110110110;
            sine_reg0   <= 36'sb11110001110110011101110111101011011;
        end
        3226: begin
            cosine_reg0 <= 36'sb1010011110101100001001010101110000;
            sine_reg0   <= 36'sb11110001111000100001101000011110100;
        end
        3227: begin
            cosine_reg0 <= 36'sb1010011101111100101001100010110100;
            sine_reg0   <= 36'sb11110001111010100101001111111100111;
        end
        3228: begin
            cosine_reg0 <= 36'sb1010011101001101001001010110000010;
            sine_reg0   <= 36'sb11110001111100101000101110000110010;
        end
        3229: begin
            cosine_reg0 <= 36'sb1010011100011101101000101111011110;
            sine_reg0   <= 36'sb11110001111110101100000010111010101;
        end
        3230: begin
            cosine_reg0 <= 36'sb1010011011101110000111101111001000;
            sine_reg0   <= 36'sb11110010000000101111001110011010000;
        end
        3231: begin
            cosine_reg0 <= 36'sb1010011010111110100110010101000010;
            sine_reg0   <= 36'sb11110010000010110010010000100100010;
        end
        3232: begin
            cosine_reg0 <= 36'sb1010011010001111000100100001001111;
            sine_reg0   <= 36'sb11110010000100110101001001011001010;
        end
        3233: begin
            cosine_reg0 <= 36'sb1010011001011111100010010011110000;
            sine_reg0   <= 36'sb11110010000110110111111000111001000;
        end
        3234: begin
            cosine_reg0 <= 36'sb1010011000101111111111101100100110;
            sine_reg0   <= 36'sb11110010001000111010011111000011010;
        end
        3235: begin
            cosine_reg0 <= 36'sb1010011000000000011100101011110101;
            sine_reg0   <= 36'sb11110010001010111100111011111000001;
        end
        3236: begin
            cosine_reg0 <= 36'sb1010010111010000111001010001011101;
            sine_reg0   <= 36'sb11110010001100111111001111010111100;
        end
        3237: begin
            cosine_reg0 <= 36'sb1010010110100001010101011101100001;
            sine_reg0   <= 36'sb11110010001111000001011001100001010;
        end
        3238: begin
            cosine_reg0 <= 36'sb1010010101110001110001010000000010;
            sine_reg0   <= 36'sb11110010010001000011011010010101010;
        end
        3239: begin
            cosine_reg0 <= 36'sb1010010101000010001100101001000010;
            sine_reg0   <= 36'sb11110010010011000101010001110011100;
        end
        3240: begin
            cosine_reg0 <= 36'sb1010010100010010100111101000100011;
            sine_reg0   <= 36'sb11110010010101000110111111111100000;
        end
        3241: begin
            cosine_reg0 <= 36'sb1010010011100011000010001110100111;
            sine_reg0   <= 36'sb11110010010111001000100100101110011;
        end
        3242: begin
            cosine_reg0 <= 36'sb1010010010110011011100011011001111;
            sine_reg0   <= 36'sb11110010011001001010000000001010111;
        end
        3243: begin
            cosine_reg0 <= 36'sb1010010010000011110110001110011110;
            sine_reg0   <= 36'sb11110010011011001011010010010001011;
        end
        3244: begin
            cosine_reg0 <= 36'sb1010010001010100001111101000010110;
            sine_reg0   <= 36'sb11110010011101001100011011000001101;
        end
        3245: begin
            cosine_reg0 <= 36'sb1010010000100100101000101000110111;
            sine_reg0   <= 36'sb11110010011111001101011010011011101;
        end
        3246: begin
            cosine_reg0 <= 36'sb1010001111110101000001010000000101;
            sine_reg0   <= 36'sb11110010100001001110010000011111010;
        end
        3247: begin
            cosine_reg0 <= 36'sb1010001111000101011001011110000000;
            sine_reg0   <= 36'sb11110010100011001110111101001100101;
        end
        3248: begin
            cosine_reg0 <= 36'sb1010001110010101110001010010101011;
            sine_reg0   <= 36'sb11110010100101001111100000100011100;
        end
        3249: begin
            cosine_reg0 <= 36'sb1010001101100110001000101110000111;
            sine_reg0   <= 36'sb11110010100111001111111010100011110;
        end
        3250: begin
            cosine_reg0 <= 36'sb1010001100110110011111110000010111;
            sine_reg0   <= 36'sb11110010101001010000001011001101011;
        end
        3251: begin
            cosine_reg0 <= 36'sb1010001100000110110110011001011011;
            sine_reg0   <= 36'sb11110010101011010000010010100000011;
        end
        3252: begin
            cosine_reg0 <= 36'sb1010001011010111001100101001010111;
            sine_reg0   <= 36'sb11110010101101010000010000011100101;
        end
        3253: begin
            cosine_reg0 <= 36'sb1010001010100111100010100000001100;
            sine_reg0   <= 36'sb11110010101111010000000101000001111;
        end
        3254: begin
            cosine_reg0 <= 36'sb1010001001110111110111111101111011;
            sine_reg0   <= 36'sb11110010110001001111110000010000011;
        end
        3255: begin
            cosine_reg0 <= 36'sb1010001001001000001101000010100111;
            sine_reg0   <= 36'sb11110010110011001111010010000111110;
        end
        3256: begin
            cosine_reg0 <= 36'sb1010001000011000100001101110010001;
            sine_reg0   <= 36'sb11110010110101001110101010101000000;
        end
        3257: begin
            cosine_reg0 <= 36'sb1010000111101000110110000000111011;
            sine_reg0   <= 36'sb11110010110111001101111001110001001;
        end
        3258: begin
            cosine_reg0 <= 36'sb1010000110111001001001111010100111;
            sine_reg0   <= 36'sb11110010111001001100111111100011001;
        end
        3259: begin
            cosine_reg0 <= 36'sb1010000110001001011101011011011000;
            sine_reg0   <= 36'sb11110010111011001011111011111101101;
        end
        3260: begin
            cosine_reg0 <= 36'sb1010000101011001110000100011001101;
            sine_reg0   <= 36'sb11110010111101001010101111000000111;
        end
        3261: begin
            cosine_reg0 <= 36'sb1010000100101010000011010010001011;
            sine_reg0   <= 36'sb11110010111111001001011000101100101;
        end
        3262: begin
            cosine_reg0 <= 36'sb1010000011111010010101101000010010;
            sine_reg0   <= 36'sb11110011000001000111111001000000110;
        end
        3263: begin
            cosine_reg0 <= 36'sb1010000011001010100111100101100100;
            sine_reg0   <= 36'sb11110011000011000110001111111101010;
        end
        3264: begin
            cosine_reg0 <= 36'sb1010000010011010111001001010000011;
            sine_reg0   <= 36'sb11110011000101000100011101100010001;
        end
        3265: begin
            cosine_reg0 <= 36'sb1010000001101011001010010101110001;
            sine_reg0   <= 36'sb11110011000111000010100001101111010;
        end
        3266: begin
            cosine_reg0 <= 36'sb1010000000111011011011001000101111;
            sine_reg0   <= 36'sb11110011001001000000011100100100100;
        end
        3267: begin
            cosine_reg0 <= 36'sb1010000000001011101011100011000000;
            sine_reg0   <= 36'sb11110011001010111110001110000001110;
        end
        3268: begin
            cosine_reg0 <= 36'sb1001111111011011111011100100100110;
            sine_reg0   <= 36'sb11110011001100111011110110000111001;
        end
        3269: begin
            cosine_reg0 <= 36'sb1001111110101100001011001101100010;
            sine_reg0   <= 36'sb11110011001110111001010100110100011;
        end
        3270: begin
            cosine_reg0 <= 36'sb1001111101111100011010011101110110;
            sine_reg0   <= 36'sb11110011010000110110101010001001011;
        end
        3271: begin
            cosine_reg0 <= 36'sb1001111101001100101001010101100100;
            sine_reg0   <= 36'sb11110011010010110011110110000110010;
        end
        3272: begin
            cosine_reg0 <= 36'sb1001111100011100110111110100101110;
            sine_reg0   <= 36'sb11110011010100110000111000101010110;
        end
        3273: begin
            cosine_reg0 <= 36'sb1001111011101101000101111011010101;
            sine_reg0   <= 36'sb11110011010110101101110001110111000;
        end
        3274: begin
            cosine_reg0 <= 36'sb1001111010111101010011101001011100;
            sine_reg0   <= 36'sb11110011011000101010100001101010101;
        end
        3275: begin
            cosine_reg0 <= 36'sb1001111010001101100000111111000100;
            sine_reg0   <= 36'sb11110011011010100111001000000101111;
        end
        3276: begin
            cosine_reg0 <= 36'sb1001111001011101101101111100001111;
            sine_reg0   <= 36'sb11110011011100100011100101001000100;
        end
        3277: begin
            cosine_reg0 <= 36'sb1001111000101101111010100000111111;
            sine_reg0   <= 36'sb11110011011110011111111000110010011;
        end
        3278: begin
            cosine_reg0 <= 36'sb1001110111111110000110101101010110;
            sine_reg0   <= 36'sb11110011100000011100000011000011100;
        end
        3279: begin
            cosine_reg0 <= 36'sb1001110111001110010010100001010110;
            sine_reg0   <= 36'sb11110011100010011000000011111011110;
        end
        3280: begin
            cosine_reg0 <= 36'sb1001110110011110011101111101000000;
            sine_reg0   <= 36'sb11110011100100010011111011011011010;
        end
        3281: begin
            cosine_reg0 <= 36'sb1001110101101110101001000000010111;
            sine_reg0   <= 36'sb11110011100110001111101001100001101;
        end
        3282: begin
            cosine_reg0 <= 36'sb1001110100111110110011101011011100;
            sine_reg0   <= 36'sb11110011101000001011001110001111000;
        end
        3283: begin
            cosine_reg0 <= 36'sb1001110100001110111101111110010000;
            sine_reg0   <= 36'sb11110011101010000110101001100011010;
        end
        3284: begin
            cosine_reg0 <= 36'sb1001110011011111000111111000110111;
            sine_reg0   <= 36'sb11110011101100000001111011011110011;
        end
        3285: begin
            cosine_reg0 <= 36'sb1001110010101111010001011011010010;
            sine_reg0   <= 36'sb11110011101101111101000100000000001;
        end
        3286: begin
            cosine_reg0 <= 36'sb1001110001111111011010100101100010;
            sine_reg0   <= 36'sb11110011101111111000000011001000100;
        end
        3287: begin
            cosine_reg0 <= 36'sb1001110001001111100011010111101001;
            sine_reg0   <= 36'sb11110011110001110010111000110111100;
        end
        3288: begin
            cosine_reg0 <= 36'sb1001110000011111101011110001101010;
            sine_reg0   <= 36'sb11110011110011101101100101001101000;
        end
        3289: begin
            cosine_reg0 <= 36'sb1001101111101111110011110011100110;
            sine_reg0   <= 36'sb11110011110101101000001000001001000;
        end
        3290: begin
            cosine_reg0 <= 36'sb1001101110111111111011011101011111;
            sine_reg0   <= 36'sb11110011110111100010100001101011010;
        end
        3291: begin
            cosine_reg0 <= 36'sb1001101110010000000010101111010111;
            sine_reg0   <= 36'sb11110011111001011100110001110011111;
        end
        3292: begin
            cosine_reg0 <= 36'sb1001101101100000001001101001001111;
            sine_reg0   <= 36'sb11110011111011010110111000100010101;
        end
        3293: begin
            cosine_reg0 <= 36'sb1001101100110000010000001011001010;
            sine_reg0   <= 36'sb11110011111101010000110101110111100;
        end
        3294: begin
            cosine_reg0 <= 36'sb1001101100000000010110010101001001;
            sine_reg0   <= 36'sb11110011111111001010101001110010100;
        end
        3295: begin
            cosine_reg0 <= 36'sb1001101011010000011100000111001110;
            sine_reg0   <= 36'sb11110100000001000100010100010011011;
        end
        3296: begin
            cosine_reg0 <= 36'sb1001101010100000100001100001011100;
            sine_reg0   <= 36'sb11110100000010111101110101011010010;
        end
        3297: begin
            cosine_reg0 <= 36'sb1001101001110000100110100011110011;
            sine_reg0   <= 36'sb11110100000100110111001101000111000;
        end
        3298: begin
            cosine_reg0 <= 36'sb1001101001000000101011001110010110;
            sine_reg0   <= 36'sb11110100000110110000011011011001100;
        end
        3299: begin
            cosine_reg0 <= 36'sb1001101000010000101111100001000111;
            sine_reg0   <= 36'sb11110100001000101001100000010001101;
        end
        3300: begin
            cosine_reg0 <= 36'sb1001100111100000110011011100000111;
            sine_reg0   <= 36'sb11110100001010100010011011101111011;
        end
        3301: begin
            cosine_reg0 <= 36'sb1001100110110000110110111111011000;
            sine_reg0   <= 36'sb11110100001100011011001101110010110;
        end
        3302: begin
            cosine_reg0 <= 36'sb1001100110000000111010001010111101;
            sine_reg0   <= 36'sb11110100001110010011110110011011100;
        end
        3303: begin
            cosine_reg0 <= 36'sb1001100101010000111100111110110110;
            sine_reg0   <= 36'sb11110100010000001100010101101001110;
        end
        3304: begin
            cosine_reg0 <= 36'sb1001100100100000111111011011000111;
            sine_reg0   <= 36'sb11110100010010000100101011011101010;
        end
        3305: begin
            cosine_reg0 <= 36'sb1001100011110001000001011111110000;
            sine_reg0   <= 36'sb11110100010011111100110111110110001;
        end
        3306: begin
            cosine_reg0 <= 36'sb1001100011000001000011001100110011;
            sine_reg0   <= 36'sb11110100010101110100111010110100001;
        end
        3307: begin
            cosine_reg0 <= 36'sb1001100010010001000100100010010011;
            sine_reg0   <= 36'sb11110100010111101100110100010111001;
        end
        3308: begin
            cosine_reg0 <= 36'sb1001100001100001000101100000010001;
            sine_reg0   <= 36'sb11110100011001100100100100011111010;
        end
        3309: begin
            cosine_reg0 <= 36'sb1001100000110001000110000110110000;
            sine_reg0   <= 36'sb11110100011011011100001011001100011;
        end
        3310: begin
            cosine_reg0 <= 36'sb1001100000000001000110010101110000;
            sine_reg0   <= 36'sb11110100011101010011101000011110011;
        end
        3311: begin
            cosine_reg0 <= 36'sb1001011111010001000110001101010100;
            sine_reg0   <= 36'sb11110100011111001010111100010101010;
        end
        3312: begin
            cosine_reg0 <= 36'sb1001011110100001000101101101011101;
            sine_reg0   <= 36'sb11110100100001000010000110110000111;
        end
        3313: begin
            cosine_reg0 <= 36'sb1001011101110001000100110110001110;
            sine_reg0   <= 36'sb11110100100010111001000111110001001;
        end
        3314: begin
            cosine_reg0 <= 36'sb1001011101000001000011100111101001;
            sine_reg0   <= 36'sb11110100100100101111111111010110000;
        end
        3315: begin
            cosine_reg0 <= 36'sb1001011100010001000010000001101110;
            sine_reg0   <= 36'sb11110100100110100110101101011111011;
        end
        3316: begin
            cosine_reg0 <= 36'sb1001011011100001000000000100100001;
            sine_reg0   <= 36'sb11110100101000011101010010001101010;
        end
        3317: begin
            cosine_reg0 <= 36'sb1001011010110000111101110000000010;
            sine_reg0   <= 36'sb11110100101010010011101101011111100;
        end
        3318: begin
            cosine_reg0 <= 36'sb1001011010000000111011000100010100;
            sine_reg0   <= 36'sb11110100101100001001111111010110001;
        end
        3319: begin
            cosine_reg0 <= 36'sb1001011001010000111000000001011001;
            sine_reg0   <= 36'sb11110100101110000000000111110000111;
        end
        3320: begin
            cosine_reg0 <= 36'sb1001011000100000110100100111010010;
            sine_reg0   <= 36'sb11110100101111110110000110101111111;
        end
        3321: begin
            cosine_reg0 <= 36'sb1001010111110000110000110110000010;
            sine_reg0   <= 36'sb11110100110001101011111100010011000;
        end
        3322: begin
            cosine_reg0 <= 36'sb1001010111000000101100101101101010;
            sine_reg0   <= 36'sb11110100110011100001101000011010010;
        end
        3323: begin
            cosine_reg0 <= 36'sb1001010110010000101000001110001011;
            sine_reg0   <= 36'sb11110100110101010111001011000101011;
        end
        3324: begin
            cosine_reg0 <= 36'sb1001010101100000100011010111101001;
            sine_reg0   <= 36'sb11110100110111001100100100010100011;
        end
        3325: begin
            cosine_reg0 <= 36'sb1001010100110000011110001010000100;
            sine_reg0   <= 36'sb11110100111001000001110100000111010;
        end
        3326: begin
            cosine_reg0 <= 36'sb1001010100000000011000100101011111;
            sine_reg0   <= 36'sb11110100111010110110111010011101111;
        end
        3327: begin
            cosine_reg0 <= 36'sb1001010011010000010010101001111011;
            sine_reg0   <= 36'sb11110100111100101011110111011000001;
        end
        3328: begin
            cosine_reg0 <= 36'sb1001010010100000001100010111011010;
            sine_reg0   <= 36'sb11110100111110100000101010110110001;
        end
        3329: begin
            cosine_reg0 <= 36'sb1001010001110000000101101101111111;
            sine_reg0   <= 36'sb11110101000000010101010100110111100;
        end
        3330: begin
            cosine_reg0 <= 36'sb1001010000111111111110101101101011;
            sine_reg0   <= 36'sb11110101000010001001110101011100100;
        end
        3331: begin
            cosine_reg0 <= 36'sb1001010000001111110111010110011111;
            sine_reg0   <= 36'sb11110101000011111110001100100100110;
        end
        3332: begin
            cosine_reg0 <= 36'sb1001001111011111101111101000011110;
            sine_reg0   <= 36'sb11110101000101110010011010010000100;
        end
        3333: begin
            cosine_reg0 <= 36'sb1001001110101111100111100011101010;
            sine_reg0   <= 36'sb11110101000111100110011110011111011;
        end
        3334: begin
            cosine_reg0 <= 36'sb1001001101111111011111001000000100;
            sine_reg0   <= 36'sb11110101001001011010011001010001100;
        end
        3335: begin
            cosine_reg0 <= 36'sb1001001101001111010110010101101110;
            sine_reg0   <= 36'sb11110101001011001110001010100110110;
        end
        3336: begin
            cosine_reg0 <= 36'sb1001001100011111001101001100101010;
            sine_reg0   <= 36'sb11110101001101000001110010011111001;
        end
        3337: begin
            cosine_reg0 <= 36'sb1001001011101111000011101100111011;
            sine_reg0   <= 36'sb11110101001110110101010000111010011;
        end
        3338: begin
            cosine_reg0 <= 36'sb1001001010111110111001110110100001;
            sine_reg0   <= 36'sb11110101010000101000100101111000101;
        end
        3339: begin
            cosine_reg0 <= 36'sb1001001010001110101111101001011111;
            sine_reg0   <= 36'sb11110101010010011011110001011001101;
        end
        3340: begin
            cosine_reg0 <= 36'sb1001001001011110100101000101110110;
            sine_reg0   <= 36'sb11110101010100001110110011011101100;
        end
        3341: begin
            cosine_reg0 <= 36'sb1001001000101110011010001011101001;
            sine_reg0   <= 36'sb11110101010110000001101100000100000;
        end
        3342: begin
            cosine_reg0 <= 36'sb1001000111111110001110111010111001;
            sine_reg0   <= 36'sb11110101010111110100011011001101001;
        end
        3343: begin
            cosine_reg0 <= 36'sb1001000111001110000011010011101000;
            sine_reg0   <= 36'sb11110101011001100111000000111000111;
        end
        3344: begin
            cosine_reg0 <= 36'sb1001000110011101110111010101111000;
            sine_reg0   <= 36'sb11110101011011011001011101000111001;
        end
        3345: begin
            cosine_reg0 <= 36'sb1001000101101101101011000001101011;
            sine_reg0   <= 36'sb11110101011101001011101111110111110;
        end
        3346: begin
            cosine_reg0 <= 36'sb1001000100111101011110010111000011;
            sine_reg0   <= 36'sb11110101011110111101111001001010111;
        end
        3347: begin
            cosine_reg0 <= 36'sb1001000100001101010001010110000001;
            sine_reg0   <= 36'sb11110101100000101111111001000000001;
        end
        3348: begin
            cosine_reg0 <= 36'sb1001000011011101000011111110100111;
            sine_reg0   <= 36'sb11110101100010100001101111010111101;
        end
        3349: begin
            cosine_reg0 <= 36'sb1001000010101100110110010000111000;
            sine_reg0   <= 36'sb11110101100100010011011100010001011;
        end
        3350: begin
            cosine_reg0 <= 36'sb1001000001111100101000001100110101;
            sine_reg0   <= 36'sb11110101100110000100111111101101001;
        end
        3351: begin
            cosine_reg0 <= 36'sb1001000001001100011001110010100000;
            sine_reg0   <= 36'sb11110101100111110110011001101011000;
        end
        3352: begin
            cosine_reg0 <= 36'sb1001000000011100001011000001111011;
            sine_reg0   <= 36'sb11110101101001100111101010001010110;
        end
        3353: begin
            cosine_reg0 <= 36'sb1000111111101011111011111011000111;
            sine_reg0   <= 36'sb11110101101011011000110001001100011;
        end
        3354: begin
            cosine_reg0 <= 36'sb1000111110111011101100011110000111;
            sine_reg0   <= 36'sb11110101101101001001101110101111111;
        end
        3355: begin
            cosine_reg0 <= 36'sb1000111110001011011100101010111100;
            sine_reg0   <= 36'sb11110101101110111010100010110101000;
        end
        3356: begin
            cosine_reg0 <= 36'sb1000111101011011001100100001101001;
            sine_reg0   <= 36'sb11110101110000101011001101011011111;
        end
        3357: begin
            cosine_reg0 <= 36'sb1000111100101010111100000010001111;
            sine_reg0   <= 36'sb11110101110010011011101110100100011;
        end
        3358: begin
            cosine_reg0 <= 36'sb1000111011111010101011001100101111;
            sine_reg0   <= 36'sb11110101110100001100000110001110011;
        end
        3359: begin
            cosine_reg0 <= 36'sb1000111011001010011010000001001101;
            sine_reg0   <= 36'sb11110101110101111100010100011010000;
        end
        3360: begin
            cosine_reg0 <= 36'sb1000111010011010001000011111101001;
            sine_reg0   <= 36'sb11110101110111101100011001000110111;
        end
        3361: begin
            cosine_reg0 <= 36'sb1000111001101001110110101000000110;
            sine_reg0   <= 36'sb11110101111001011100010100010101001;
        end
        3362: begin
            cosine_reg0 <= 36'sb1000111000111001100100011010100110;
            sine_reg0   <= 36'sb11110101111011001100000110000100101;
        end
        3363: begin
            cosine_reg0 <= 36'sb1000111000001001010001110111001001;
            sine_reg0   <= 36'sb11110101111100111011101110010101011;
        end
        3364: begin
            cosine_reg0 <= 36'sb1000110111011000111110111101110011;
            sine_reg0   <= 36'sb11110101111110101011001101000111010;
        end
        3365: begin
            cosine_reg0 <= 36'sb1000110110101000101011101110100101;
            sine_reg0   <= 36'sb11110110000000011010100010011010001;
        end
        3366: begin
            cosine_reg0 <= 36'sb1000110101111000011000001001100000;
            sine_reg0   <= 36'sb11110110000010001001101110001110001;
        end
        3367: begin
            cosine_reg0 <= 36'sb1000110101001000000100001110101000;
            sine_reg0   <= 36'sb11110110000011111000110000100011000;
        end
        3368: begin
            cosine_reg0 <= 36'sb1000110100010111101111111101111101;
            sine_reg0   <= 36'sb11110110000101100111101001011000110;
        end
        3369: begin
            cosine_reg0 <= 36'sb1000110011100111011011010111100001;
            sine_reg0   <= 36'sb11110110000111010110011000101111010;
        end
        3370: begin
            cosine_reg0 <= 36'sb1000110010110111000110011011010111;
            sine_reg0   <= 36'sb11110110001001000100111110100110100;
        end
        3371: begin
            cosine_reg0 <= 36'sb1000110010000110110001001001100000;
            sine_reg0   <= 36'sb11110110001010110011011010111110100;
        end
        3372: begin
            cosine_reg0 <= 36'sb1000110001010110011011100001111110;
            sine_reg0   <= 36'sb11110110001100100001101101110111001;
        end
        3373: begin
            cosine_reg0 <= 36'sb1000110000100110000101100100110011;
            sine_reg0   <= 36'sb11110110001110001111110111010000001;
        end
        3374: begin
            cosine_reg0 <= 36'sb1000101111110101101111010010000001;
            sine_reg0   <= 36'sb11110110001111111101110111001001110;
        end
        3375: begin
            cosine_reg0 <= 36'sb1000101111000101011000101001101010;
            sine_reg0   <= 36'sb11110110010001101011101101100011110;
        end
        3376: begin
            cosine_reg0 <= 36'sb1000101110010101000001101011101111;
            sine_reg0   <= 36'sb11110110010011011001011010011110000;
        end
        3377: begin
            cosine_reg0 <= 36'sb1000101101100100101010011000010010;
            sine_reg0   <= 36'sb11110110010101000110111101111000101;
        end
        3378: begin
            cosine_reg0 <= 36'sb1000101100110100010010101111010101;
            sine_reg0   <= 36'sb11110110010110110100010111110011011;
        end
        3379: begin
            cosine_reg0 <= 36'sb1000101100000011111010110000111011;
            sine_reg0   <= 36'sb11110110011000100001101000001110010;
        end
        3380: begin
            cosine_reg0 <= 36'sb1000101011010011100010011101000101;
            sine_reg0   <= 36'sb11110110011010001110101111001001010;
        end
        3381: begin
            cosine_reg0 <= 36'sb1000101010100011001001110011110100;
            sine_reg0   <= 36'sb11110110011011111011101100100100010;
        end
        3382: begin
            cosine_reg0 <= 36'sb1000101001110010110000110101001100;
            sine_reg0   <= 36'sb11110110011101101000100000011111010;
        end
        3383: begin
            cosine_reg0 <= 36'sb1000101001000010010111100001001100;
            sine_reg0   <= 36'sb11110110011111010101001010111010000;
        end
        3384: begin
            cosine_reg0 <= 36'sb1000101000010001111101110111111001;
            sine_reg0   <= 36'sb11110110100001000001101011110100101;
        end
        3385: begin
            cosine_reg0 <= 36'sb1000100111100001100011111001010010;
            sine_reg0   <= 36'sb11110110100010101110000011001111000;
        end
        3386: begin
            cosine_reg0 <= 36'sb1000100110110001001001100101011011;
            sine_reg0   <= 36'sb11110110100100011010010001001001001;
        end
        3387: begin
            cosine_reg0 <= 36'sb1000100110000000101110111100010100;
            sine_reg0   <= 36'sb11110110100110000110010101100010110;
        end
        3388: begin
            cosine_reg0 <= 36'sb1000100101010000010011111110000001;
            sine_reg0   <= 36'sb11110110100111110010010000011100000;
        end
        3389: begin
            cosine_reg0 <= 36'sb1000100100011111111000101010100011;
            sine_reg0   <= 36'sb11110110101001011110000001110100110;
        end
        3390: begin
            cosine_reg0 <= 36'sb1000100011101111011101000001111011;
            sine_reg0   <= 36'sb11110110101011001001101001101100111;
        end
        3391: begin
            cosine_reg0 <= 36'sb1000100010111111000001000100001011;
            sine_reg0   <= 36'sb11110110101100110101001000000100011;
        end
        3392: begin
            cosine_reg0 <= 36'sb1000100010001110100100110001010110;
            sine_reg0   <= 36'sb11110110101110100000011100111011001;
        end
        3393: begin
            cosine_reg0 <= 36'sb1000100001011110001000001001011101;
            sine_reg0   <= 36'sb11110110110000001011101000010001001;
        end
        3394: begin
            cosine_reg0 <= 36'sb1000100000101101101011001100100010;
            sine_reg0   <= 36'sb11110110110001110110101010000110011;
        end
        3395: begin
            cosine_reg0 <= 36'sb1000011111111101001101111010101000;
            sine_reg0   <= 36'sb11110110110011100001100010011010101;
        end
        3396: begin
            cosine_reg0 <= 36'sb1000011111001100110000010011101111;
            sine_reg0   <= 36'sb11110110110101001100010001001101111;
        end
        3397: begin
            cosine_reg0 <= 36'sb1000011110011100010010010111111001;
            sine_reg0   <= 36'sb11110110110110110110110110100000001;
        end
        3398: begin
            cosine_reg0 <= 36'sb1000011101101011110100000111001010;
            sine_reg0   <= 36'sb11110110111000100001010010010001011;
        end
        3399: begin
            cosine_reg0 <= 36'sb1000011100111011010101100001100010;
            sine_reg0   <= 36'sb11110110111010001011100100100001011;
        end
        3400: begin
            cosine_reg0 <= 36'sb1000011100001010110110100111000011;
            sine_reg0   <= 36'sb11110110111011110101101101010000001;
        end
        3401: begin
            cosine_reg0 <= 36'sb1000011011011010010111010111101111;
            sine_reg0   <= 36'sb11110110111101011111101100011101101;
        end
        3402: begin
            cosine_reg0 <= 36'sb1000011010101001110111110011101000;
            sine_reg0   <= 36'sb11110110111111001001100010001001110;
        end
        3403: begin
            cosine_reg0 <= 36'sb1000011001111001010111111010110001;
            sine_reg0   <= 36'sb11110111000000110011001110010100100;
        end
        3404: begin
            cosine_reg0 <= 36'sb1000011001001000110111101101001010;
            sine_reg0   <= 36'sb11110111000010011100110000111101110;
        end
        3405: begin
            cosine_reg0 <= 36'sb1000011000011000010111001010110101;
            sine_reg0   <= 36'sb11110111000100000110001010000101100;
        end
        3406: begin
            cosine_reg0 <= 36'sb1000010111100111110110010011110110;
            sine_reg0   <= 36'sb11110111000101101111011001101011101;
        end
        3407: begin
            cosine_reg0 <= 36'sb1000010110110111010101001000001100;
            sine_reg0   <= 36'sb11110111000111011000011111110000000;
        end
        3408: begin
            cosine_reg0 <= 36'sb1000010110000110110011100111111011;
            sine_reg0   <= 36'sb11110111001001000001011100010010110;
        end
        3409: begin
            cosine_reg0 <= 36'sb1000010101010110010001110011000100;
            sine_reg0   <= 36'sb11110111001010101010001111010011101;
        end
        3410: begin
            cosine_reg0 <= 36'sb1000010100100101101111101001101001;
            sine_reg0   <= 36'sb11110111001100010010111000110010101;
        end
        3411: begin
            cosine_reg0 <= 36'sb1000010011110101001101001011101100;
            sine_reg0   <= 36'sb11110111001101111011011000101111110;
        end
        3412: begin
            cosine_reg0 <= 36'sb1000010011000100101010011001001111;
            sine_reg0   <= 36'sb11110111001111100011101111001010111;
        end
        3413: begin
            cosine_reg0 <= 36'sb1000010010010100000111010010010100;
            sine_reg0   <= 36'sb11110111010001001011111100000100000;
        end
        3414: begin
            cosine_reg0 <= 36'sb1000010001100011100011110110111011;
            sine_reg0   <= 36'sb11110111010010110011111111011011000;
        end
        3415: begin
            cosine_reg0 <= 36'sb1000010000110011000000000111001001;
            sine_reg0   <= 36'sb11110111010100011011111001001111111;
        end
        3416: begin
            cosine_reg0 <= 36'sb1000010000000010011100000010111101;
            sine_reg0   <= 36'sb11110111010110000011101001100010011;
        end
        3417: begin
            cosine_reg0 <= 36'sb1000001111010001110111101010011011;
            sine_reg0   <= 36'sb11110111010111101011010000010010101;
        end
        3418: begin
            cosine_reg0 <= 36'sb1000001110100001010010111101100011;
            sine_reg0   <= 36'sb11110111011001010010101101100000101;
        end
        3419: begin
            cosine_reg0 <= 36'sb1000001101110000101101111100011001;
            sine_reg0   <= 36'sb11110111011010111010000001001100001;
        end
        3420: begin
            cosine_reg0 <= 36'sb1000001101000000001000100110111101;
            sine_reg0   <= 36'sb11110111011100100001001011010101001;
        end
        3421: begin
            cosine_reg0 <= 36'sb1000001100001111100010111101010010;
            sine_reg0   <= 36'sb11110111011110001000001011111011100;
        end
        3422: begin
            cosine_reg0 <= 36'sb1000001011011110111100111111011001;
            sine_reg0   <= 36'sb11110111011111101111000010111111011;
        end
        3423: begin
            cosine_reg0 <= 36'sb1000001010101110010110101101010101;
            sine_reg0   <= 36'sb11110111100001010101110000100000101;
        end
        3424: begin
            cosine_reg0 <= 36'sb1000001001111101110000000111000111;
            sine_reg0   <= 36'sb11110111100010111100010100011111000;
        end
        3425: begin
            cosine_reg0 <= 36'sb1000001001001101001001001100110001;
            sine_reg0   <= 36'sb11110111100100100010101110111010101;
        end
        3426: begin
            cosine_reg0 <= 36'sb1000001000011100100001111110010101;
            sine_reg0   <= 36'sb11110111100110001000111111110011100;
        end
        3427: begin
            cosine_reg0 <= 36'sb1000000111101011111010011011110101;
            sine_reg0   <= 36'sb11110111100111101111000111001001011;
        end
        3428: begin
            cosine_reg0 <= 36'sb1000000110111011010010100101010010;
            sine_reg0   <= 36'sb11110111101001010101000100111100010;
        end
        3429: begin
            cosine_reg0 <= 36'sb1000000110001010101010011010101111;
            sine_reg0   <= 36'sb11110111101010111010111001001100001;
        end
        3430: begin
            cosine_reg0 <= 36'sb1000000101011010000001111100001110;
            sine_reg0   <= 36'sb11110111101100100000100011111000111;
        end
        3431: begin
            cosine_reg0 <= 36'sb1000000100101001011001001001110000;
            sine_reg0   <= 36'sb11110111101110000110000101000010011;
        end
        3432: begin
            cosine_reg0 <= 36'sb1000000011111000110000000011010111;
            sine_reg0   <= 36'sb11110111101111101011011100101000110;
        end
        3433: begin
            cosine_reg0 <= 36'sb1000000011001000000110101001000101;
            sine_reg0   <= 36'sb11110111110001010000101010101011111;
        end
        3434: begin
            cosine_reg0 <= 36'sb1000000010010111011100111010111101;
            sine_reg0   <= 36'sb11110111110010110101101111001011101;
        end
        3435: begin
            cosine_reg0 <= 36'sb1000000001100110110010111000111111;
            sine_reg0   <= 36'sb11110111110100011010101010000111111;
        end
        3436: begin
            cosine_reg0 <= 36'sb1000000000110110001000100011001110;
            sine_reg0   <= 36'sb11110111110101111111011011100000110;
        end
        3437: begin
            cosine_reg0 <= 36'sb1000000000000101011101111001101011;
            sine_reg0   <= 36'sb11110111110111100100000011010110001;
        end
        3438: begin
            cosine_reg0 <= 36'sb111111111010100110010111100011001;
            sine_reg0   <= 36'sb11110111111001001000100001100111110;
        end
        3439: begin
            cosine_reg0 <= 36'sb111111110100100000111101011011001;
            sine_reg0   <= 36'sb11110111111010101100110110010101111;
        end
        3440: begin
            cosine_reg0 <= 36'sb111111101110011011100000110101110;
            sine_reg0   <= 36'sb11110111111100010001000001100000010;
        end
        3441: begin
            cosine_reg0 <= 36'sb111111101000010110000001110011000;
            sine_reg0   <= 36'sb11110111111101110101000011000110111;
        end
        3442: begin
            cosine_reg0 <= 36'sb111111100010010000100000010011011;
            sine_reg0   <= 36'sb11110111111111011000111011001001101;
        end
        3443: begin
            cosine_reg0 <= 36'sb111111011100001010111100010110111;
            sine_reg0   <= 36'sb11111000000000111100101001101000100;
        end
        3444: begin
            cosine_reg0 <= 36'sb111111010110000101010101111110000;
            sine_reg0   <= 36'sb11111000000010100000001110100011011;
        end
        3445: begin
            cosine_reg0 <= 36'sb111111001111111111101101001000110;
            sine_reg0   <= 36'sb11111000000100000011101001111010010;
        end
        3446: begin
            cosine_reg0 <= 36'sb111111001001111010000001110111011;
            sine_reg0   <= 36'sb11111000000101100110111011101101001;
        end
        3447: begin
            cosine_reg0 <= 36'sb111111000011110100010100001010010;
            sine_reg0   <= 36'sb11111000000111001010000011111011111;
        end
        3448: begin
            cosine_reg0 <= 36'sb111110111101101110100100000001100;
            sine_reg0   <= 36'sb11111000001000101101000010100110011;
        end
        3449: begin
            cosine_reg0 <= 36'sb111110110111101000110001011101011;
            sine_reg0   <= 36'sb11111000001010001111110111101100101;
        end
        3450: begin
            cosine_reg0 <= 36'sb111110110001100010111100011110001;
            sine_reg0   <= 36'sb11111000001011110010100011001110101;
        end
        3451: begin
            cosine_reg0 <= 36'sb111110101011011101000101000100000;
            sine_reg0   <= 36'sb11111000001101010101000101001100001;
        end
        3452: begin
            cosine_reg0 <= 36'sb111110100101010111001011001111010;
            sine_reg0   <= 36'sb11111000001110110111011101100101011;
        end
        3453: begin
            cosine_reg0 <= 36'sb111110011111010001001111000000000;
            sine_reg0   <= 36'sb11111000010000011001101100011010000;
        end
        3454: begin
            cosine_reg0 <= 36'sb111110011001001011010000010110101;
            sine_reg0   <= 36'sb11111000010001111011110001101010001;
        end
        3455: begin
            cosine_reg0 <= 36'sb111110010011000101001111010011010;
            sine_reg0   <= 36'sb11111000010011011101101101010101101;
        end
        3456: begin
            cosine_reg0 <= 36'sb111110001100111111001011110110010;
            sine_reg0   <= 36'sb11111000010100111111011111011100100;
        end
        3457: begin
            cosine_reg0 <= 36'sb111110000110111001000101111111110;
            sine_reg0   <= 36'sb11111000010110100001000111111110101;
        end
        3458: begin
            cosine_reg0 <= 36'sb111110000000110010111101101111111;
            sine_reg0   <= 36'sb11111000011000000010100110111011111;
        end
        3459: begin
            cosine_reg0 <= 36'sb111101111010101100110011000111001;
            sine_reg0   <= 36'sb11111000011001100011111100010100011;
        end
        3460: begin
            cosine_reg0 <= 36'sb111101110100100110100110000101101;
            sine_reg0   <= 36'sb11111000011011000101001000001000000;
        end
        3461: begin
            cosine_reg0 <= 36'sb111101101110100000010110101011100;
            sine_reg0   <= 36'sb11111000011100100110001010010110101;
        end
        3462: begin
            cosine_reg0 <= 36'sb111101101000011010000100111001001;
            sine_reg0   <= 36'sb11111000011110000111000011000000010;
        end
        3463: begin
            cosine_reg0 <= 36'sb111101100010010011110000101110101;
            sine_reg0   <= 36'sb11111000011111100111110010000100110;
        end
        3464: begin
            cosine_reg0 <= 36'sb111101011100001101011010001100011;
            sine_reg0   <= 36'sb11111000100001001000010111100100001;
        end
        3465: begin
            cosine_reg0 <= 36'sb111101010110000111000001010010011;
            sine_reg0   <= 36'sb11111000100010101000110011011110011;
        end
        3466: begin
            cosine_reg0 <= 36'sb111101010000000000100110000001001;
            sine_reg0   <= 36'sb11111000100100001001000101110011011;
        end
        3467: begin
            cosine_reg0 <= 36'sb111101001001111010001000011000110;
            sine_reg0   <= 36'sb11111000100101101001001110100011000;
        end
        3468: begin
            cosine_reg0 <= 36'sb111101000011110011101000011001100;
            sine_reg0   <= 36'sb11111000100111001001001101101101010;
        end
        3469: begin
            cosine_reg0 <= 36'sb111100111101101101000110000011100;
            sine_reg0   <= 36'sb11111000101000101001000011010010001;
        end
        3470: begin
            cosine_reg0 <= 36'sb111100110111100110100001010111001;
            sine_reg0   <= 36'sb11111000101010001000101111010001100;
        end
        3471: begin
            cosine_reg0 <= 36'sb111100110001011111111010010100101;
            sine_reg0   <= 36'sb11111000101011101000010001101011011;
        end
        3472: begin
            cosine_reg0 <= 36'sb111100101011011001010000111100001;
            sine_reg0   <= 36'sb11111000101101000111101010011111101;
        end
        3473: begin
            cosine_reg0 <= 36'sb111100100101010010100101001101111;
            sine_reg0   <= 36'sb11111000101110100110111001101110001;
        end
        3474: begin
            cosine_reg0 <= 36'sb111100011111001011110111001010001;
            sine_reg0   <= 36'sb11111000110000000101111111010111000;
        end
        3475: begin
            cosine_reg0 <= 36'sb111100011001000101000110110001010;
            sine_reg0   <= 36'sb11111000110001100100111011011010001;
        end
        3476: begin
            cosine_reg0 <= 36'sb111100010010111110010100000011010;
            sine_reg0   <= 36'sb11111000110011000011101101110111100;
        end
        3477: begin
            cosine_reg0 <= 36'sb111100001100110111011111000000100;
            sine_reg0   <= 36'sb11111000110100100010010110101110111;
        end
        3478: begin
            cosine_reg0 <= 36'sb111100000110110000100111101001010;
            sine_reg0   <= 36'sb11111000110110000000110110000000010;
        end
        3479: begin
            cosine_reg0 <= 36'sb111100000000101001101101111101101;
            sine_reg0   <= 36'sb11111000110111011111001011101011110;
        end
        3480: begin
            cosine_reg0 <= 36'sb111011111010100010110001111110000;
            sine_reg0   <= 36'sb11111000111000111101010111110001001;
        end
        3481: begin
            cosine_reg0 <= 36'sb111011110100011011110011101010100;
            sine_reg0   <= 36'sb11111000111010011011011010010000011;
        end
        3482: begin
            cosine_reg0 <= 36'sb111011101110010100110011000011011;
            sine_reg0   <= 36'sb11111000111011111001010011001001100;
        end
        3483: begin
            cosine_reg0 <= 36'sb111011101000001101110000001001000;
            sine_reg0   <= 36'sb11111000111101010111000010011100100;
        end
        3484: begin
            cosine_reg0 <= 36'sb111011100010000110101010111011011;
            sine_reg0   <= 36'sb11111000111110110100101000001001000;
        end
        3485: begin
            cosine_reg0 <= 36'sb111011011011111111100011011010111;
            sine_reg0   <= 36'sb11111001000000010010000100001111011;
        end
        3486: begin
            cosine_reg0 <= 36'sb111011010101111000011001100111110;
            sine_reg0   <= 36'sb11111001000001101111010110101111010;
        end
        3487: begin
            cosine_reg0 <= 36'sb111011001111110001001101100010010;
            sine_reg0   <= 36'sb11111001000011001100011111101000101;
        end
        3488: begin
            cosine_reg0 <= 36'sb111011001001101001111111001010100;
            sine_reg0   <= 36'sb11111001000100101001011110111011101;
        end
        3489: begin
            cosine_reg0 <= 36'sb111011000011100010101110100000111;
            sine_reg0   <= 36'sb11111001000110000110010100101000000;
        end
        3490: begin
            cosine_reg0 <= 36'sb111010111101011011011011100101100;
            sine_reg0   <= 36'sb11111001000111100011000000101101101;
        end
        3491: begin
            cosine_reg0 <= 36'sb111010110111010100000110011000101;
            sine_reg0   <= 36'sb11111001001000111111100011001100110;
        end
        3492: begin
            cosine_reg0 <= 36'sb111010110001001100101110111010100;
            sine_reg0   <= 36'sb11111001001010011011111100000101001;
        end
        3493: begin
            cosine_reg0 <= 36'sb111010101011000101010101001011011;
            sine_reg0   <= 36'sb11111001001011111000001011010110101;
        end
        3494: begin
            cosine_reg0 <= 36'sb111010100100111101111001001011100;
            sine_reg0   <= 36'sb11111001001101010100010001000001011;
        end
        3495: begin
            cosine_reg0 <= 36'sb111010011110110110011010111011000;
            sine_reg0   <= 36'sb11111001001110110000001101000101010;
        end
        3496: begin
            cosine_reg0 <= 36'sb111010011000101110111010011010011;
            sine_reg0   <= 36'sb11111001010000001011111111100010001;
        end
        3497: begin
            cosine_reg0 <= 36'sb111010010010100111010111101001100;
            sine_reg0   <= 36'sb11111001010001100111101000010111111;
        end
        3498: begin
            cosine_reg0 <= 36'sb111010001100011111110010101000111;
            sine_reg0   <= 36'sb11111001010011000011000111100110110;
        end
        3499: begin
            cosine_reg0 <= 36'sb111010000110011000001011011000110;
            sine_reg0   <= 36'sb11111001010100011110011101001110011;
        end
        3500: begin
            cosine_reg0 <= 36'sb111010000000010000100001111001001;
            sine_reg0   <= 36'sb11111001010101111001101001001110111;
        end
        3501: begin
            cosine_reg0 <= 36'sb111001111010001000110110001010100;
            sine_reg0   <= 36'sb11111001010111010100101011101000010;
        end
        3502: begin
            cosine_reg0 <= 36'sb111001110100000001001000001101000;
            sine_reg0   <= 36'sb11111001011000101111100100011010010;
        end
        3503: begin
            cosine_reg0 <= 36'sb111001101101111001011000000000110;
            sine_reg0   <= 36'sb11111001011010001010010011100100111;
        end
        3504: begin
            cosine_reg0 <= 36'sb111001100111110001100101100110001;
            sine_reg0   <= 36'sb11111001011011100100111001001000001;
        end
        3505: begin
            cosine_reg0 <= 36'sb111001100001101001110000111101011;
            sine_reg0   <= 36'sb11111001011100111111010101000100000;
        end
        3506: begin
            cosine_reg0 <= 36'sb111001011011100001111010000110101;
            sine_reg0   <= 36'sb11111001011110011001100111011000010;
        end
        3507: begin
            cosine_reg0 <= 36'sb111001010101011010000001000010001;
            sine_reg0   <= 36'sb11111001011111110011110000000101001;
        end
        3508: begin
            cosine_reg0 <= 36'sb111001001111010010000101110000010;
            sine_reg0   <= 36'sb11111001100001001101101111001010010;
        end
        3509: begin
            cosine_reg0 <= 36'sb111001001001001010001000010001001;
            sine_reg0   <= 36'sb11111001100010100111100100100111110;
        end
        3510: begin
            cosine_reg0 <= 36'sb111001000011000010001000100101000;
            sine_reg0   <= 36'sb11111001100100000001010000011101100;
        end
        3511: begin
            cosine_reg0 <= 36'sb111000111100111010000110101100001;
            sine_reg0   <= 36'sb11111001100101011010110010101011100;
        end
        3512: begin
            cosine_reg0 <= 36'sb111000110110110010000010100110110;
            sine_reg0   <= 36'sb11111001100110110100001011010001110;
        end
        3513: begin
            cosine_reg0 <= 36'sb111000110000101001111100010101000;
            sine_reg0   <= 36'sb11111001101000001101011010010000000;
        end
        3514: begin
            cosine_reg0 <= 36'sb111000101010100001110011110111010;
            sine_reg0   <= 36'sb11111001101001100110011111100110011;
        end
        3515: begin
            cosine_reg0 <= 36'sb111000100100011001101001001101110;
            sine_reg0   <= 36'sb11111001101010111111011011010100110;
        end
        3516: begin
            cosine_reg0 <= 36'sb111000011110010001011100011000101;
            sine_reg0   <= 36'sb11111001101100011000001101011011001;
        end
        3517: begin
            cosine_reg0 <= 36'sb111000011000001001001101011000001;
            sine_reg0   <= 36'sb11111001101101110000110101111001011;
        end
        3518: begin
            cosine_reg0 <= 36'sb111000010010000000111100001100100;
            sine_reg0   <= 36'sb11111001101111001001010100101111100;
        end
        3519: begin
            cosine_reg0 <= 36'sb111000001011111000101000110110000;
            sine_reg0   <= 36'sb11111001110000100001101001111101011;
        end
        3520: begin
            cosine_reg0 <= 36'sb111000000101110000010011010101000;
            sine_reg0   <= 36'sb11111001110001111001110101100011000;
        end
        3521: begin
            cosine_reg0 <= 36'sb110111111111100111111011101001100;
            sine_reg0   <= 36'sb11111001110011010001110111100000011;
        end
        3522: begin
            cosine_reg0 <= 36'sb110111111001011111100001110011111;
            sine_reg0   <= 36'sb11111001110100101001101111110101011;
        end
        3523: begin
            cosine_reg0 <= 36'sb110111110011010111000101110100010;
            sine_reg0   <= 36'sb11111001110110000001011110100001111;
        end
        3524: begin
            cosine_reg0 <= 36'sb110111101101001110100111101011000;
            sine_reg0   <= 36'sb11111001110111011001000011100110000;
        end
        3525: begin
            cosine_reg0 <= 36'sb110111100111000110000111011000010;
            sine_reg0   <= 36'sb11111001111000110000011111000001101;
        end
        3526: begin
            cosine_reg0 <= 36'sb110111100000111101100100111100011;
            sine_reg0   <= 36'sb11111001111010000111110000110100101;
        end
        3527: begin
            cosine_reg0 <= 36'sb110111011010110101000000010111100;
            sine_reg0   <= 36'sb11111001111011011110111000111111000;
        end
        3528: begin
            cosine_reg0 <= 36'sb110111010100101100011001101001111;
            sine_reg0   <= 36'sb11111001111100110101110111100000110;
        end
        3529: begin
            cosine_reg0 <= 36'sb110111001110100011110000110011110;
            sine_reg0   <= 36'sb11111001111110001100101100011001110;
        end
        3530: begin
            cosine_reg0 <= 36'sb110111001000011011000101110101010;
            sine_reg0   <= 36'sb11111001111111100011010111101010000;
        end
        3531: begin
            cosine_reg0 <= 36'sb110111000010010010011000101110111;
            sine_reg0   <= 36'sb11111010000000111001111001010001011;
        end
        3532: begin
            cosine_reg0 <= 36'sb110110111100001001101001100000101;
            sine_reg0   <= 36'sb11111010000010010000010001001111110;
        end
        3533: begin
            cosine_reg0 <= 36'sb110110110110000000111000001010111;
            sine_reg0   <= 36'sb11111010000011100110011111100101011;
        end
        3534: begin
            cosine_reg0 <= 36'sb110110101111111000000100101101110;
            sine_reg0   <= 36'sb11111010000100111100100100010001111;
        end
        3535: begin
            cosine_reg0 <= 36'sb110110101001101111001111001001100;
            sine_reg0   <= 36'sb11111010000110010010011111010101011;
        end
        3536: begin
            cosine_reg0 <= 36'sb110110100011100110010111011110100;
            sine_reg0   <= 36'sb11111010000111101000010000101111111;
        end
        3537: begin
            cosine_reg0 <= 36'sb110110011101011101011101101100110;
            sine_reg0   <= 36'sb11111010001000111101111000100001001;
        end
        3538: begin
            cosine_reg0 <= 36'sb110110010111010100100001110100110;
            sine_reg0   <= 36'sb11111010001010010011010110101001010;
        end
        3539: begin
            cosine_reg0 <= 36'sb110110010001001011100011110110101;
            sine_reg0   <= 36'sb11111010001011101000101011001000001;
        end
        3540: begin
            cosine_reg0 <= 36'sb110110001011000010100011110010100;
            sine_reg0   <= 36'sb11111010001100111101110101111101101;
        end
        3541: begin
            cosine_reg0 <= 36'sb110110000100111001100001101000110;
            sine_reg0   <= 36'sb11111010001110010010110111001001110;
        end
        3542: begin
            cosine_reg0 <= 36'sb110101111110110000011101011001101;
            sine_reg0   <= 36'sb11111010001111100111101110101100101;
        end
        3543: begin
            cosine_reg0 <= 36'sb110101111000100111010111000101010;
            sine_reg0   <= 36'sb11111010010000111100011100100110000;
        end
        3544: begin
            cosine_reg0 <= 36'sb110101110010011110001110101011111;
            sine_reg0   <= 36'sb11111010010010010001000000110101110;
        end
        3545: begin
            cosine_reg0 <= 36'sb110101101100010101000100001101111;
            sine_reg0   <= 36'sb11111010010011100101011011011100000;
        end
        3546: begin
            cosine_reg0 <= 36'sb110101100110001011110111101011011;
            sine_reg0   <= 36'sb11111010010100111001101100011000110;
        end
        3547: begin
            cosine_reg0 <= 36'sb110101100000000010101001000100100;
            sine_reg0   <= 36'sb11111010010110001101110011101011110;
        end
        3548: begin
            cosine_reg0 <= 36'sb110101011001111001011000011001110;
            sine_reg0   <= 36'sb11111010010111100001110001010101000;
        end
        3549: begin
            cosine_reg0 <= 36'sb110101010011110000000101101011010;
            sine_reg0   <= 36'sb11111010011000110101100101010100101;
        end
        3550: begin
            cosine_reg0 <= 36'sb110101001101100110110000111001001;
            sine_reg0   <= 36'sb11111010011010001001001111101010011;
        end
        3551: begin
            cosine_reg0 <= 36'sb110101000111011101011010000011110;
            sine_reg0   <= 36'sb11111010011011011100110000010110010;
        end
        3552: begin
            cosine_reg0 <= 36'sb110101000001010100000001001011011;
            sine_reg0   <= 36'sb11111010011100110000000111011000010;
        end
        3553: begin
            cosine_reg0 <= 36'sb110100111011001010100110010000001;
            sine_reg0   <= 36'sb11111010011110000011010100110000010;
        end
        3554: begin
            cosine_reg0 <= 36'sb110100110101000001001001010010010;
            sine_reg0   <= 36'sb11111010011111010110011000011110010;
        end
        3555: begin
            cosine_reg0 <= 36'sb110100101110110111101010010010000;
            sine_reg0   <= 36'sb11111010100000101001010010100010010;
        end
        3556: begin
            cosine_reg0 <= 36'sb110100101000101110001001001111110;
            sine_reg0   <= 36'sb11111010100001111100000010111100000;
        end
        3557: begin
            cosine_reg0 <= 36'sb110100100010100100100110001011101;
            sine_reg0   <= 36'sb11111010100011001110101001101011110;
        end
        3558: begin
            cosine_reg0 <= 36'sb110100011100011011000001000101110;
            sine_reg0   <= 36'sb11111010100100100001000110110001010;
        end
        3559: begin
            cosine_reg0 <= 36'sb110100010110010001011001111110100;
            sine_reg0   <= 36'sb11111010100101110011011010001100100;
        end
        3560: begin
            cosine_reg0 <= 36'sb110100010000000111110000110110001;
            sine_reg0   <= 36'sb11111010100111000101100011111101011;
        end
        3561: begin
            cosine_reg0 <= 36'sb110100001001111110000101101100111;
            sine_reg0   <= 36'sb11111010101000010111100100000011111;
        end
        3562: begin
            cosine_reg0 <= 36'sb110100000011110100011000100010111;
            sine_reg0   <= 36'sb11111010101001101001011010100000000;
        end
        3563: begin
            cosine_reg0 <= 36'sb110011111101101010101001011000011;
            sine_reg0   <= 36'sb11111010101010111011000111010001110;
        end
        3564: begin
            cosine_reg0 <= 36'sb110011110111100000111000001101110;
            sine_reg0   <= 36'sb11111010101100001100101010011000111;
        end
        3565: begin
            cosine_reg0 <= 36'sb110011110001010111000101000011001;
            sine_reg0   <= 36'sb11111010101101011110000011110101101;
        end
        3566: begin
            cosine_reg0 <= 36'sb110011101011001101001111111000110;
            sine_reg0   <= 36'sb11111010101110101111010011100111101;
        end
        3567: begin
            cosine_reg0 <= 36'sb110011100101000011011000101110111;
            sine_reg0   <= 36'sb11111010110000000000011001101111000;
        end
        3568: begin
            cosine_reg0 <= 36'sb110011011110111001011111100101110;
            sine_reg0   <= 36'sb11111010110001010001010110001011101;
        end
        3569: begin
            cosine_reg0 <= 36'sb110011011000101111100100011101100;
            sine_reg0   <= 36'sb11111010110010100010001000111101101;
        end
        3570: begin
            cosine_reg0 <= 36'sb110011010010100101100111010110100;
            sine_reg0   <= 36'sb11111010110011110010110010000100110;
        end
        3571: begin
            cosine_reg0 <= 36'sb110011001100011011101000010001000;
            sine_reg0   <= 36'sb11111010110101000011010001100001000;
        end
        3572: begin
            cosine_reg0 <= 36'sb110011000110010001100111001101001;
            sine_reg0   <= 36'sb11111010110110010011100111010010011;
        end
        3573: begin
            cosine_reg0 <= 36'sb110011000000000111100100001011010;
            sine_reg0   <= 36'sb11111010110111100011110011011000110;
        end
        3574: begin
            cosine_reg0 <= 36'sb110010111001111101011111001011100;
            sine_reg0   <= 36'sb11111010111000110011110101110100010;
        end
        3575: begin
            cosine_reg0 <= 36'sb110010110011110011011000001110001;
            sine_reg0   <= 36'sb11111010111010000011101110100100101;
        end
        3576: begin
            cosine_reg0 <= 36'sb110010101101101001001111010011011;
            sine_reg0   <= 36'sb11111010111011010011011101101010000;
        end
        3577: begin
            cosine_reg0 <= 36'sb110010100111011111000100011011100;
            sine_reg0   <= 36'sb11111010111100100011000011000100001;
        end
        3578: begin
            cosine_reg0 <= 36'sb110010100001010100110111100110110;
            sine_reg0   <= 36'sb11111010111101110010011110110011001;
        end
        3579: begin
            cosine_reg0 <= 36'sb110010011011001010101000110101011;
            sine_reg0   <= 36'sb11111010111111000001110000110110111;
        end
        3580: begin
            cosine_reg0 <= 36'sb110010010101000000011000000111100;
            sine_reg0   <= 36'sb11111011000000010000111001001111011;
        end
        3581: begin
            cosine_reg0 <= 36'sb110010001110110110000101011101100;
            sine_reg0   <= 36'sb11111011000001011111110111111100101;
        end
        3582: begin
            cosine_reg0 <= 36'sb110010001000101011110000110111101;
            sine_reg0   <= 36'sb11111011000010101110101100111110011;
        end
        3583: begin
            cosine_reg0 <= 36'sb110010000010100001011010010101111;
            sine_reg0   <= 36'sb11111011000011111101011000010100110;
        end
        3584: begin
            cosine_reg0 <= 36'sb110001111100010111000001111000110;
            sine_reg0   <= 36'sb11111011000101001011111001111111101;
        end
        3585: begin
            cosine_reg0 <= 36'sb110001110110001100100111100000100;
            sine_reg0   <= 36'sb11111011000110011010010001111111000;
        end
        3586: begin
            cosine_reg0 <= 36'sb110001110000000010001011001101001;
            sine_reg0   <= 36'sb11111011000111101000100000010010110;
        end
        3587: begin
            cosine_reg0 <= 36'sb110001101001110111101100111111000;
            sine_reg0   <= 36'sb11111011001000110110100100111011000;
        end
        3588: begin
            cosine_reg0 <= 36'sb110001100011101101001100110110011;
            sine_reg0   <= 36'sb11111011001010000100011111110111100;
        end
        3589: begin
            cosine_reg0 <= 36'sb110001011101100010101010110011100;
            sine_reg0   <= 36'sb11111011001011010010010001001000011;
        end
        3590: begin
            cosine_reg0 <= 36'sb110001010111011000000110110110100;
            sine_reg0   <= 36'sb11111011001100011111111000101101011;
        end
        3591: begin
            cosine_reg0 <= 36'sb110001010001001101100000111111111;
            sine_reg0   <= 36'sb11111011001101101101010110100110110;
        end
        3592: begin
            cosine_reg0 <= 36'sb110001001011000010111001001111100;
            sine_reg0   <= 36'sb11111011001110111010101010110100001;
        end
        3593: begin
            cosine_reg0 <= 36'sb110001000100111000001111100101111;
            sine_reg0   <= 36'sb11111011010000000111110101010101101;
        end
        3594: begin
            cosine_reg0 <= 36'sb110000111110101101100100000011001;
            sine_reg0   <= 36'sb11111011010001010100110110001011010;
        end
        3595: begin
            cosine_reg0 <= 36'sb110000111000100010110110100111101;
            sine_reg0   <= 36'sb11111011010010100001101101010100111;
        end
        3596: begin
            cosine_reg0 <= 36'sb110000110010011000000111010011011;
            sine_reg0   <= 36'sb11111011010011101110011010110010100;
        end
        3597: begin
            cosine_reg0 <= 36'sb110000101100001101010110000110110;
            sine_reg0   <= 36'sb11111011010100111010111110100100000;
        end
        3598: begin
            cosine_reg0 <= 36'sb110000100110000010100011000010001;
            sine_reg0   <= 36'sb11111011010110000111011000101001011;
        end
        3599: begin
            cosine_reg0 <= 36'sb110000011111110111101110000101100;
            sine_reg0   <= 36'sb11111011010111010011101001000010101;
        end
        3600: begin
            cosine_reg0 <= 36'sb110000011001101100110111010001010;
            sine_reg0   <= 36'sb11111011011000011111101111101111100;
        end
        3601: begin
            cosine_reg0 <= 36'sb110000010011100001111110100101100;
            sine_reg0   <= 36'sb11111011011001101011101100110000010;
        end
        3602: begin
            cosine_reg0 <= 36'sb110000001101010111000100000010101;
            sine_reg0   <= 36'sb11111011011010110111100000000100110;
        end
        3603: begin
            cosine_reg0 <= 36'sb110000000111001100000111101000110;
            sine_reg0   <= 36'sb11111011011100000011001001101100110;
        end
        3604: begin
            cosine_reg0 <= 36'sb110000000001000001001001011000010;
            sine_reg0   <= 36'sb11111011011101001110101001101000100;
        end
        3605: begin
            cosine_reg0 <= 36'sb101111111010110110001001010001001;
            sine_reg0   <= 36'sb11111011011110011001111111110111101;
        end
        3606: begin
            cosine_reg0 <= 36'sb101111110100101011000111010011111;
            sine_reg0   <= 36'sb11111011011111100101001100011010011;
        end
        3607: begin
            cosine_reg0 <= 36'sb101111101110100000000011100000101;
            sine_reg0   <= 36'sb11111011100000110000001111010000101;
        end
        3608: begin
            cosine_reg0 <= 36'sb101111101000010100111101110111101;
            sine_reg0   <= 36'sb11111011100001111011001000011010010;
        end
        3609: begin
            cosine_reg0 <= 36'sb101111100010001001110110011001001;
            sine_reg0   <= 36'sb11111011100011000101110111110111010;
        end
        3610: begin
            cosine_reg0 <= 36'sb101111011011111110101101000101010;
            sine_reg0   <= 36'sb11111011100100010000011101100111100;
        end
        3611: begin
            cosine_reg0 <= 36'sb101111010101110011100001111100011;
            sine_reg0   <= 36'sb11111011100101011010111001101011001;
        end
        3612: begin
            cosine_reg0 <= 36'sb101111001111101000010100111110101;
            sine_reg0   <= 36'sb11111011100110100101001100000010000;
        end
        3613: begin
            cosine_reg0 <= 36'sb101111001001011101000110001100011;
            sine_reg0   <= 36'sb11111011100111101111010100101100000;
        end
        3614: begin
            cosine_reg0 <= 36'sb101111000011010001110101100101111;
            sine_reg0   <= 36'sb11111011101000111001010011101001010;
        end
        3615: begin
            cosine_reg0 <= 36'sb101110111101000110100011001011001;
            sine_reg0   <= 36'sb11111011101010000011001000111001100;
        end
        3616: begin
            cosine_reg0 <= 36'sb101110110110111011001110111100101;
            sine_reg0   <= 36'sb11111011101011001100110100011100111;
        end
        3617: begin
            cosine_reg0 <= 36'sb101110110000101111111000111010100;
            sine_reg0   <= 36'sb11111011101100010110010110010011010;
        end
        3618: begin
            cosine_reg0 <= 36'sb101110101010100100100001000100111;
            sine_reg0   <= 36'sb11111011101101011111101110011100101;
        end
        3619: begin
            cosine_reg0 <= 36'sb101110100100011001000111011100010;
            sine_reg0   <= 36'sb11111011101110101000111100111000111;
        end
        3620: begin
            cosine_reg0 <= 36'sb101110011110001101101100000000101;
            sine_reg0   <= 36'sb11111011101111110010000001101000001;
        end
        3621: begin
            cosine_reg0 <= 36'sb101110011000000010001110110010011;
            sine_reg0   <= 36'sb11111011110000111010111100101010001;
        end
        3622: begin
            cosine_reg0 <= 36'sb101110010001110110101111110001110;
            sine_reg0   <= 36'sb11111011110010000011101101111110111;
        end
        3623: begin
            cosine_reg0 <= 36'sb101110001011101011001110111110111;
            sine_reg0   <= 36'sb11111011110011001100010101100110011;
        end
        3624: begin
            cosine_reg0 <= 36'sb101110000101011111101100011010000;
            sine_reg0   <= 36'sb11111011110100010100110011100000110;
        end
        3625: begin
            cosine_reg0 <= 36'sb101101111111010100001000000011100;
            sine_reg0   <= 36'sb11111011110101011101000111101101101;
        end
        3626: begin
            cosine_reg0 <= 36'sb101101111001001000100001111011100;
            sine_reg0   <= 36'sb11111011110110100101010010001101001;
        end
        3627: begin
            cosine_reg0 <= 36'sb101101110010111100111010000010010;
            sine_reg0   <= 36'sb11111011110111101101010010111111010;
        end
        3628: begin
            cosine_reg0 <= 36'sb101101101100110001010000011000000;
            sine_reg0   <= 36'sb11111011111000110101001010000100000;
        end
        3629: begin
            cosine_reg0 <= 36'sb101101100110100101100100111101000;
            sine_reg0   <= 36'sb11111011111001111100110111011011001;
        end
        3630: begin
            cosine_reg0 <= 36'sb101101100000011001110111110001100;
            sine_reg0   <= 36'sb11111011111011000100011011000100110;
        end
        3631: begin
            cosine_reg0 <= 36'sb101101011010001110001000110101110;
            sine_reg0   <= 36'sb11111011111100001011110101000000110;
        end
        3632: begin
            cosine_reg0 <= 36'sb101101010100000010011000001001111;
            sine_reg0   <= 36'sb11111011111101010011000101001111001;
        end
        3633: begin
            cosine_reg0 <= 36'sb101101001101110110100101101110010;
            sine_reg0   <= 36'sb11111011111110011010001011101111110;
        end
        3634: begin
            cosine_reg0 <= 36'sb101101000111101010110001100011000;
            sine_reg0   <= 36'sb11111011111111100001001000100010110;
        end
        3635: begin
            cosine_reg0 <= 36'sb101101000001011110111011101000100;
            sine_reg0   <= 36'sb11111100000000100111111011100111111;
        end
        3636: begin
            cosine_reg0 <= 36'sb101100111011010011000011111110111;
            sine_reg0   <= 36'sb11111100000001101110100100111111010;
        end
        3637: begin
            cosine_reg0 <= 36'sb101100110101000111001010100110011;
            sine_reg0   <= 36'sb11111100000010110101000100101000111;
        end
        3638: begin
            cosine_reg0 <= 36'sb101100101110111011001111011111010;
            sine_reg0   <= 36'sb11111100000011111011011010100100100;
        end
        3639: begin
            cosine_reg0 <= 36'sb101100101000101111010010101001111;
            sine_reg0   <= 36'sb11111100000101000001100110110010001;
        end
        3640: begin
            cosine_reg0 <= 36'sb101100100010100011010100000110010;
            sine_reg0   <= 36'sb11111100000110000111101001010001111;
        end
        3641: begin
            cosine_reg0 <= 36'sb101100011100010111010011110100110;
            sine_reg0   <= 36'sb11111100000111001101100010000011101;
        end
        3642: begin
            cosine_reg0 <= 36'sb101100010110001011010001110101100;
            sine_reg0   <= 36'sb11111100001000010011010001000111010;
        end
        3643: begin
            cosine_reg0 <= 36'sb101100001111111111001110001001000;
            sine_reg0   <= 36'sb11111100001001011000110110011100110;
        end
        3644: begin
            cosine_reg0 <= 36'sb101100001001110011001000101111001;
            sine_reg0   <= 36'sb11111100001010011110010010000100001;
        end
        3645: begin
            cosine_reg0 <= 36'sb101100000011100111000001101000100;
            sine_reg0   <= 36'sb11111100001011100011100011111101011;
        end
        3646: begin
            cosine_reg0 <= 36'sb101011111101011010111000110101000;
            sine_reg0   <= 36'sb11111100001100101000101100001000011;
        end
        3647: begin
            cosine_reg0 <= 36'sb101011110111001110101110010101001;
            sine_reg0   <= 36'sb11111100001101101101101010100101000;
        end
        3648: begin
            cosine_reg0 <= 36'sb101011110001000010100010001001001;
            sine_reg0   <= 36'sb11111100001110110010011111010011011;
        end
        3649: begin
            cosine_reg0 <= 36'sb101011101010110110010100010001000;
            sine_reg0   <= 36'sb11111100001111110111001010010011100;
        end
        3650: begin
            cosine_reg0 <= 36'sb101011100100101010000100101101001;
            sine_reg0   <= 36'sb11111100010000111011101011100101001;
        end
        3651: begin
            cosine_reg0 <= 36'sb101011011110011101110011011101110;
            sine_reg0   <= 36'sb11111100010010000000000011001000010;
        end
        3652: begin
            cosine_reg0 <= 36'sb101011011000010001100000100011001;
            sine_reg0   <= 36'sb11111100010011000100010000111101000;
        end
        3653: begin
            cosine_reg0 <= 36'sb101011010010000101001011111101100;
            sine_reg0   <= 36'sb11111100010100001000010101000011001;
        end
        3654: begin
            cosine_reg0 <= 36'sb101011001011111000110101101101000;
            sine_reg0   <= 36'sb11111100010101001100001111011010110;
        end
        3655: begin
            cosine_reg0 <= 36'sb101011000101101100011101110010000;
            sine_reg0   <= 36'sb11111100010110010000000000000011111;
        end
        3656: begin
            cosine_reg0 <= 36'sb101010111111100000000100001100101;
            sine_reg0   <= 36'sb11111100010111010011100110111110010;
        end
        3657: begin
            cosine_reg0 <= 36'sb101010111001010011101000111101010;
            sine_reg0   <= 36'sb11111100011000010111000100001001111;
        end
        3658: begin
            cosine_reg0 <= 36'sb101010110011000111001100000100000;
            sine_reg0   <= 36'sb11111100011001011010010111100110111;
        end
        3659: begin
            cosine_reg0 <= 36'sb101010101100111010101101100001001;
            sine_reg0   <= 36'sb11111100011010011101100001010101001;
        end
        3660: begin
            cosine_reg0 <= 36'sb101010100110101110001101010100111;
            sine_reg0   <= 36'sb11111100011011100000100001010100100;
        end
        3661: begin
            cosine_reg0 <= 36'sb101010100000100001101011011111100;
            sine_reg0   <= 36'sb11111100011100100011010111100101001;
        end
        3662: begin
            cosine_reg0 <= 36'sb101010011010010101001000000001011;
            sine_reg0   <= 36'sb11111100011101100110000100000110110;
        end
        3663: begin
            cosine_reg0 <= 36'sb101010010100001000100010111010100;
            sine_reg0   <= 36'sb11111100011110101000100110111001100;
        end
        3664: begin
            cosine_reg0 <= 36'sb101010001101111011111100001011001;
            sine_reg0   <= 36'sb11111100011111101010111111111101011;
        end
        3665: begin
            cosine_reg0 <= 36'sb101010000111101111010011110011110;
            sine_reg0   <= 36'sb11111100100000101101001111010010001;
        end
        3666: begin
            cosine_reg0 <= 36'sb101010000001100010101001110100011;
            sine_reg0   <= 36'sb11111100100001101111010100110111111;
        end
        3667: begin
            cosine_reg0 <= 36'sb101001111011010101111110001101010;
            sine_reg0   <= 36'sb11111100100010110001010000101110100;
        end
        3668: begin
            cosine_reg0 <= 36'sb101001110101001001010000111110110;
            sine_reg0   <= 36'sb11111100100011110011000010110110000;
        end
        3669: begin
            cosine_reg0 <= 36'sb101001101110111100100010001001000;
            sine_reg0   <= 36'sb11111100100100110100101011001110011;
        end
        3670: begin
            cosine_reg0 <= 36'sb101001101000101111110001101100010;
            sine_reg0   <= 36'sb11111100100101110110001001110111100;
        end
        3671: begin
            cosine_reg0 <= 36'sb101001100010100010111111101000111;
            sine_reg0   <= 36'sb11111100100110110111011110110001011;
        end
        3672: begin
            cosine_reg0 <= 36'sb101001011100010110001011111110111;
            sine_reg0   <= 36'sb11111100100111111000101001111100000;
        end
        3673: begin
            cosine_reg0 <= 36'sb101001010110001001010110101110110;
            sine_reg0   <= 36'sb11111100101000111001101011010111011;
        end
        3674: begin
            cosine_reg0 <= 36'sb101001001111111100011111111000100;
            sine_reg0   <= 36'sb11111100101001111010100011000011010;
        end
        3675: begin
            cosine_reg0 <= 36'sb101001001001101111100111011100100;
            sine_reg0   <= 36'sb11111100101010111011010000111111111;
        end
        3676: begin
            cosine_reg0 <= 36'sb101001000011100010101101011011000;
            sine_reg0   <= 36'sb11111100101011111011110101001100111;
        end
        3677: begin
            cosine_reg0 <= 36'sb101000111101010101110001110100010;
            sine_reg0   <= 36'sb11111100101100111100001111101010100;
        end
        3678: begin
            cosine_reg0 <= 36'sb101000110111001000110100101000010;
            sine_reg0   <= 36'sb11111100101101111100100000011000101;
        end
        3679: begin
            cosine_reg0 <= 36'sb101000110000111011110101110111101;
            sine_reg0   <= 36'sb11111100101110111100100111010111010;
        end
        3680: begin
            cosine_reg0 <= 36'sb101000101010101110110101100010010;
            sine_reg0   <= 36'sb11111100101111111100100100100110001;
        end
        3681: begin
            cosine_reg0 <= 36'sb101000100100100001110011101000101;
            sine_reg0   <= 36'sb11111100110000111100011000000101100;
        end
        3682: begin
            cosine_reg0 <= 36'sb101000011110010100110000001010111;
            sine_reg0   <= 36'sb11111100110001111100000001110101001;
        end
        3683: begin
            cosine_reg0 <= 36'sb101000011000000111101011001001011;
            sine_reg0   <= 36'sb11111100110010111011100001110101000;
        end
        3684: begin
            cosine_reg0 <= 36'sb101000010001111010100100100100001;
            sine_reg0   <= 36'sb11111100110011111010111000000101010;
        end
        3685: begin
            cosine_reg0 <= 36'sb101000001011101101011100011011100;
            sine_reg0   <= 36'sb11111100110100111010000100100101101;
        end
        3686: begin
            cosine_reg0 <= 36'sb101000000101100000010010101111110;
            sine_reg0   <= 36'sb11111100110101111001000111010110010;
        end
        3687: begin
            cosine_reg0 <= 36'sb100111111111010011000111100001000;
            sine_reg0   <= 36'sb11111100110110111000000000010110111;
        end
        3688: begin
            cosine_reg0 <= 36'sb100111111001000101111010101111110;
            sine_reg0   <= 36'sb11111100110111110110101111100111110;
        end
        3689: begin
            cosine_reg0 <= 36'sb100111110010111000101100011011111;
            sine_reg0   <= 36'sb11111100111000110101010101001000101;
        end
        3690: begin
            cosine_reg0 <= 36'sb100111101100101011011100100110000;
            sine_reg0   <= 36'sb11111100111001110011110000111001100;
        end
        3691: begin
            cosine_reg0 <= 36'sb100111100110011110001011001110000;
            sine_reg0   <= 36'sb11111100111010110010000010111010011;
        end
        3692: begin
            cosine_reg0 <= 36'sb100111100000010000111000010100011;
            sine_reg0   <= 36'sb11111100111011110000001011001011010;
        end
        3693: begin
            cosine_reg0 <= 36'sb100111011010000011100011111001011;
            sine_reg0   <= 36'sb11111100111100101110001001101100000;
        end
        3694: begin
            cosine_reg0 <= 36'sb100111010011110110001101111101000;
            sine_reg0   <= 36'sb11111100111101101011111110011100101;
        end
        3695: begin
            cosine_reg0 <= 36'sb100111001101101000110110011111101;
            sine_reg0   <= 36'sb11111100111110101001101001011101000;
        end
        3696: begin
            cosine_reg0 <= 36'sb100111000111011011011101100001101;
            sine_reg0   <= 36'sb11111100111111100111001010101101010;
        end
        3697: begin
            cosine_reg0 <= 36'sb100111000001001110000011000011000;
            sine_reg0   <= 36'sb11111101000000100100100010001101011;
        end
        3698: begin
            cosine_reg0 <= 36'sb100110111011000000100111000100001;
            sine_reg0   <= 36'sb11111101000001100001101111111101001;
        end
        3699: begin
            cosine_reg0 <= 36'sb100110110100110011001001100101010;
            sine_reg0   <= 36'sb11111101000010011110110011111100100;
        end
        3700: begin
            cosine_reg0 <= 36'sb100110101110100101101010100110100;
            sine_reg0   <= 36'sb11111101000011011011101110001011101;
        end
        3701: begin
            cosine_reg0 <= 36'sb100110101000011000001010001000010;
            sine_reg0   <= 36'sb11111101000100011000011110101010010;
        end
        3702: begin
            cosine_reg0 <= 36'sb100110100010001010101000001010101;
            sine_reg0   <= 36'sb11111101000101010101000101011000100;
        end
        3703: begin
            cosine_reg0 <= 36'sb100110011011111101000100101110000;
            sine_reg0   <= 36'sb11111101000110010001100010010110011;
        end
        3704: begin
            cosine_reg0 <= 36'sb100110010101101111011111110010100;
            sine_reg0   <= 36'sb11111101000111001101110101100011110;
        end
        3705: begin
            cosine_reg0 <= 36'sb100110001111100001111001011000011;
            sine_reg0   <= 36'sb11111101001000001001111111000000100;
        end
        3706: begin
            cosine_reg0 <= 36'sb100110001001010100010001100000000;
            sine_reg0   <= 36'sb11111101001001000101111110101100110;
        end
        3707: begin
            cosine_reg0 <= 36'sb100110000011000110101000001001011;
            sine_reg0   <= 36'sb11111101001010000001110100101000011;
        end
        3708: begin
            cosine_reg0 <= 36'sb100101111100111000111101010101000;
            sine_reg0   <= 36'sb11111101001010111101100000110011011;
        end
        3709: begin
            cosine_reg0 <= 36'sb100101110110101011010001000010111;
            sine_reg0   <= 36'sb11111101001011111001000011001101101;
        end
        3710: begin
            cosine_reg0 <= 36'sb100101110000011101100011010011011;
            sine_reg0   <= 36'sb11111101001100110100011011110111010;
        end
        3711: begin
            cosine_reg0 <= 36'sb100101101010001111110100000110101;
            sine_reg0   <= 36'sb11111101001101101111101010110000001;
        end
        3712: begin
            cosine_reg0 <= 36'sb100101100100000010000011011101001;
            sine_reg0   <= 36'sb11111101001110101010101111111000001;
        end
        3713: begin
            cosine_reg0 <= 36'sb100101011101110100010001010110111;
            sine_reg0   <= 36'sb11111101001111100101101011001111011;
        end
        3714: begin
            cosine_reg0 <= 36'sb100101010111100110011101110100001;
            sine_reg0   <= 36'sb11111101010000100000011100110101110;
        end
        3715: begin
            cosine_reg0 <= 36'sb100101010001011000101000110101010;
            sine_reg0   <= 36'sb11111101010001011011000100101011010;
        end
        3716: begin
            cosine_reg0 <= 36'sb100101001011001010110010011010011;
            sine_reg0   <= 36'sb11111101010010010101100010101111111;
        end
        3717: begin
            cosine_reg0 <= 36'sb100101000100111100111010100011110;
            sine_reg0   <= 36'sb11111101010011001111110111000011100;
        end
        3718: begin
            cosine_reg0 <= 36'sb100100111110101111000001010001101;
            sine_reg0   <= 36'sb11111101010100001010000001100110001;
        end
        3719: begin
            cosine_reg0 <= 36'sb100100111000100001000110100100010;
            sine_reg0   <= 36'sb11111101010101000100000010010111110;
        end
        3720: begin
            cosine_reg0 <= 36'sb100100110010010011001010011100000;
            sine_reg0   <= 36'sb11111101010101111101111001011000010;
        end
        3721: begin
            cosine_reg0 <= 36'sb100100101100000101001100111000111;
            sine_reg0   <= 36'sb11111101010110110111100110100111110;
        end
        3722: begin
            cosine_reg0 <= 36'sb100100100101110111001101111011010;
            sine_reg0   <= 36'sb11111101010111110001001010000110000;
        end
        3723: begin
            cosine_reg0 <= 36'sb100100011111101001001101100011010;
            sine_reg0   <= 36'sb11111101011000101010100011110011001;
        end
        3724: begin
            cosine_reg0 <= 36'sb100100011001011011001011110001011;
            sine_reg0   <= 36'sb11111101011001100011110011101111001;
        end
        3725: begin
            cosine_reg0 <= 36'sb100100010011001101001000100101101;
            sine_reg0   <= 36'sb11111101011010011100111001111001110;
        end
        3726: begin
            cosine_reg0 <= 36'sb100100001100111111000100000000010;
            sine_reg0   <= 36'sb11111101011011010101110110010011010;
        end
        3727: begin
            cosine_reg0 <= 36'sb100100000110110000111110000001101;
            sine_reg0   <= 36'sb11111101011100001110101000111011011;
        end
        3728: begin
            cosine_reg0 <= 36'sb100100000000100010110110101001111;
            sine_reg0   <= 36'sb11111101011101000111010001110010001;
        end
        3729: begin
            cosine_reg0 <= 36'sb100011111010010100101101111001010;
            sine_reg0   <= 36'sb11111101011101111111110000110111100;
        end
        3730: begin
            cosine_reg0 <= 36'sb100011110100000110100011110000000;
            sine_reg0   <= 36'sb11111101011110111000000110001011100;
        end
        3731: begin
            cosine_reg0 <= 36'sb100011101101111000011000001110100;
            sine_reg0   <= 36'sb11111101011111110000010001101110000;
        end
        3732: begin
            cosine_reg0 <= 36'sb100011100111101010001011010100110;
            sine_reg0   <= 36'sb11111101100000101000010011011111001;
        end
        3733: begin
            cosine_reg0 <= 36'sb100011100001011011111101000011001;
            sine_reg0   <= 36'sb11111101100001100000001011011110101;
        end
        3734: begin
            cosine_reg0 <= 36'sb100011011011001101101101011001111;
            sine_reg0   <= 36'sb11111101100010010111111001101100101;
        end
        3735: begin
            cosine_reg0 <= 36'sb100011010100111111011100011001010;
            sine_reg0   <= 36'sb11111101100011001111011110001001001;
        end
        3736: begin
            cosine_reg0 <= 36'sb100011001110110001001010000001100;
            sine_reg0   <= 36'sb11111101100100000110111000110011111;
        end
        3737: begin
            cosine_reg0 <= 36'sb100011001000100010110110010010110;
            sine_reg0   <= 36'sb11111101100100111110001001101101001;
        end
        3738: begin
            cosine_reg0 <= 36'sb100011000010010100100001001101010;
            sine_reg0   <= 36'sb11111101100101110101010000110100101;
        end
        3739: begin
            cosine_reg0 <= 36'sb100010111100000110001010110001011;
            sine_reg0   <= 36'sb11111101100110101100001110001010011;
        end
        3740: begin
            cosine_reg0 <= 36'sb100010110101110111110010111111011;
            sine_reg0   <= 36'sb11111101100111100011000001101110100;
        end
        3741: begin
            cosine_reg0 <= 36'sb100010101111101001011001110111010;
            sine_reg0   <= 36'sb11111101101000011001101011100000110;
        end
        3742: begin
            cosine_reg0 <= 36'sb100010101001011010111111011001100;
            sine_reg0   <= 36'sb11111101101001010000001011100001010;
        end
        3743: begin
            cosine_reg0 <= 36'sb100010100011001100100011100110010;
            sine_reg0   <= 36'sb11111101101010000110100001101111111;
        end
        3744: begin
            cosine_reg0 <= 36'sb100010011100111110000110011101110;
            sine_reg0   <= 36'sb11111101101010111100101110001100100;
        end
        3745: begin
            cosine_reg0 <= 36'sb100010010110101111101000000000001;
            sine_reg0   <= 36'sb11111101101011110010110000110111011;
        end
        3746: begin
            cosine_reg0 <= 36'sb100010010000100001001000001101111;
            sine_reg0   <= 36'sb11111101101100101000101001110000010;
        end
        3747: begin
            cosine_reg0 <= 36'sb100010001010010010100111000111000;
            sine_reg0   <= 36'sb11111101101101011110011000110111010;
        end
        3748: begin
            cosine_reg0 <= 36'sb100010000100000100000100101011111;
            sine_reg0   <= 36'sb11111101101110010011111110001100001;
        end
        3749: begin
            cosine_reg0 <= 36'sb100001111101110101100000111100110;
            sine_reg0   <= 36'sb11111101101111001001011001101111000;
        end
        3750: begin
            cosine_reg0 <= 36'sb100001110111100110111011111001110;
            sine_reg0   <= 36'sb11111101101111111110101011011111110;
        end
        3751: begin
            cosine_reg0 <= 36'sb100001110001011000010101100011010;
            sine_reg0   <= 36'sb11111101110000110011110011011110100;
        end
        3752: begin
            cosine_reg0 <= 36'sb100001101011001001101101111001011;
            sine_reg0   <= 36'sb11111101110001101000110001101011001;
        end
        3753: begin
            cosine_reg0 <= 36'sb100001100100111011000100111100011;
            sine_reg0   <= 36'sb11111101110010011101100110000101100;
        end
        3754: begin
            cosine_reg0 <= 36'sb100001011110101100011010101100101;
            sine_reg0   <= 36'sb11111101110011010010010000101101110;
        end
        3755: begin
            cosine_reg0 <= 36'sb100001011000011101101111001010010;
            sine_reg0   <= 36'sb11111101110100000110110001100011101;
        end
        3756: begin
            cosine_reg0 <= 36'sb100001010010001111000010010101011;
            sine_reg0   <= 36'sb11111101110100111011001000100111011;
        end
        3757: begin
            cosine_reg0 <= 36'sb100001001100000000010100001110100;
            sine_reg0   <= 36'sb11111101110101101111010101111000110;
        end
        3758: begin
            cosine_reg0 <= 36'sb100001000101110001100100110101110;
            sine_reg0   <= 36'sb11111101110110100011011001010111111;
        end
        3759: begin
            cosine_reg0 <= 36'sb100000111111100010110100001011010;
            sine_reg0   <= 36'sb11111101110111010111010011000100101;
        end
        3760: begin
            cosine_reg0 <= 36'sb100000111001010100000010001111100;
            sine_reg0   <= 36'sb11111101111000001011000010111111000;
        end
        3761: begin
            cosine_reg0 <= 36'sb100000110011000101001111000010011;
            sine_reg0   <= 36'sb11111101111000111110101001000111000;
        end
        3762: begin
            cosine_reg0 <= 36'sb100000101100110110011010100100100;
            sine_reg0   <= 36'sb11111101111001110010000101011100011;
        end
        3763: begin
            cosine_reg0 <= 36'sb100000100110100111100100110101111;
            sine_reg0   <= 36'sb11111101111010100101010111111111100;
        end
        3764: begin
            cosine_reg0 <= 36'sb100000100000011000101101110110110;
            sine_reg0   <= 36'sb11111101111011011000100000110000000;
        end
        3765: begin
            cosine_reg0 <= 36'sb100000011010001001110101100111100;
            sine_reg0   <= 36'sb11111101111100001011011111101101111;
        end
        3766: begin
            cosine_reg0 <= 36'sb100000010011111010111100001000010;
            sine_reg0   <= 36'sb11111101111100111110010100111001010;
        end
        3767: begin
            cosine_reg0 <= 36'sb100000001101101100000001011001010;
            sine_reg0   <= 36'sb11111101111101110001000000010010000;
        end
        3768: begin
            cosine_reg0 <= 36'sb100000000111011101000101011010111;
            sine_reg0   <= 36'sb11111101111110100011100001111000010;
        end
        3769: begin
            cosine_reg0 <= 36'sb100000000001001110001000001101001;
            sine_reg0   <= 36'sb11111101111111010101111001101011110;
        end
        3770: begin
            cosine_reg0 <= 36'sb11111111010111111001001110000100;
            sine_reg0   <= 36'sb11111110000000001000000111101100100;
        end
        3771: begin
            cosine_reg0 <= 36'sb11111110100110000001010000101000;
            sine_reg0   <= 36'sb11111110000000111010001011111010100;
        end
        3772: begin
            cosine_reg0 <= 36'sb11111101110100001001001001011000;
            sine_reg0   <= 36'sb11111110000001101100000110010101111;
        end
        3773: begin
            cosine_reg0 <= 36'sb11111101000010010000111000010110;
            sine_reg0   <= 36'sb11111110000010011101110110111110011;
        end
        3774: begin
            cosine_reg0 <= 36'sb11111100010000011000011101100011;
            sine_reg0   <= 36'sb11111110000011001111011101110100001;
        end
        3775: begin
            cosine_reg0 <= 36'sb11111011011110011111111001000011;
            sine_reg0   <= 36'sb11111110000100000000111010110111000;
        end
        3776: begin
            cosine_reg0 <= 36'sb11111010101100100111001010110101;
            sine_reg0   <= 36'sb11111110000100110010001110000110111;
        end
        3777: begin
            cosine_reg0 <= 36'sb11111001111010101110010010111101;
            sine_reg0   <= 36'sb11111110000101100011010111100100000;
        end
        3778: begin
            cosine_reg0 <= 36'sb11111001001000110101010001011101;
            sine_reg0   <= 36'sb11111110000110010100010111001110001;
        end
        3779: begin
            cosine_reg0 <= 36'sb11111000010110111100000110010101;
            sine_reg0   <= 36'sb11111110000111000101001101000101011;
        end
        3780: begin
            cosine_reg0 <= 36'sb11110111100101000010110001101001;
            sine_reg0   <= 36'sb11111110000111110101111001001001100;
        end
        3781: begin
            cosine_reg0 <= 36'sb11110110110011001001010011011010;
            sine_reg0   <= 36'sb11111110001000100110011011011010110;
        end
        3782: begin
            cosine_reg0 <= 36'sb11110110000001001111101011101010;
            sine_reg0   <= 36'sb11111110001001010110110011111000111;
        end
        3783: begin
            cosine_reg0 <= 36'sb11110101001111010101111010011011;
            sine_reg0   <= 36'sb11111110001010000111000010100011111;
        end
        3784: begin
            cosine_reg0 <= 36'sb11110100011101011011111111101111;
            sine_reg0   <= 36'sb11111110001010110111000111011011110;
        end
        3785: begin
            cosine_reg0 <= 36'sb11110011101011100001111011101000;
            sine_reg0   <= 36'sb11111110001011100111000010100000101;
        end
        3786: begin
            cosine_reg0 <= 36'sb11110010111001100111101110000111;
            sine_reg0   <= 36'sb11111110001100010110110011110010010;
        end
        3787: begin
            cosine_reg0 <= 36'sb11110010000111101101010111001111;
            sine_reg0   <= 36'sb11111110001101000110011011010000101;
        end
        3788: begin
            cosine_reg0 <= 36'sb11110001010101110010110111000010;
            sine_reg0   <= 36'sb11111110001101110101111000111011111;
        end
        3789: begin
            cosine_reg0 <= 36'sb11110000100011111000001101100001;
            sine_reg0   <= 36'sb11111110001110100101001100110011110;
        end
        3790: begin
            cosine_reg0 <= 36'sb11101111110001111101011010101111;
            sine_reg0   <= 36'sb11111110001111010100010110111000100;
        end
        3791: begin
            cosine_reg0 <= 36'sb11101111000000000010011110101101;
            sine_reg0   <= 36'sb11111110010000000011010111001001111;
        end
        3792: begin
            cosine_reg0 <= 36'sb11101110001110000111011001011101;
            sine_reg0   <= 36'sb11111110010000110010001101100111111;
        end
        3793: begin
            cosine_reg0 <= 36'sb11101101011100001100001011000010;
            sine_reg0   <= 36'sb11111110010001100000111010010010100;
        end
        3794: begin
            cosine_reg0 <= 36'sb11101100101010010000110011011101;
            sine_reg0   <= 36'sb11111110010010001111011101001001110;
        end
        3795: begin
            cosine_reg0 <= 36'sb11101011111000010101010010101111;
            sine_reg0   <= 36'sb11111110010010111101110110001101101;
        end
        3796: begin
            cosine_reg0 <= 36'sb11101011000110011001101000111100;
            sine_reg0   <= 36'sb11111110010011101100000101011110000;
        end
        3797: begin
            cosine_reg0 <= 36'sb11101010010100011101110110000101;
            sine_reg0   <= 36'sb11111110010100011010001010111010111;
        end
        3798: begin
            cosine_reg0 <= 36'sb11101001100010100001111010001011;
            sine_reg0   <= 36'sb11111110010101001000000110100100010;
        end
        3799: begin
            cosine_reg0 <= 36'sb11101000110000100101110101010001;
            sine_reg0   <= 36'sb11111110010101110101111000011010001;
        end
        3800: begin
            cosine_reg0 <= 36'sb11100111111110101001100111011001;
            sine_reg0   <= 36'sb11111110010110100011100000011100011;
        end
        3801: begin
            cosine_reg0 <= 36'sb11100111001100101101010000100101;
            sine_reg0   <= 36'sb11111110010111010000111110101011001;
        end
        3802: begin
            cosine_reg0 <= 36'sb11100110011010110000110000110110;
            sine_reg0   <= 36'sb11111110010111111110010011000110010;
        end
        3803: begin
            cosine_reg0 <= 36'sb11100101101000110100001000001111;
            sine_reg0   <= 36'sb11111110011000101011011101101101101;
        end
        3804: begin
            cosine_reg0 <= 36'sb11100100110110110111010110110001;
            sine_reg0   <= 36'sb11111110011001011000011110100001100;
        end
        3805: begin
            cosine_reg0 <= 36'sb11100100000100111010011100011110;
            sine_reg0   <= 36'sb11111110011010000101010101100001100;
        end
        3806: begin
            cosine_reg0 <= 36'sb11100011010010111101011001011000;
            sine_reg0   <= 36'sb11111110011010110010000010101101111;
        end
        3807: begin
            cosine_reg0 <= 36'sb11100010100001000000001101100010;
            sine_reg0   <= 36'sb11111110011011011110100110000110100;
        end
        3808: begin
            cosine_reg0 <= 36'sb11100001101111000010111000111101;
            sine_reg0   <= 36'sb11111110011100001010111111101011010;
        end
        3809: begin
            cosine_reg0 <= 36'sb11100000111101000101011011101011;
            sine_reg0   <= 36'sb11111110011100110111001111011100011;
        end
        3810: begin
            cosine_reg0 <= 36'sb11100000001011000111110101101101;
            sine_reg0   <= 36'sb11111110011101100011010101011001100;
        end
        3811: begin
            cosine_reg0 <= 36'sb11011111011001001010000111000111;
            sine_reg0   <= 36'sb11111110011110001111010001100010111;
        end
        3812: begin
            cosine_reg0 <= 36'sb11011110100111001100001111111001;
            sine_reg0   <= 36'sb11111110011110111011000011111000010;
        end
        3813: begin
            cosine_reg0 <= 36'sb11011101110101001110010000000111;
            sine_reg0   <= 36'sb11111110011111100110101100011001110;
        end
        3814: begin
            cosine_reg0 <= 36'sb11011101000011010000000111110000;
            sine_reg0   <= 36'sb11111110100000010010001011000111011;
        end
        3815: begin
            cosine_reg0 <= 36'sb11011100010001010001110110111001;
            sine_reg0   <= 36'sb11111110100000111101100000000001000;
        end
        3816: begin
            cosine_reg0 <= 36'sb11011011011111010011011101100010;
            sine_reg0   <= 36'sb11111110100001101000101011000110101;
        end
        3817: begin
            cosine_reg0 <= 36'sb11011010101101010100111011101101;
            sine_reg0   <= 36'sb11111110100010010011101100011000010;
        end
        3818: begin
            cosine_reg0 <= 36'sb11011001111011010110010001011101;
            sine_reg0   <= 36'sb11111110100010111110100011110101111;
        end
        3819: begin
            cosine_reg0 <= 36'sb11011001001001010111011110110011;
            sine_reg0   <= 36'sb11111110100011101001010001011111011;
        end
        3820: begin
            cosine_reg0 <= 36'sb11011000010111011000100011110001;
            sine_reg0   <= 36'sb11111110100100010011110101010100110;
        end
        3821: begin
            cosine_reg0 <= 36'sb11010111100101011001100000011001;
            sine_reg0   <= 36'sb11111110100100111110001111010110000;
        end
        3822: begin
            cosine_reg0 <= 36'sb11010110110011011010010100101110;
            sine_reg0   <= 36'sb11111110100101101000011111100011001;
        end
        3823: begin
            cosine_reg0 <= 36'sb11010110000001011011000000110000;
            sine_reg0   <= 36'sb11111110100110010010100101111100001;
        end
        3824: begin
            cosine_reg0 <= 36'sb11010101001111011011100100100010;
            sine_reg0   <= 36'sb11111110100110111100100010100001000;
        end
        3825: begin
            cosine_reg0 <= 36'sb11010100011101011100000000000110;
            sine_reg0   <= 36'sb11111110100111100110010101010001100;
        end
        3826: begin
            cosine_reg0 <= 36'sb11010011101011011100010011011110;
            sine_reg0   <= 36'sb11111110101000001111111110001101110;
        end
        3827: begin
            cosine_reg0 <= 36'sb11010010111001011100011110101100;
            sine_reg0   <= 36'sb11111110101000111001011101010101111;
        end
        3828: begin
            cosine_reg0 <= 36'sb11010010000111011100100001110001;
            sine_reg0   <= 36'sb11111110101001100010110010101001101;
        end
        3829: begin
            cosine_reg0 <= 36'sb11010001010101011100011100110000;
            sine_reg0   <= 36'sb11111110101010001011111110001001000;
        end
        3830: begin
            cosine_reg0 <= 36'sb11010000100011011100001111101010;
            sine_reg0   <= 36'sb11111110101010110100111111110100001;
        end
        3831: begin
            cosine_reg0 <= 36'sb11001111110001011011111010100010;
            sine_reg0   <= 36'sb11111110101011011101110111101010110;
        end
        3832: begin
            cosine_reg0 <= 36'sb11001110111111011011011101011001;
            sine_reg0   <= 36'sb11111110101100000110100101101101001;
        end
        3833: begin
            cosine_reg0 <= 36'sb11001110001101011010111000010001;
            sine_reg0   <= 36'sb11111110101100101111001001111011000;
        end
        3834: begin
            cosine_reg0 <= 36'sb11001101011011011010001011001101;
            sine_reg0   <= 36'sb11111110101101010111100100010100100;
        end
        3835: begin
            cosine_reg0 <= 36'sb11001100101001011001010110001110;
            sine_reg0   <= 36'sb11111110101101111111110100111001011;
        end
        3836: begin
            cosine_reg0 <= 36'sb11001011110111011000011001010101;
            sine_reg0   <= 36'sb11111110101110100111111011101001111;
        end
        3837: begin
            cosine_reg0 <= 36'sb11001011000101010111010100100110;
            sine_reg0   <= 36'sb11111110101111001111111000100101111;
        end
        3838: begin
            cosine_reg0 <= 36'sb11001010010011010110001000000010;
            sine_reg0   <= 36'sb11111110101111110111101011101101010;
        end
        3839: begin
            cosine_reg0 <= 36'sb11001001100001010100110011101010;
            sine_reg0   <= 36'sb11111110110000011111010101000000001;
        end
        3840: begin
            cosine_reg0 <= 36'sb11001000101111010011010111100001;
            sine_reg0   <= 36'sb11111110110001000110110100011110011;
        end
        3841: begin
            cosine_reg0 <= 36'sb11000111111101010001110011101001;
            sine_reg0   <= 36'sb11111110110001101110001010001000001;
        end
        3842: begin
            cosine_reg0 <= 36'sb11000111001011010000001000000100;
            sine_reg0   <= 36'sb11111110110010010101010101111101001;
        end
        3843: begin
            cosine_reg0 <= 36'sb11000110011001001110010100110011;
            sine_reg0   <= 36'sb11111110110010111100010111111101100;
        end
        3844: begin
            cosine_reg0 <= 36'sb11000101100111001100011001111000;
            sine_reg0   <= 36'sb11111110110011100011010000001001001;
        end
        3845: begin
            cosine_reg0 <= 36'sb11000100110101001010010111010110;
            sine_reg0   <= 36'sb11111110110100001001111110100000001;
        end
        3846: begin
            cosine_reg0 <= 36'sb11000100000011001000001101001111;
            sine_reg0   <= 36'sb11111110110100110000100011000010011;
        end
        3847: begin
            cosine_reg0 <= 36'sb11000011010001000101111011100011;
            sine_reg0   <= 36'sb11111110110101010110111101101111110;
        end
        3848: begin
            cosine_reg0 <= 36'sb11000010011111000011100010010110;
            sine_reg0   <= 36'sb11111110110101111101001110101000100;
        end
        3849: begin
            cosine_reg0 <= 36'sb11000001101101000001000001101001;
            sine_reg0   <= 36'sb11111110110110100011010101101100011;
        end
        3850: begin
            cosine_reg0 <= 36'sb11000000111010111110011001011110;
            sine_reg0   <= 36'sb11111110110111001001010010111011100;
        end
        3851: begin
            cosine_reg0 <= 36'sb11000000001000111011101001110111;
            sine_reg0   <= 36'sb11111110110111101111000110010101110;
        end
        3852: begin
            cosine_reg0 <= 36'sb10111111010110111000110010110110;
            sine_reg0   <= 36'sb11111110111000010100101111111011001;
        end
        3853: begin
            cosine_reg0 <= 36'sb10111110100100110101110100011100;
            sine_reg0   <= 36'sb11111110111000111010001111101011101;
        end
        3854: begin
            cosine_reg0 <= 36'sb10111101110010110010101110101101;
            sine_reg0   <= 36'sb11111110111001011111100101100111001;
        end
        3855: begin
            cosine_reg0 <= 36'sb10111101000000101111100001101001;
            sine_reg0   <= 36'sb11111110111010000100110001101101110;
        end
        3856: begin
            cosine_reg0 <= 36'sb10111100001110101100001101010011;
            sine_reg0   <= 36'sb11111110111010101001110011111111011;
        end
        3857: begin
            cosine_reg0 <= 36'sb10111011011100101000110001101100;
            sine_reg0   <= 36'sb11111110111011001110101100011100001;
        end
        3858: begin
            cosine_reg0 <= 36'sb10111010101010100101001110110111;
            sine_reg0   <= 36'sb11111110111011110011011011000011110;
        end
        3859: begin
            cosine_reg0 <= 36'sb10111001111000100001100100110101;
            sine_reg0   <= 36'sb11111110111100010111111111110110100;
        end
        3860: begin
            cosine_reg0 <= 36'sb10111001000110011101110011101001;
            sine_reg0   <= 36'sb11111110111100111100011010110100001;
        end
        3861: begin
            cosine_reg0 <= 36'sb10111000010100011001111011010100;
            sine_reg0   <= 36'sb11111110111101100000101011111100101;
        end
        3862: begin
            cosine_reg0 <= 36'sb10110111100010010101111011111000;
            sine_reg0   <= 36'sb11111110111110000100110011010000001;
        end
        3863: begin
            cosine_reg0 <= 36'sb10110110110000010001110101010111;
            sine_reg0   <= 36'sb11111110111110101000110000101110011;
        end
        3864: begin
            cosine_reg0 <= 36'sb10110101111110001101100111110100;
            sine_reg0   <= 36'sb11111110111111001100100100010111101;
        end
        3865: begin
            cosine_reg0 <= 36'sb10110101001100001001010011001111;
            sine_reg0   <= 36'sb11111110111111110000001110001011101;
        end
        3866: begin
            cosine_reg0 <= 36'sb10110100011010000100110111101011;
            sine_reg0   <= 36'sb11111111000000010011101110001010100;
        end
        3867: begin
            cosine_reg0 <= 36'sb10110011101000000000010101001011;
            sine_reg0   <= 36'sb11111111000000110111000100010100001;
        end
        3868: begin
            cosine_reg0 <= 36'sb10110010110101111011101011101110;
            sine_reg0   <= 36'sb11111111000001011010010000101000101;
        end
        3869: begin
            cosine_reg0 <= 36'sb10110010000011110110111011011001;
            sine_reg0   <= 36'sb11111111000001111101010011000111111;
        end
        3870: begin
            cosine_reg0 <= 36'sb10110001010001110010000100001100;
            sine_reg0   <= 36'sb11111111000010100000001011110001110;
        end
        3871: begin
            cosine_reg0 <= 36'sb10110000011111101101000110001010;
            sine_reg0   <= 36'sb11111111000011000010111010100110100;
        end
        3872: begin
            cosine_reg0 <= 36'sb10101111101101101000000001010101;
            sine_reg0   <= 36'sb11111111000011100101011111100101110;
        end
        3873: begin
            cosine_reg0 <= 36'sb10101110111011100010110101101110;
            sine_reg0   <= 36'sb11111111000100000111111010101111111;
        end
        3874: begin
            cosine_reg0 <= 36'sb10101110001001011101100011010111;
            sine_reg0   <= 36'sb11111111000100101010001100000100100;
        end
        3875: begin
            cosine_reg0 <= 36'sb10101101010111011000001010010010;
            sine_reg0   <= 36'sb11111111000101001100010011100011111;
        end
        3876: begin
            cosine_reg0 <= 36'sb10101100100101010010101010100010;
            sine_reg0   <= 36'sb11111111000101101110010001001101110;
        end
        3877: begin
            cosine_reg0 <= 36'sb10101011110011001101000100001000;
            sine_reg0   <= 36'sb11111111000110010000000101000010010;
        end
        3878: begin
            cosine_reg0 <= 36'sb10101011000001000111010111000110;
            sine_reg0   <= 36'sb11111111000110110001101111000001011;
        end
        3879: begin
            cosine_reg0 <= 36'sb10101010001111000001100011011110;
            sine_reg0   <= 36'sb11111111000111010011001111001011000;
        end
        3880: begin
            cosine_reg0 <= 36'sb10101001011100111011101001010010;
            sine_reg0   <= 36'sb11111111000111110100100101011111001;
        end
        3881: begin
            cosine_reg0 <= 36'sb10101000101010110101101000100100;
            sine_reg0   <= 36'sb11111111001000010101110001111101111;
        end
        3882: begin
            cosine_reg0 <= 36'sb10100111111000101111100001010110;
            sine_reg0   <= 36'sb11111111001000110110110100100111000;
        end
        3883: begin
            cosine_reg0 <= 36'sb10100111000110101001010011101010;
            sine_reg0   <= 36'sb11111111001001010111101101011010110;
        end
        3884: begin
            cosine_reg0 <= 36'sb10100110010100100010111111100001;
            sine_reg0   <= 36'sb11111111001001111000011100011000110;
        end
        3885: begin
            cosine_reg0 <= 36'sb10100101100010011100100100111110;
            sine_reg0   <= 36'sb11111111001010011001000001100001011;
        end
        3886: begin
            cosine_reg0 <= 36'sb10100100110000010110000100000010;
            sine_reg0   <= 36'sb11111111001010111001011100110100010;
        end
        3887: begin
            cosine_reg0 <= 36'sb10100011111110001111011100110000;
            sine_reg0   <= 36'sb11111111001011011001101110010001101;
        end
        3888: begin
            cosine_reg0 <= 36'sb10100011001100001000101111001001;
            sine_reg0   <= 36'sb11111111001011111001110101111001011;
        end
        3889: begin
            cosine_reg0 <= 36'sb10100010011010000001111011010000;
            sine_reg0   <= 36'sb11111111001100011001110011101011011;
        end
        3890: begin
            cosine_reg0 <= 36'sb10100001100111111011000001000110;
            sine_reg0   <= 36'sb11111111001100111001100111100111110;
        end
        3891: begin
            cosine_reg0 <= 36'sb10100000110101110100000000101101;
            sine_reg0   <= 36'sb11111111001101011001010001101110100;
        end
        3892: begin
            cosine_reg0 <= 36'sb10100000000011101100111010000111;
            sine_reg0   <= 36'sb11111111001101111000110001111111100;
        end
        3893: begin
            cosine_reg0 <= 36'sb10011111010001100101101101010110;
            sine_reg0   <= 36'sb11111111001110011000001000011010110;
        end
        3894: begin
            cosine_reg0 <= 36'sb10011110011111011110011010011101;
            sine_reg0   <= 36'sb11111111001110110111010101000000011;
        end
        3895: begin
            cosine_reg0 <= 36'sb10011101101101010111000001011100;
            sine_reg0   <= 36'sb11111111001111010110010111110000001;
        end
        3896: begin
            cosine_reg0 <= 36'sb10011100111011001111100010010110;
            sine_reg0   <= 36'sb11111111001111110101010000101010001;
        end
        3897: begin
            cosine_reg0 <= 36'sb10011100001001000111111101001101;
            sine_reg0   <= 36'sb11111111010000010011111111101110011;
        end
        3898: begin
            cosine_reg0 <= 36'sb10011011010111000000010010000011;
            sine_reg0   <= 36'sb11111111010000110010100100111100110;
        end
        3899: begin
            cosine_reg0 <= 36'sb10011010100100111000100000111001;
            sine_reg0   <= 36'sb11111111010001010001000000010101010;
        end
        3900: begin
            cosine_reg0 <= 36'sb10011001110010110000101001110010;
            sine_reg0   <= 36'sb11111111010001101111010001111000000;
        end
        3901: begin
            cosine_reg0 <= 36'sb10011001000000101000101100101111;
            sine_reg0   <= 36'sb11111111010010001101011001100100111;
        end
        3902: begin
            cosine_reg0 <= 36'sb10011000001110100000101001110011;
            sine_reg0   <= 36'sb11111111010010101011010111011011110;
        end
        3903: begin
            cosine_reg0 <= 36'sb10010111011100011000100001000000;
            sine_reg0   <= 36'sb11111111010011001001001011011100110;
        end
        3904: begin
            cosine_reg0 <= 36'sb10010110101010010000010010010110;
            sine_reg0   <= 36'sb11111111010011100110110101100111111;
        end
        3905: begin
            cosine_reg0 <= 36'sb10010101111000000111111101111001;
            sine_reg0   <= 36'sb11111111010100000100010101111101001;
        end
        3906: begin
            cosine_reg0 <= 36'sb10010101000101111111100011101010;
            sine_reg0   <= 36'sb11111111010100100001101100011100010;
        end
        3907: begin
            cosine_reg0 <= 36'sb10010100010011110111000011101100;
            sine_reg0   <= 36'sb11111111010100111110111001000101100;
        end
        3908: begin
            cosine_reg0 <= 36'sb10010011100001101110011101111111;
            sine_reg0   <= 36'sb11111111010101011011111011111000110;
        end
        3909: begin
            cosine_reg0 <= 36'sb10010010101111100101110010100110;
            sine_reg0   <= 36'sb11111111010101111000110100110110000;
        end
        3910: begin
            cosine_reg0 <= 36'sb10010001111101011101000001100011;
            sine_reg0   <= 36'sb11111111010110010101100011111101001;
        end
        3911: begin
            cosine_reg0 <= 36'sb10010001001011010100001010111000;
            sine_reg0   <= 36'sb11111111010110110010001001001110010;
        end
        3912: begin
            cosine_reg0 <= 36'sb10010000011001001011001110100111;
            sine_reg0   <= 36'sb11111111010111001110100100101001011;
        end
        3913: begin
            cosine_reg0 <= 36'sb10001111100111000010001100110010;
            sine_reg0   <= 36'sb11111111010111101010110110001110011;
        end
        3914: begin
            cosine_reg0 <= 36'sb10001110110100111001000101011010;
            sine_reg0   <= 36'sb11111111011000000110111101111101010;
        end
        3915: begin
            cosine_reg0 <= 36'sb10001110000010101111111000100010;
            sine_reg0   <= 36'sb11111111011000100010111011110110000;
        end
        3916: begin
            cosine_reg0 <= 36'sb10001101010000100110100110001011;
            sine_reg0   <= 36'sb11111111011000111110101111111000101;
        end
        3917: begin
            cosine_reg0 <= 36'sb10001100011110011101001110011000;
            sine_reg0   <= 36'sb11111111011001011010011010000101001;
        end
        3918: begin
            cosine_reg0 <= 36'sb10001011101100010011110001001010;
            sine_reg0   <= 36'sb11111111011001110101111010011011100;
        end
        3919: begin
            cosine_reg0 <= 36'sb10001010111010001010001110100100;
            sine_reg0   <= 36'sb11111111011010010001010000111011101;
        end
        3920: begin
            cosine_reg0 <= 36'sb10001010001000000000100110100111;
            sine_reg0   <= 36'sb11111111011010101100011101100101101;
        end
        3921: begin
            cosine_reg0 <= 36'sb10001001010101110110111001010101;
            sine_reg0   <= 36'sb11111111011011000111100000011001010;
        end
        3922: begin
            cosine_reg0 <= 36'sb10001000100011101101000110110000;
            sine_reg0   <= 36'sb11111111011011100010011001010110110;
        end
        3923: begin
            cosine_reg0 <= 36'sb10000111110001100011001110111010;
            sine_reg0   <= 36'sb11111111011011111101001000011110000;
        end
        3924: begin
            cosine_reg0 <= 36'sb10000110111111011001010001110101;
            sine_reg0   <= 36'sb11111111011100010111101101101111000;
        end
        3925: begin
            cosine_reg0 <= 36'sb10000110001101001111001111100011;
            sine_reg0   <= 36'sb11111111011100110010001001001001110;
        end
        3926: begin
            cosine_reg0 <= 36'sb10000101011011000101001000000110;
            sine_reg0   <= 36'sb11111111011101001100011010101110001;
        end
        3927: begin
            cosine_reg0 <= 36'sb10000100101000111010111011100000;
            sine_reg0   <= 36'sb11111111011101100110100010011100010;
        end
        3928: begin
            cosine_reg0 <= 36'sb10000011110110110000101001110010;
            sine_reg0   <= 36'sb11111111011110000000100000010100000;
        end
        3929: begin
            cosine_reg0 <= 36'sb10000011000100100110010010111111;
            sine_reg0   <= 36'sb11111111011110011010010100010101011;
        end
        3930: begin
            cosine_reg0 <= 36'sb10000010010010011011110111001001;
            sine_reg0   <= 36'sb11111111011110110011111110100000011;
        end
        3931: begin
            cosine_reg0 <= 36'sb10000001100000010001010110010001;
            sine_reg0   <= 36'sb11111111011111001101011110110101001;
        end
        3932: begin
            cosine_reg0 <= 36'sb10000000101110000110110000011010;
            sine_reg0   <= 36'sb11111111011111100110110101010011011;
        end
        3933: begin
            cosine_reg0 <= 36'sb1111111111011111100000101100101;
            sine_reg0   <= 36'sb11111111100000000000000001111011010;
        end
        3934: begin
            cosine_reg0 <= 36'sb1111111001001110001010101110100;
            sine_reg0   <= 36'sb11111111100000011001000100101100110;
        end
        3935: begin
            cosine_reg0 <= 36'sb1111110010111100110100001001010;
            sine_reg0   <= 36'sb11111111100000110001111101100111110;
        end
        3936: begin
            cosine_reg0 <= 36'sb1111101100101011011100111101000;
            sine_reg0   <= 36'sb11111111100001001010101100101100011;
        end
        3937: begin
            cosine_reg0 <= 36'sb1111100110011010000101001010000;
            sine_reg0   <= 36'sb11111111100001100011010001111010011;
        end
        3938: begin
            cosine_reg0 <= 36'sb1111100000001000101100110000100;
            sine_reg0   <= 36'sb11111111100001111011101101010010000;
        end
        3939: begin
            cosine_reg0 <= 36'sb1111011001110111010011110000110;
            sine_reg0   <= 36'sb11111111100010010011111110110011010;
        end
        3940: begin
            cosine_reg0 <= 36'sb1111010011100101111010001011000;
            sine_reg0   <= 36'sb11111111100010101100000110011101111;
        end
        3941: begin
            cosine_reg0 <= 36'sb1111001101010100011111111111100;
            sine_reg0   <= 36'sb11111111100011000100000100010001111;
        end
        3942: begin
            cosine_reg0 <= 36'sb1111000111000011000101001110011;
            sine_reg0   <= 36'sb11111111100011011011111000001111100;
        end
        3943: begin
            cosine_reg0 <= 36'sb1111000000110001101001111000001;
            sine_reg0   <= 36'sb11111111100011110011100010010110100;
        end
        3944: begin
            cosine_reg0 <= 36'sb1110111010100000001101111100110;
            sine_reg0   <= 36'sb11111111100100001011000010100110111;
        end
        3945: begin
            cosine_reg0 <= 36'sb1110110100001110110001011100101;
            sine_reg0   <= 36'sb11111111100100100010011001000000110;
        end
        3946: begin
            cosine_reg0 <= 36'sb1110101101111101010100010111111;
            sine_reg0   <= 36'sb11111111100100111001100101100100000;
        end
        3947: begin
            cosine_reg0 <= 36'sb1110100111101011110110101110111;
            sine_reg0   <= 36'sb11111111100101010000101000010000101;
        end
        3948: begin
            cosine_reg0 <= 36'sb1110100001011010011000100001110;
            sine_reg0   <= 36'sb11111111100101100111100001000110110;
        end
        3949: begin
            cosine_reg0 <= 36'sb1110011011001000111001110000110;
            sine_reg0   <= 36'sb11111111100101111110010000000110001;
        end
        3950: begin
            cosine_reg0 <= 36'sb1110010100110111011010011100010;
            sine_reg0   <= 36'sb11111111100110010100110101001110111;
        end
        3951: begin
            cosine_reg0 <= 36'sb1110001110100101111010100100011;
            sine_reg0   <= 36'sb11111111100110101011010000100000111;
        end
        3952: begin
            cosine_reg0 <= 36'sb1110001000010100011010001001011;
            sine_reg0   <= 36'sb11111111100111000001100001111100010;
        end
        3953: begin
            cosine_reg0 <= 36'sb1110000010000010111001001011100;
            sine_reg0   <= 36'sb11111111100111010111101001100001000;
        end
        3954: begin
            cosine_reg0 <= 36'sb1101111011110001010111101011000;
            sine_reg0   <= 36'sb11111111100111101101100111001111000;
        end
        3955: begin
            cosine_reg0 <= 36'sb1101110101011111110101101000010;
            sine_reg0   <= 36'sb11111111101000000011011011000110010;
        end
        3956: begin
            cosine_reg0 <= 36'sb1101101111001110010011000011010;
            sine_reg0   <= 36'sb11111111101000011001000101000110111;
        end
        3957: begin
            cosine_reg0 <= 36'sb1101101000111100101111111100010;
            sine_reg0   <= 36'sb11111111101000101110100101010000101;
        end
        3958: begin
            cosine_reg0 <= 36'sb1101100010101011001100010011110;
            sine_reg0   <= 36'sb11111111101001000011111011100011101;
        end
        3959: begin
            cosine_reg0 <= 36'sb1101011100011001101000001001110;
            sine_reg0   <= 36'sb11111111101001011001001000000000000;
        end
        3960: begin
            cosine_reg0 <= 36'sb1101010110001000000011011110101;
            sine_reg0   <= 36'sb11111111101001101110001010100101011;
        end
        3961: begin
            cosine_reg0 <= 36'sb1101001111110110011110010010101;
            sine_reg0   <= 36'sb11111111101010000011000011010100001;
        end
        3962: begin
            cosine_reg0 <= 36'sb1101001001100100111000100101111;
            sine_reg0   <= 36'sb11111111101010010111110010001100000;
        end
        3963: begin
            cosine_reg0 <= 36'sb1101000011010011010010011000101;
            sine_reg0   <= 36'sb11111111101010101100010111001101001;
        end
        3964: begin
            cosine_reg0 <= 36'sb1100111101000001101011101011010;
            sine_reg0   <= 36'sb11111111101011000000110010010111011;
        end
        3965: begin
            cosine_reg0 <= 36'sb1100110110110000000100011101111;
            sine_reg0   <= 36'sb11111111101011010101000011101010110;
        end
        3966: begin
            cosine_reg0 <= 36'sb1100110000011110011100110000111;
            sine_reg0   <= 36'sb11111111101011101001001011000111010;
        end
        3967: begin
            cosine_reg0 <= 36'sb1100101010001100110100100100010;
            sine_reg0   <= 36'sb11111111101011111101001000101100111;
        end
        3968: begin
            cosine_reg0 <= 36'sb1100100011111011001011111000100;
            sine_reg0   <= 36'sb11111111101100010000111100011011101;
        end
        3969: begin
            cosine_reg0 <= 36'sb1100011101101001100010101101110;
            sine_reg0   <= 36'sb11111111101100100100100110010011100;
        end
        3970: begin
            cosine_reg0 <= 36'sb1100010111010111111001000100010;
            sine_reg0   <= 36'sb11111111101100111000000110010100100;
        end
        3971: begin
            cosine_reg0 <= 36'sb1100010001000110001110111100001;
            sine_reg0   <= 36'sb11111111101101001011011100011110101;
        end
        3972: begin
            cosine_reg0 <= 36'sb1100001010110100100100010101111;
            sine_reg0   <= 36'sb11111111101101011110101000110001110;
        end
        3973: begin
            cosine_reg0 <= 36'sb1100000100100010111001010001100;
            sine_reg0   <= 36'sb11111111101101110001101011001101111;
        end
        3974: begin
            cosine_reg0 <= 36'sb1011111110010001001101101111011;
            sine_reg0   <= 36'sb11111111101110000100100011110011001;
        end
        3975: begin
            cosine_reg0 <= 36'sb1011110111111111100001101111110;
            sine_reg0   <= 36'sb11111111101110010111010010100001011;
        end
        3976: begin
            cosine_reg0 <= 36'sb1011110001101101110101010010110;
            sine_reg0   <= 36'sb11111111101110101001110111011000110;
        end
        3977: begin
            cosine_reg0 <= 36'sb1011101011011100001000011000110;
            sine_reg0   <= 36'sb11111111101110111100010010011001000;
        end
        3978: begin
            cosine_reg0 <= 36'sb1011100101001010011011000001111;
            sine_reg0   <= 36'sb11111111101111001110100011100010011;
        end
        3979: begin
            cosine_reg0 <= 36'sb1011011110111000101101001110100;
            sine_reg0   <= 36'sb11111111101111100000101010110100101;
        end
        3980: begin
            cosine_reg0 <= 36'sb1011011000100110111110111110110;
            sine_reg0   <= 36'sb11111111101111110010101000010000000;
        end
        3981: begin
            cosine_reg0 <= 36'sb1011010010010101010000010010111;
            sine_reg0   <= 36'sb11111111110000000100011011110100010;
        end
        3982: begin
            cosine_reg0 <= 36'sb1011001100000011100001001011010;
            sine_reg0   <= 36'sb11111111110000010110000101100001100;
        end
        3983: begin
            cosine_reg0 <= 36'sb1011000101110001110001100111111;
            sine_reg0   <= 36'sb11111111110000100111100101010111101;
        end
        3984: begin
            cosine_reg0 <= 36'sb1010111111100000000001101001010;
            sine_reg0   <= 36'sb11111111110000111000111011010110110;
        end
        3985: begin
            cosine_reg0 <= 36'sb1010111001001110010001001111100;
            sine_reg0   <= 36'sb11111111110001001010000111011110110;
        end
        3986: begin
            cosine_reg0 <= 36'sb1010110010111100100000011010111;
            sine_reg0   <= 36'sb11111111110001011011001001101111110;
        end
        3987: begin
            cosine_reg0 <= 36'sb1010101100101010101111001011100;
            sine_reg0   <= 36'sb11111111110001101100000010001001101;
        end
        3988: begin
            cosine_reg0 <= 36'sb1010100110011000111101100001111;
            sine_reg0   <= 36'sb11111111110001111100110000101100011;
        end
        3989: begin
            cosine_reg0 <= 36'sb1010100000000111001011011110000;
            sine_reg0   <= 36'sb11111111110010001101010101011000000;
        end
        3990: begin
            cosine_reg0 <= 36'sb1010011001110101011001000000010;
            sine_reg0   <= 36'sb11111111110010011101110000001100100;
        end
        3991: begin
            cosine_reg0 <= 36'sb1010010011100011100110001000111;
            sine_reg0   <= 36'sb11111111110010101110000001001001111;
        end
        3992: begin
            cosine_reg0 <= 36'sb1010001101010001110010111000000;
            sine_reg0   <= 36'sb11111111110010111110001000010000001;
        end
        3993: begin
            cosine_reg0 <= 36'sb1010000110111111111111001110000;
            sine_reg0   <= 36'sb11111111110011001110000101011111010;
        end
        3994: begin
            cosine_reg0 <= 36'sb1010000000101110001011001011000;
            sine_reg0   <= 36'sb11111111110011011101111000110111001;
        end
        3995: begin
            cosine_reg0 <= 36'sb1001111010011100010110101111010;
            sine_reg0   <= 36'sb11111111110011101101100010010111111;
        end
        3996: begin
            cosine_reg0 <= 36'sb1001110100001010100001111011001;
            sine_reg0   <= 36'sb11111111110011111101000010000001100;
        end
        3997: begin
            cosine_reg0 <= 36'sb1001101101111000101100101110110;
            sine_reg0   <= 36'sb11111111110100001100010111110011111;
        end
        3998: begin
            cosine_reg0 <= 36'sb1001100111100110110111001010011;
            sine_reg0   <= 36'sb11111111110100011011100011101111001;
        end
        3999: begin
            cosine_reg0 <= 36'sb1001100001010101000001001110011;
            sine_reg0   <= 36'sb11111111110100101010100101110011001;
        end
        4000: begin
            cosine_reg0 <= 36'sb1001011011000011001010111010110;
            sine_reg0   <= 36'sb11111111110100111001011101111111111;
        end
        4001: begin
            cosine_reg0 <= 36'sb1001010100110001010100010000000;
            sine_reg0   <= 36'sb11111111110101001000001100010101011;
        end
        4002: begin
            cosine_reg0 <= 36'sb1001001110011111011101001110001;
            sine_reg0   <= 36'sb11111111110101010110110000110011101;
        end
        4003: begin
            cosine_reg0 <= 36'sb1001001000001101100101110101101;
            sine_reg0   <= 36'sb11111111110101100101001011011010110;
        end
        4004: begin
            cosine_reg0 <= 36'sb1001000001111011101110000110100;
            sine_reg0   <= 36'sb11111111110101110011011100001010100;
        end
        4005: begin
            cosine_reg0 <= 36'sb1000111011101001110110000001001;
            sine_reg0   <= 36'sb11111111110110000001100011000011001;
        end
        4006: begin
            cosine_reg0 <= 36'sb1000110101010111111101100101101;
            sine_reg0   <= 36'sb11111111110110001111100000000100011;
        end
        4007: begin
            cosine_reg0 <= 36'sb1000101111000110000100110100011;
            sine_reg0   <= 36'sb11111111110110011101010011001110011;
        end
        4008: begin
            cosine_reg0 <= 36'sb1000101000110100001011101101101;
            sine_reg0   <= 36'sb11111111110110101010111100100001000;
        end
        4009: begin
            cosine_reg0 <= 36'sb1000100010100010010010010001100;
            sine_reg0   <= 36'sb11111111110110111000011011111100100;
        end
        4010: begin
            cosine_reg0 <= 36'sb1000011100010000011000100000011;
            sine_reg0   <= 36'sb11111111110111000101110001100000101;
        end
        4011: begin
            cosine_reg0 <= 36'sb1000010101111110011110011010011;
            sine_reg0   <= 36'sb11111111110111010010111101001101011;
        end
        4012: begin
            cosine_reg0 <= 36'sb1000001111101100100011111111110;
            sine_reg0   <= 36'sb11111111110111011111111111000010111;
        end
        4013: begin
            cosine_reg0 <= 36'sb1000001001011010101001010000111;
            sine_reg0   <= 36'sb11111111110111101100110111000001000;
        end
        4014: begin
            cosine_reg0 <= 36'sb1000000011001000101110001101111;
            sine_reg0   <= 36'sb11111111110111111001100101000111111;
        end
        4015: begin
            cosine_reg0 <= 36'sb111111100110110110010110111000;
            sine_reg0   <= 36'sb11111111111000000110001001010111010;
        end
        4016: begin
            cosine_reg0 <= 36'sb111110110100100110111001100100;
            sine_reg0   <= 36'sb11111111111000010010100011101111011;
        end
        4017: begin
            cosine_reg0 <= 36'sb111110000010010111011001110101;
            sine_reg0   <= 36'sb11111111111000011110110100010000010;
        end
        4018: begin
            cosine_reg0 <= 36'sb111101010000000111110111101100;
            sine_reg0   <= 36'sb11111111111000101010111010111001101;
        end
        4019: begin
            cosine_reg0 <= 36'sb111100011101111000010011001101;
            sine_reg0   <= 36'sb11111111111000110110110111101011101;
        end
        4020: begin
            cosine_reg0 <= 36'sb111011101011101000101100011001;
            sine_reg0   <= 36'sb11111111111001000010101010100110010;
        end
        4021: begin
            cosine_reg0 <= 36'sb111010111001011001000011010001;
            sine_reg0   <= 36'sb11111111111001001110010011101001100;
        end
        4022: begin
            cosine_reg0 <= 36'sb111010000111001001010111111000;
            sine_reg0   <= 36'sb11111111111001011001110010110101011;
        end
        4023: begin
            cosine_reg0 <= 36'sb111001010100111001101010010000;
            sine_reg0   <= 36'sb11111111111001100101001000001001111;
        end
        4024: begin
            cosine_reg0 <= 36'sb111000100010101001111010011010;
            sine_reg0   <= 36'sb11111111111001110000010011100111000;
        end
        4025: begin
            cosine_reg0 <= 36'sb110111110000011010001000011000;
            sine_reg0   <= 36'sb11111111111001111011010101001100101;
        end
        4026: begin
            cosine_reg0 <= 36'sb110110111110001010010100001101;
            sine_reg0   <= 36'sb11111111111010000110001100111010111;
        end
        4027: begin
            cosine_reg0 <= 36'sb110110001011111010011101111011;
            sine_reg0   <= 36'sb11111111111010010000111010110001101;
        end
        4028: begin
            cosine_reg0 <= 36'sb110101011001101010100101100011;
            sine_reg0   <= 36'sb11111111111010011011011110110001000;
        end
        4029: begin
            cosine_reg0 <= 36'sb110100100111011010101011000111;
            sine_reg0   <= 36'sb11111111111010100101111000111001000;
        end
        4030: begin
            cosine_reg0 <= 36'sb110011110101001010101110101001;
            sine_reg0   <= 36'sb11111111111010110000001001001001011;
        end
        4031: begin
            cosine_reg0 <= 36'sb110011000010111010110000001011;
            sine_reg0   <= 36'sb11111111111010111010001111100010100;
        end
        4032: begin
            cosine_reg0 <= 36'sb110010010000101010101111101111;
            sine_reg0   <= 36'sb11111111111011000100001100000100000;
        end
        4033: begin
            cosine_reg0 <= 36'sb110001011110011010101101011000;
            sine_reg0   <= 36'sb11111111111011001101111110101110001;
        end
        4034: begin
            cosine_reg0 <= 36'sb110000101100001010101001000110;
            sine_reg0   <= 36'sb11111111111011010111100111100000110;
        end
        4035: begin
            cosine_reg0 <= 36'sb101111111001111010100010111100;
            sine_reg0   <= 36'sb11111111111011100001000110011011111;
        end
        4036: begin
            cosine_reg0 <= 36'sb101111000111101010011010111100;
            sine_reg0   <= 36'sb11111111111011101010011011011111101;
        end
        4037: begin
            cosine_reg0 <= 36'sb101110010101011010010001000111;
            sine_reg0   <= 36'sb11111111111011110011100110101011110;
        end
        4038: begin
            cosine_reg0 <= 36'sb101101100011001010000101100001;
            sine_reg0   <= 36'sb11111111111011111100101000000000100;
        end
        4039: begin
            cosine_reg0 <= 36'sb101100110000111001111000001001;
            sine_reg0   <= 36'sb11111111111100000101011111011101110;
        end
        4040: begin
            cosine_reg0 <= 36'sb101011111110101001101001000100;
            sine_reg0   <= 36'sb11111111111100001110001101000011011;
        end
        4041: begin
            cosine_reg0 <= 36'sb101011001100011001011000010010;
            sine_reg0   <= 36'sb11111111111100010110110000110001101;
        end
        4042: begin
            cosine_reg0 <= 36'sb101010011010001001000101110101;
            sine_reg0   <= 36'sb11111111111100011111001010101000010;
        end
        4043: begin
            cosine_reg0 <= 36'sb101001100111111000110001110000;
            sine_reg0   <= 36'sb11111111111100100111011010100111011;
        end
        4044: begin
            cosine_reg0 <= 36'sb101000110101101000011100000100;
            sine_reg0   <= 36'sb11111111111100101111100000101111000;
        end
        4045: begin
            cosine_reg0 <= 36'sb101000000011011000000100110011;
            sine_reg0   <= 36'sb11111111111100110111011100111111001;
        end
        4046: begin
            cosine_reg0 <= 36'sb100111010001000111101100000000;
            sine_reg0   <= 36'sb11111111111100111111001111010111110;
        end
        4047: begin
            cosine_reg0 <= 36'sb100110011110110111010001101011;
            sine_reg0   <= 36'sb11111111111101000110110111111000110;
        end
        4048: begin
            cosine_reg0 <= 36'sb100101101100100110110101111000;
            sine_reg0   <= 36'sb11111111111101001110010110100010010;
        end
        4049: begin
            cosine_reg0 <= 36'sb100100111010010110011000100111;
            sine_reg0   <= 36'sb11111111111101010101101011010100001;
        end
        4050: begin
            cosine_reg0 <= 36'sb100100001000000101111001111100;
            sine_reg0   <= 36'sb11111111111101011100110110001110100;
        end
        4051: begin
            cosine_reg0 <= 36'sb100011010101110101011001110111;
            sine_reg0   <= 36'sb11111111111101100011110111010001011;
        end
        4052: begin
            cosine_reg0 <= 36'sb100010100011100100111000011011;
            sine_reg0   <= 36'sb11111111111101101010101110011100101;
        end
        4053: begin
            cosine_reg0 <= 36'sb100001110001010100010101101010;
            sine_reg0   <= 36'sb11111111111101110001011011110000011;
        end
        4054: begin
            cosine_reg0 <= 36'sb100000111111000011110001100110;
            sine_reg0   <= 36'sb11111111111101110111111111001100100;
        end
        4055: begin
            cosine_reg0 <= 36'sb100000001100110011001100010000;
            sine_reg0   <= 36'sb11111111111101111110011000110001000;
        end
        4056: begin
            cosine_reg0 <= 36'sb11111011010100010100101101011;
            sine_reg0   <= 36'sb11111111111110000100101000011110000;
        end
        4057: begin
            cosine_reg0 <= 36'sb11110101000010001111101111000;
            sine_reg0   <= 36'sb11111111111110001010101110010011100;
        end
        4058: begin
            cosine_reg0 <= 36'sb11101110110000001010100111010;
            sine_reg0   <= 36'sb11111111111110010000101010010001010;
        end
        4059: begin
            cosine_reg0 <= 36'sb11101000011110000101010110010;
            sine_reg0   <= 36'sb11111111111110010110011100010111100;
        end
        4060: begin
            cosine_reg0 <= 36'sb11100010001011111111111100010;
            sine_reg0   <= 36'sb11111111111110011100000100100110001;
        end
        4061: begin
            cosine_reg0 <= 36'sb11011011111001111010011001100;
            sine_reg0   <= 36'sb11111111111110100001100010111101010;
        end
        4062: begin
            cosine_reg0 <= 36'sb11010101100111110100101110011;
            sine_reg0   <= 36'sb11111111111110100110110111011100101;
        end
        4063: begin
            cosine_reg0 <= 36'sb11001111010101101110111011000;
            sine_reg0   <= 36'sb11111111111110101100000010000100100;
        end
        4064: begin
            cosine_reg0 <= 36'sb11001001000011101000111111101;
            sine_reg0   <= 36'sb11111111111110110001000010110100110;
        end
        4065: begin
            cosine_reg0 <= 36'sb11000010110001100010111100100;
            sine_reg0   <= 36'sb11111111111110110101111001101101011;
        end
        4066: begin
            cosine_reg0 <= 36'sb10111100011111011100110001111;
            sine_reg0   <= 36'sb11111111111110111010100110101110011;
        end
        4067: begin
            cosine_reg0 <= 36'sb10110110001101010110011111111;
            sine_reg0   <= 36'sb11111111111110111111001001110111111;
        end
        4068: begin
            cosine_reg0 <= 36'sb10101111111011010000000111000;
            sine_reg0   <= 36'sb11111111111111000011100011001001101;
        end
        4069: begin
            cosine_reg0 <= 36'sb10101001101001001001100111010;
            sine_reg0   <= 36'sb11111111111111000111110010100011110;
        end
        4070: begin
            cosine_reg0 <= 36'sb10100011010111000011000001000;
            sine_reg0   <= 36'sb11111111111111001011111000000110011;
        end
        4071: begin
            cosine_reg0 <= 36'sb10011101000100111100010100011;
            sine_reg0   <= 36'sb11111111111111001111110011110001010;
        end
        4072: begin
            cosine_reg0 <= 36'sb10010110110010110101100001110;
            sine_reg0   <= 36'sb11111111111111010011100101100100101;
        end
        4073: begin
            cosine_reg0 <= 36'sb10010000100000101110101001011;
            sine_reg0   <= 36'sb11111111111111010111001101100000010;
        end
        4074: begin
            cosine_reg0 <= 36'sb10001010001110100111101011011;
            sine_reg0   <= 36'sb11111111111111011010101011100100011;
        end
        4075: begin
            cosine_reg0 <= 36'sb10000011111100100000101000000;
            sine_reg0   <= 36'sb11111111111111011101111111110000110;
        end
        4076: begin
            cosine_reg0 <= 36'sb1111101101010011001011111101;
            sine_reg0   <= 36'sb11111111111111100001001010000101100;
        end
        4077: begin
            cosine_reg0 <= 36'sb1110111011000010010010010011;
            sine_reg0   <= 36'sb11111111111111100100001010100010110;
        end
        4078: begin
            cosine_reg0 <= 36'sb1110001000110001011000000100;
            sine_reg0   <= 36'sb11111111111111100111000001001000010;
        end
        4079: begin
            cosine_reg0 <= 36'sb1101010110100000011101010010;
            sine_reg0   <= 36'sb11111111111111101001101101110110001;
        end
        4080: begin
            cosine_reg0 <= 36'sb1100100100001111100001111111;
            sine_reg0   <= 36'sb11111111111111101100010000101100011;
        end
        4081: begin
            cosine_reg0 <= 36'sb1011110001111110100110001101;
            sine_reg0   <= 36'sb11111111111111101110101001101010111;
        end
        4082: begin
            cosine_reg0 <= 36'sb1010111111101101101001111111;
            sine_reg0   <= 36'sb11111111111111110000111000110001111;
        end
        4083: begin
            cosine_reg0 <= 36'sb1010001101011100101101010101;
            sine_reg0   <= 36'sb11111111111111110010111110000001001;
        end
        4084: begin
            cosine_reg0 <= 36'sb1001011011001011110000010001;
            sine_reg0   <= 36'sb11111111111111110100111001011000111;
        end
        4085: begin
            cosine_reg0 <= 36'sb1000101000111010110010110111;
            sine_reg0   <= 36'sb11111111111111110110101010111000111;
        end
        4086: begin
            cosine_reg0 <= 36'sb111110110101001110101000111;
            sine_reg0   <= 36'sb11111111111111111000010010100001001;
        end
        4087: begin
            cosine_reg0 <= 36'sb111000100011000110111000100;
            sine_reg0   <= 36'sb11111111111111111001110000010001111;
        end
        4088: begin
            cosine_reg0 <= 36'sb110010010000111111000110000;
            sine_reg0   <= 36'sb11111111111111111011000100001011000;
        end
        4089: begin
            cosine_reg0 <= 36'sb101011111110110111010001100;
            sine_reg0   <= 36'sb11111111111111111100001110001100011;
        end
        4090: begin
            cosine_reg0 <= 36'sb100101101100101111011011010;
            sine_reg0   <= 36'sb11111111111111111101001110010110001;
        end
        4091: begin
            cosine_reg0 <= 36'sb11111011010100111100011101;
            sine_reg0   <= 36'sb11111111111111111110000100101000010;
        end
        4092: begin
            cosine_reg0 <= 36'sb11001001000011111101010110;
            sine_reg0   <= 36'sb11111111111111111110110001000010101;
        end
        4093: begin
            cosine_reg0 <= 36'sb10010110110010111110000111;
            sine_reg0   <= 36'sb11111111111111111111010011100101011;
        end
        4094: begin
            cosine_reg0 <= 36'sb1100100100001111110110011;
            sine_reg0   <= 36'sb11111111111111111111101100010000101;
        end
        4095: begin
            cosine_reg0 <= 36'sb110010010000111111011010;
            sine_reg0   <= 36'sb11111111111111111111111011000100000;
        end
        4096: begin
            cosine_reg0 <= 36'sb0;
            sine_reg0   <= 36'sb11111111111111111111111111111111111;
        end
        4097: begin
            cosine_reg0 <= 36'sb111111111111001101101111000000100110;
            sine_reg0   <= 36'sb11111111111111111111111011000100000;
        end
        4098: begin
            cosine_reg0 <= 36'sb111111111110011011011110000001001101;
            sine_reg0   <= 36'sb11111111111111111111101100010000101;
        end
        4099: begin
            cosine_reg0 <= 36'sb111111111101101001001101000001111001;
            sine_reg0   <= 36'sb11111111111111111111010011100101011;
        end
        4100: begin
            cosine_reg0 <= 36'sb111111111100110110111100000010101010;
            sine_reg0   <= 36'sb11111111111111111110110001000010101;
        end
        4101: begin
            cosine_reg0 <= 36'sb111111111100000100101011000011100011;
            sine_reg0   <= 36'sb11111111111111111110000100101000010;
        end
        4102: begin
            cosine_reg0 <= 36'sb111111111011010010011010000100100110;
            sine_reg0   <= 36'sb11111111111111111101001110010110001;
        end
        4103: begin
            cosine_reg0 <= 36'sb111111111010100000001001000101110100;
            sine_reg0   <= 36'sb11111111111111111100001110001100011;
        end
        4104: begin
            cosine_reg0 <= 36'sb111111111001101101111000000111010000;
            sine_reg0   <= 36'sb11111111111111111011000100001011000;
        end
        4105: begin
            cosine_reg0 <= 36'sb111111111000111011100111001000111100;
            sine_reg0   <= 36'sb11111111111111111001110000010001111;
        end
        4106: begin
            cosine_reg0 <= 36'sb111111111000001001010110001010111001;
            sine_reg0   <= 36'sb11111111111111111000010010100001001;
        end
        4107: begin
            cosine_reg0 <= 36'sb111111110111010111000101001101001001;
            sine_reg0   <= 36'sb11111111111111110110101010111000111;
        end
        4108: begin
            cosine_reg0 <= 36'sb111111110110100100110100001111101111;
            sine_reg0   <= 36'sb11111111111111110100111001011000111;
        end
        4109: begin
            cosine_reg0 <= 36'sb111111110101110010100011010010101011;
            sine_reg0   <= 36'sb11111111111111110010111110000001001;
        end
        4110: begin
            cosine_reg0 <= 36'sb111111110101000000010010010110000001;
            sine_reg0   <= 36'sb11111111111111110000111000110001111;
        end
        4111: begin
            cosine_reg0 <= 36'sb111111110100001110000001011001110011;
            sine_reg0   <= 36'sb11111111111111101110101001101010111;
        end
        4112: begin
            cosine_reg0 <= 36'sb111111110011011011110000011110000001;
            sine_reg0   <= 36'sb11111111111111101100010000101100011;
        end
        4113: begin
            cosine_reg0 <= 36'sb111111110010101001011111100010101110;
            sine_reg0   <= 36'sb11111111111111101001101101110110001;
        end
        4114: begin
            cosine_reg0 <= 36'sb111111110001110111001110100111111100;
            sine_reg0   <= 36'sb11111111111111100111000001001000010;
        end
        4115: begin
            cosine_reg0 <= 36'sb111111110001000100111101101101101101;
            sine_reg0   <= 36'sb11111111111111100100001010100010110;
        end
        4116: begin
            cosine_reg0 <= 36'sb111111110000010010101100110100000011;
            sine_reg0   <= 36'sb11111111111111100001001010000101100;
        end
        4117: begin
            cosine_reg0 <= 36'sb111111101111100000011011111011000000;
            sine_reg0   <= 36'sb11111111111111011101111111110000110;
        end
        4118: begin
            cosine_reg0 <= 36'sb111111101110101110001011000010100101;
            sine_reg0   <= 36'sb11111111111111011010101011100100011;
        end
        4119: begin
            cosine_reg0 <= 36'sb111111101101111011111010001010110101;
            sine_reg0   <= 36'sb11111111111111010111001101100000010;
        end
        4120: begin
            cosine_reg0 <= 36'sb111111101101001001101001010011110010;
            sine_reg0   <= 36'sb11111111111111010011100101100100101;
        end
        4121: begin
            cosine_reg0 <= 36'sb111111101100010111011000011101011101;
            sine_reg0   <= 36'sb11111111111111001111110011110001010;
        end
        4122: begin
            cosine_reg0 <= 36'sb111111101011100101000111100111111000;
            sine_reg0   <= 36'sb11111111111111001011111000000110011;
        end
        4123: begin
            cosine_reg0 <= 36'sb111111101010110010110110110011000110;
            sine_reg0   <= 36'sb11111111111111000111110010100011110;
        end
        4124: begin
            cosine_reg0 <= 36'sb111111101010000000100101111111001000;
            sine_reg0   <= 36'sb11111111111111000011100011001001101;
        end
        4125: begin
            cosine_reg0 <= 36'sb111111101001001110010101001100000001;
            sine_reg0   <= 36'sb11111111111110111111001001110111111;
        end
        4126: begin
            cosine_reg0 <= 36'sb111111101000011100000100011001110001;
            sine_reg0   <= 36'sb11111111111110111010100110101110011;
        end
        4127: begin
            cosine_reg0 <= 36'sb111111100111101001110011101000011100;
            sine_reg0   <= 36'sb11111111111110110101111001101101011;
        end
        4128: begin
            cosine_reg0 <= 36'sb111111100110110111100010111000000011;
            sine_reg0   <= 36'sb11111111111110110001000010110100110;
        end
        4129: begin
            cosine_reg0 <= 36'sb111111100110000101010010001000101000;
            sine_reg0   <= 36'sb11111111111110101100000010000100100;
        end
        4130: begin
            cosine_reg0 <= 36'sb111111100101010011000001011010001101;
            sine_reg0   <= 36'sb11111111111110100110110111011100101;
        end
        4131: begin
            cosine_reg0 <= 36'sb111111100100100000110000101100110100;
            sine_reg0   <= 36'sb11111111111110100001100010111101010;
        end
        4132: begin
            cosine_reg0 <= 36'sb111111100011101110100000000000011110;
            sine_reg0   <= 36'sb11111111111110011100000100100110001;
        end
        4133: begin
            cosine_reg0 <= 36'sb111111100010111100001111010101001110;
            sine_reg0   <= 36'sb11111111111110010110011100010111100;
        end
        4134: begin
            cosine_reg0 <= 36'sb111111100010001001111110101011000110;
            sine_reg0   <= 36'sb11111111111110010000101010010001010;
        end
        4135: begin
            cosine_reg0 <= 36'sb111111100001010111101110000010001000;
            sine_reg0   <= 36'sb11111111111110001010101110010011100;
        end
        4136: begin
            cosine_reg0 <= 36'sb111111100000100101011101011010010101;
            sine_reg0   <= 36'sb11111111111110000100101000011110000;
        end
        4137: begin
            cosine_reg0 <= 36'sb111111011111110011001100110011110000;
            sine_reg0   <= 36'sb11111111111101111110011000110001000;
        end
        4138: begin
            cosine_reg0 <= 36'sb111111011111000000111100001110011010;
            sine_reg0   <= 36'sb11111111111101110111111111001100100;
        end
        4139: begin
            cosine_reg0 <= 36'sb111111011110001110101011101010010110;
            sine_reg0   <= 36'sb11111111111101110001011011110000011;
        end
        4140: begin
            cosine_reg0 <= 36'sb111111011101011100011011000111100101;
            sine_reg0   <= 36'sb11111111111101101010101110011100101;
        end
        4141: begin
            cosine_reg0 <= 36'sb111111011100101010001010100110001001;
            sine_reg0   <= 36'sb11111111111101100011110111010001011;
        end
        4142: begin
            cosine_reg0 <= 36'sb111111011011110111111010000110000100;
            sine_reg0   <= 36'sb11111111111101011100110110001110100;
        end
        4143: begin
            cosine_reg0 <= 36'sb111111011011000101101001100111011001;
            sine_reg0   <= 36'sb11111111111101010101101011010100001;
        end
        4144: begin
            cosine_reg0 <= 36'sb111111011010010011011001001010001000;
            sine_reg0   <= 36'sb11111111111101001110010110100010010;
        end
        4145: begin
            cosine_reg0 <= 36'sb111111011001100001001000101110010101;
            sine_reg0   <= 36'sb11111111111101000110110111111000110;
        end
        4146: begin
            cosine_reg0 <= 36'sb111111011000101110111000010100000000;
            sine_reg0   <= 36'sb11111111111100111111001111010111110;
        end
        4147: begin
            cosine_reg0 <= 36'sb111111010111111100100111111011001101;
            sine_reg0   <= 36'sb11111111111100110111011100111111001;
        end
        4148: begin
            cosine_reg0 <= 36'sb111111010111001010010111100011111100;
            sine_reg0   <= 36'sb11111111111100101111100000101111000;
        end
        4149: begin
            cosine_reg0 <= 36'sb111111010110011000000111001110010000;
            sine_reg0   <= 36'sb11111111111100100111011010100111011;
        end
        4150: begin
            cosine_reg0 <= 36'sb111111010101100101110110111010001011;
            sine_reg0   <= 36'sb11111111111100011111001010101000010;
        end
        4151: begin
            cosine_reg0 <= 36'sb111111010100110011100110100111101110;
            sine_reg0   <= 36'sb11111111111100010110110000110001101;
        end
        4152: begin
            cosine_reg0 <= 36'sb111111010100000001010110010110111100;
            sine_reg0   <= 36'sb11111111111100001110001101000011011;
        end
        4153: begin
            cosine_reg0 <= 36'sb111111010011001111000110000111110111;
            sine_reg0   <= 36'sb11111111111100000101011111011101110;
        end
        4154: begin
            cosine_reg0 <= 36'sb111111010010011100110101111010011111;
            sine_reg0   <= 36'sb11111111111011111100101000000000100;
        end
        4155: begin
            cosine_reg0 <= 36'sb111111010001101010100101101110111001;
            sine_reg0   <= 36'sb11111111111011110011100110101011110;
        end
        4156: begin
            cosine_reg0 <= 36'sb111111010000111000010101100101000100;
            sine_reg0   <= 36'sb11111111111011101010011011011111101;
        end
        4157: begin
            cosine_reg0 <= 36'sb111111010000000110000101011101000100;
            sine_reg0   <= 36'sb11111111111011100001000110011011111;
        end
        4158: begin
            cosine_reg0 <= 36'sb111111001111010011110101010110111010;
            sine_reg0   <= 36'sb11111111111011010111100111100000110;
        end
        4159: begin
            cosine_reg0 <= 36'sb111111001110100001100101010010101000;
            sine_reg0   <= 36'sb11111111111011001101111110101110001;
        end
        4160: begin
            cosine_reg0 <= 36'sb111111001101101111010101010000010001;
            sine_reg0   <= 36'sb11111111111011000100001100000100000;
        end
        4161: begin
            cosine_reg0 <= 36'sb111111001100111101000101001111110101;
            sine_reg0   <= 36'sb11111111111010111010001111100010100;
        end
        4162: begin
            cosine_reg0 <= 36'sb111111001100001010110101010001010111;
            sine_reg0   <= 36'sb11111111111010110000001001001001011;
        end
        4163: begin
            cosine_reg0 <= 36'sb111111001011011000100101010100111001;
            sine_reg0   <= 36'sb11111111111010100101111000111001000;
        end
        4164: begin
            cosine_reg0 <= 36'sb111111001010100110010101011010011101;
            sine_reg0   <= 36'sb11111111111010011011011110110001000;
        end
        4165: begin
            cosine_reg0 <= 36'sb111111001001110100000101100010000101;
            sine_reg0   <= 36'sb11111111111010010000111010110001101;
        end
        4166: begin
            cosine_reg0 <= 36'sb111111001001000001110101101011110011;
            sine_reg0   <= 36'sb11111111111010000110001100111010111;
        end
        4167: begin
            cosine_reg0 <= 36'sb111111001000001111100101110111101000;
            sine_reg0   <= 36'sb11111111111001111011010101001100101;
        end
        4168: begin
            cosine_reg0 <= 36'sb111111000111011101010110000101100110;
            sine_reg0   <= 36'sb11111111111001110000010011100111000;
        end
        4169: begin
            cosine_reg0 <= 36'sb111111000110101011000110010101110000;
            sine_reg0   <= 36'sb11111111111001100101001000001001111;
        end
        4170: begin
            cosine_reg0 <= 36'sb111111000101111000110110101000001000;
            sine_reg0   <= 36'sb11111111111001011001110010110101011;
        end
        4171: begin
            cosine_reg0 <= 36'sb111111000101000110100110111100101111;
            sine_reg0   <= 36'sb11111111111001001110010011101001100;
        end
        4172: begin
            cosine_reg0 <= 36'sb111111000100010100010111010011100111;
            sine_reg0   <= 36'sb11111111111001000010101010100110010;
        end
        4173: begin
            cosine_reg0 <= 36'sb111111000011100010000111101100110011;
            sine_reg0   <= 36'sb11111111111000110110110111101011101;
        end
        4174: begin
            cosine_reg0 <= 36'sb111111000010101111111000001000010100;
            sine_reg0   <= 36'sb11111111111000101010111010111001101;
        end
        4175: begin
            cosine_reg0 <= 36'sb111111000001111101101000100110001011;
            sine_reg0   <= 36'sb11111111111000011110110100010000010;
        end
        4176: begin
            cosine_reg0 <= 36'sb111111000001001011011001000110011100;
            sine_reg0   <= 36'sb11111111111000010010100011101111011;
        end
        4177: begin
            cosine_reg0 <= 36'sb111111000000011001001001101001001000;
            sine_reg0   <= 36'sb11111111111000000110001001010111010;
        end
        4178: begin
            cosine_reg0 <= 36'sb111110111111100110111010001110010001;
            sine_reg0   <= 36'sb11111111110111111001100101000111111;
        end
        4179: begin
            cosine_reg0 <= 36'sb111110111110110100101010110101111001;
            sine_reg0   <= 36'sb11111111110111101100110111000001000;
        end
        4180: begin
            cosine_reg0 <= 36'sb111110111110000010011011100000000010;
            sine_reg0   <= 36'sb11111111110111011111111111000010111;
        end
        4181: begin
            cosine_reg0 <= 36'sb111110111101010000001100001100101101;
            sine_reg0   <= 36'sb11111111110111010010111101001101011;
        end
        4182: begin
            cosine_reg0 <= 36'sb111110111100011101111100111011111101;
            sine_reg0   <= 36'sb11111111110111000101110001100000101;
        end
        4183: begin
            cosine_reg0 <= 36'sb111110111011101011101101101101110100;
            sine_reg0   <= 36'sb11111111110110111000011011111100100;
        end
        4184: begin
            cosine_reg0 <= 36'sb111110111010111001011110100010010011;
            sine_reg0   <= 36'sb11111111110110101010111100100001000;
        end
        4185: begin
            cosine_reg0 <= 36'sb111110111010000111001111011001011101;
            sine_reg0   <= 36'sb11111111110110011101010011001110011;
        end
        4186: begin
            cosine_reg0 <= 36'sb111110111001010101000000010011010011;
            sine_reg0   <= 36'sb11111111110110001111100000000100011;
        end
        4187: begin
            cosine_reg0 <= 36'sb111110111000100010110001001111110111;
            sine_reg0   <= 36'sb11111111110110000001100011000011001;
        end
        4188: begin
            cosine_reg0 <= 36'sb111110110111110000100010001111001100;
            sine_reg0   <= 36'sb11111111110101110011011100001010100;
        end
        4189: begin
            cosine_reg0 <= 36'sb111110110110111110010011010001010011;
            sine_reg0   <= 36'sb11111111110101100101001011011010110;
        end
        4190: begin
            cosine_reg0 <= 36'sb111110110110001100000100010110001111;
            sine_reg0   <= 36'sb11111111110101010110110000110011101;
        end
        4191: begin
            cosine_reg0 <= 36'sb111110110101011001110101011110000000;
            sine_reg0   <= 36'sb11111111110101001000001100010101011;
        end
        4192: begin
            cosine_reg0 <= 36'sb111110110100100111100110101000101010;
            sine_reg0   <= 36'sb11111111110100111001011101111111111;
        end
        4193: begin
            cosine_reg0 <= 36'sb111110110011110101010111110110001101;
            sine_reg0   <= 36'sb11111111110100101010100101110011001;
        end
        4194: begin
            cosine_reg0 <= 36'sb111110110011000011001001000110101101;
            sine_reg0   <= 36'sb11111111110100011011100011101111001;
        end
        4195: begin
            cosine_reg0 <= 36'sb111110110010010000111010011010001010;
            sine_reg0   <= 36'sb11111111110100001100010111110011111;
        end
        4196: begin
            cosine_reg0 <= 36'sb111110110001011110101011110000100111;
            sine_reg0   <= 36'sb11111111110011111101000010000001100;
        end
        4197: begin
            cosine_reg0 <= 36'sb111110110000101100011101001010000110;
            sine_reg0   <= 36'sb11111111110011101101100010010111111;
        end
        4198: begin
            cosine_reg0 <= 36'sb111110101111111010001110100110101000;
            sine_reg0   <= 36'sb11111111110011011101111000110111001;
        end
        4199: begin
            cosine_reg0 <= 36'sb111110101111001000000000000110010000;
            sine_reg0   <= 36'sb11111111110011001110000101011111010;
        end
        4200: begin
            cosine_reg0 <= 36'sb111110101110010101110001101001000000;
            sine_reg0   <= 36'sb11111111110010111110001000010000001;
        end
        4201: begin
            cosine_reg0 <= 36'sb111110101101100011100011001110111001;
            sine_reg0   <= 36'sb11111111110010101110000001001001111;
        end
        4202: begin
            cosine_reg0 <= 36'sb111110101100110001010100110111111110;
            sine_reg0   <= 36'sb11111111110010011101110000001100100;
        end
        4203: begin
            cosine_reg0 <= 36'sb111110101011111111000110100100010000;
            sine_reg0   <= 36'sb11111111110010001101010101011000000;
        end
        4204: begin
            cosine_reg0 <= 36'sb111110101011001100111000010011110001;
            sine_reg0   <= 36'sb11111111110001111100110000101100011;
        end
        4205: begin
            cosine_reg0 <= 36'sb111110101010011010101010000110100100;
            sine_reg0   <= 36'sb11111111110001101100000010001001101;
        end
        4206: begin
            cosine_reg0 <= 36'sb111110101001101000011011111100101001;
            sine_reg0   <= 36'sb11111111110001011011001001101111110;
        end
        4207: begin
            cosine_reg0 <= 36'sb111110101000110110001101110110000100;
            sine_reg0   <= 36'sb11111111110001001010000111011110110;
        end
        4208: begin
            cosine_reg0 <= 36'sb111110101000000011111111110010110110;
            sine_reg0   <= 36'sb11111111110000111000111011010110110;
        end
        4209: begin
            cosine_reg0 <= 36'sb111110100111010001110001110011000001;
            sine_reg0   <= 36'sb11111111110000100111100101010111101;
        end
        4210: begin
            cosine_reg0 <= 36'sb111110100110011111100011110110100110;
            sine_reg0   <= 36'sb11111111110000010110000101100001100;
        end
        4211: begin
            cosine_reg0 <= 36'sb111110100101101101010101111101101001;
            sine_reg0   <= 36'sb11111111110000000100011011110100010;
        end
        4212: begin
            cosine_reg0 <= 36'sb111110100100111011001000001000001010;
            sine_reg0   <= 36'sb11111111101111110010101000010000000;
        end
        4213: begin
            cosine_reg0 <= 36'sb111110100100001000111010010110001100;
            sine_reg0   <= 36'sb11111111101111100000101010110100101;
        end
        4214: begin
            cosine_reg0 <= 36'sb111110100011010110101100100111110001;
            sine_reg0   <= 36'sb11111111101111001110100011100010011;
        end
        4215: begin
            cosine_reg0 <= 36'sb111110100010100100011110111100111010;
            sine_reg0   <= 36'sb11111111101110111100010010011001000;
        end
        4216: begin
            cosine_reg0 <= 36'sb111110100001110010010001010101101010;
            sine_reg0   <= 36'sb11111111101110101001110111011000110;
        end
        4217: begin
            cosine_reg0 <= 36'sb111110100001000000000011110010000010;
            sine_reg0   <= 36'sb11111111101110010111010010100001011;
        end
        4218: begin
            cosine_reg0 <= 36'sb111110100000001101110110010010000101;
            sine_reg0   <= 36'sb11111111101110000100100011110011001;
        end
        4219: begin
            cosine_reg0 <= 36'sb111110011111011011101000110101110100;
            sine_reg0   <= 36'sb11111111101101110001101011001101111;
        end
        4220: begin
            cosine_reg0 <= 36'sb111110011110101001011011011101010001;
            sine_reg0   <= 36'sb11111111101101011110101000110001110;
        end
        4221: begin
            cosine_reg0 <= 36'sb111110011101110111001110001000011111;
            sine_reg0   <= 36'sb11111111101101001011011100011110101;
        end
        4222: begin
            cosine_reg0 <= 36'sb111110011101000101000000110111011110;
            sine_reg0   <= 36'sb11111111101100111000000110010100100;
        end
        4223: begin
            cosine_reg0 <= 36'sb111110011100010010110011101010010010;
            sine_reg0   <= 36'sb11111111101100100100100110010011100;
        end
        4224: begin
            cosine_reg0 <= 36'sb111110011011100000100110100000111100;
            sine_reg0   <= 36'sb11111111101100010000111100011011101;
        end
        4225: begin
            cosine_reg0 <= 36'sb111110011010101110011001011011011110;
            sine_reg0   <= 36'sb11111111101011111101001000101100111;
        end
        4226: begin
            cosine_reg0 <= 36'sb111110011001111100001100011001111001;
            sine_reg0   <= 36'sb11111111101011101001001011000111010;
        end
        4227: begin
            cosine_reg0 <= 36'sb111110011001001001111111011100010001;
            sine_reg0   <= 36'sb11111111101011010101000011101010110;
        end
        4228: begin
            cosine_reg0 <= 36'sb111110011000010111110010100010100110;
            sine_reg0   <= 36'sb11111111101011000000110010010111011;
        end
        4229: begin
            cosine_reg0 <= 36'sb111110010111100101100101101100111011;
            sine_reg0   <= 36'sb11111111101010101100010111001101001;
        end
        4230: begin
            cosine_reg0 <= 36'sb111110010110110011011000111011010001;
            sine_reg0   <= 36'sb11111111101010010111110010001100000;
        end
        4231: begin
            cosine_reg0 <= 36'sb111110010110000001001100001101101011;
            sine_reg0   <= 36'sb11111111101010000011000011010100001;
        end
        4232: begin
            cosine_reg0 <= 36'sb111110010101001110111111100100001011;
            sine_reg0   <= 36'sb11111111101001101110001010100101011;
        end
        4233: begin
            cosine_reg0 <= 36'sb111110010100011100110010111110110010;
            sine_reg0   <= 36'sb11111111101001011001001000000000000;
        end
        4234: begin
            cosine_reg0 <= 36'sb111110010011101010100110011101100010;
            sine_reg0   <= 36'sb11111111101001000011111011100011101;
        end
        4235: begin
            cosine_reg0 <= 36'sb111110010010111000011010000000011110;
            sine_reg0   <= 36'sb11111111101000101110100101010000101;
        end
        4236: begin
            cosine_reg0 <= 36'sb111110010010000110001101100111100110;
            sine_reg0   <= 36'sb11111111101000011001000101000110111;
        end
        4237: begin
            cosine_reg0 <= 36'sb111110010001010100000001010010111110;
            sine_reg0   <= 36'sb11111111101000000011011011000110010;
        end
        4238: begin
            cosine_reg0 <= 36'sb111110010000100001110101000010101000;
            sine_reg0   <= 36'sb11111111100111101101100111001111000;
        end
        4239: begin
            cosine_reg0 <= 36'sb111110001111101111101000110110100100;
            sine_reg0   <= 36'sb11111111100111010111101001100001000;
        end
        4240: begin
            cosine_reg0 <= 36'sb111110001110111101011100101110110101;
            sine_reg0   <= 36'sb11111111100111000001100001111100010;
        end
        4241: begin
            cosine_reg0 <= 36'sb111110001110001011010000101011011101;
            sine_reg0   <= 36'sb11111111100110101011010000100000111;
        end
        4242: begin
            cosine_reg0 <= 36'sb111110001101011001000100101100011110;
            sine_reg0   <= 36'sb11111111100110010100110101001110111;
        end
        4243: begin
            cosine_reg0 <= 36'sb111110001100100110111000110001111010;
            sine_reg0   <= 36'sb11111111100101111110010000000110001;
        end
        4244: begin
            cosine_reg0 <= 36'sb111110001011110100101100111011110010;
            sine_reg0   <= 36'sb11111111100101100111100001000110110;
        end
        4245: begin
            cosine_reg0 <= 36'sb111110001011000010100001001010001001;
            sine_reg0   <= 36'sb11111111100101010000101000010000101;
        end
        4246: begin
            cosine_reg0 <= 36'sb111110001010010000010101011101000001;
            sine_reg0   <= 36'sb11111111100100111001100101100100000;
        end
        4247: begin
            cosine_reg0 <= 36'sb111110001001011110001001110100011011;
            sine_reg0   <= 36'sb11111111100100100010011001000000110;
        end
        4248: begin
            cosine_reg0 <= 36'sb111110001000101011111110010000011010;
            sine_reg0   <= 36'sb11111111100100001011000010100110111;
        end
        4249: begin
            cosine_reg0 <= 36'sb111110000111111001110010110000111111;
            sine_reg0   <= 36'sb11111111100011110011100010010110100;
        end
        4250: begin
            cosine_reg0 <= 36'sb111110000111000111100111010110001101;
            sine_reg0   <= 36'sb11111111100011011011111000001111100;
        end
        4251: begin
            cosine_reg0 <= 36'sb111110000110010101011100000000000100;
            sine_reg0   <= 36'sb11111111100011000100000100010001111;
        end
        4252: begin
            cosine_reg0 <= 36'sb111110000101100011010000101110101000;
            sine_reg0   <= 36'sb11111111100010101100000110011101111;
        end
        4253: begin
            cosine_reg0 <= 36'sb111110000100110001000101100001111010;
            sine_reg0   <= 36'sb11111111100010010011111110110011010;
        end
        4254: begin
            cosine_reg0 <= 36'sb111110000011111110111010011001111100;
            sine_reg0   <= 36'sb11111111100001111011101101010010000;
        end
        4255: begin
            cosine_reg0 <= 36'sb111110000011001100101111010110110000;
            sine_reg0   <= 36'sb11111111100001100011010001111010011;
        end
        4256: begin
            cosine_reg0 <= 36'sb111110000010011010100100011000011000;
            sine_reg0   <= 36'sb11111111100001001010101100101100011;
        end
        4257: begin
            cosine_reg0 <= 36'sb111110000001101000011001011110110110;
            sine_reg0   <= 36'sb11111111100000110001111101100111110;
        end
        4258: begin
            cosine_reg0 <= 36'sb111110000000110110001110101010001100;
            sine_reg0   <= 36'sb11111111100000011001000100101100110;
        end
        4259: begin
            cosine_reg0 <= 36'sb111110000000000100000011111010011011;
            sine_reg0   <= 36'sb11111111100000000000000001111011010;
        end
        4260: begin
            cosine_reg0 <= 36'sb111101111111010001111001001111100110;
            sine_reg0   <= 36'sb11111111011111100110110101010011011;
        end
        4261: begin
            cosine_reg0 <= 36'sb111101111110011111101110101001101111;
            sine_reg0   <= 36'sb11111111011111001101011110110101001;
        end
        4262: begin
            cosine_reg0 <= 36'sb111101111101101101100100001000110111;
            sine_reg0   <= 36'sb11111111011110110011111110100000011;
        end
        4263: begin
            cosine_reg0 <= 36'sb111101111100111011011001101101000001;
            sine_reg0   <= 36'sb11111111011110011010010100010101011;
        end
        4264: begin
            cosine_reg0 <= 36'sb111101111100001001001111010110001110;
            sine_reg0   <= 36'sb11111111011110000000100000010100000;
        end
        4265: begin
            cosine_reg0 <= 36'sb111101111011010111000101000100100000;
            sine_reg0   <= 36'sb11111111011101100110100010011100010;
        end
        4266: begin
            cosine_reg0 <= 36'sb111101111010100100111010110111111010;
            sine_reg0   <= 36'sb11111111011101001100011010101110001;
        end
        4267: begin
            cosine_reg0 <= 36'sb111101111001110010110000110000011101;
            sine_reg0   <= 36'sb11111111011100110010001001001001110;
        end
        4268: begin
            cosine_reg0 <= 36'sb111101111001000000100110101110001011;
            sine_reg0   <= 36'sb11111111011100010111101101101111000;
        end
        4269: begin
            cosine_reg0 <= 36'sb111101111000001110011100110001000110;
            sine_reg0   <= 36'sb11111111011011111101001000011110000;
        end
        4270: begin
            cosine_reg0 <= 36'sb111101110111011100010010111001010000;
            sine_reg0   <= 36'sb11111111011011100010011001010110110;
        end
        4271: begin
            cosine_reg0 <= 36'sb111101110110101010001001000110101011;
            sine_reg0   <= 36'sb11111111011011000111100000011001010;
        end
        4272: begin
            cosine_reg0 <= 36'sb111101110101110111111111011001011001;
            sine_reg0   <= 36'sb11111111011010101100011101100101101;
        end
        4273: begin
            cosine_reg0 <= 36'sb111101110101000101110101110001011100;
            sine_reg0   <= 36'sb11111111011010010001010000111011101;
        end
        4274: begin
            cosine_reg0 <= 36'sb111101110100010011101100001110110110;
            sine_reg0   <= 36'sb11111111011001110101111010011011100;
        end
        4275: begin
            cosine_reg0 <= 36'sb111101110011100001100010110001101000;
            sine_reg0   <= 36'sb11111111011001011010011010000101001;
        end
        4276: begin
            cosine_reg0 <= 36'sb111101110010101111011001011001110101;
            sine_reg0   <= 36'sb11111111011000111110101111111000101;
        end
        4277: begin
            cosine_reg0 <= 36'sb111101110001111101010000000111011110;
            sine_reg0   <= 36'sb11111111011000100010111011110110000;
        end
        4278: begin
            cosine_reg0 <= 36'sb111101110001001011000110111010100110;
            sine_reg0   <= 36'sb11111111011000000110111101111101010;
        end
        4279: begin
            cosine_reg0 <= 36'sb111101110000011000111101110011001110;
            sine_reg0   <= 36'sb11111111010111101010110110001110011;
        end
        4280: begin
            cosine_reg0 <= 36'sb111101101111100110110100110001011001;
            sine_reg0   <= 36'sb11111111010111001110100100101001011;
        end
        4281: begin
            cosine_reg0 <= 36'sb111101101110110100101011110101001000;
            sine_reg0   <= 36'sb11111111010110110010001001001110010;
        end
        4282: begin
            cosine_reg0 <= 36'sb111101101110000010100010111110011101;
            sine_reg0   <= 36'sb11111111010110010101100011111101001;
        end
        4283: begin
            cosine_reg0 <= 36'sb111101101101010000011010001101011010;
            sine_reg0   <= 36'sb11111111010101111000110100110110000;
        end
        4284: begin
            cosine_reg0 <= 36'sb111101101100011110010001100010000001;
            sine_reg0   <= 36'sb11111111010101011011111011111000110;
        end
        4285: begin
            cosine_reg0 <= 36'sb111101101011101100001000111100010100;
            sine_reg0   <= 36'sb11111111010100111110111001000101100;
        end
        4286: begin
            cosine_reg0 <= 36'sb111101101010111010000000011100010110;
            sine_reg0   <= 36'sb11111111010100100001101100011100010;
        end
        4287: begin
            cosine_reg0 <= 36'sb111101101010000111111000000010000111;
            sine_reg0   <= 36'sb11111111010100000100010101111101001;
        end
        4288: begin
            cosine_reg0 <= 36'sb111101101001010101101111101101101010;
            sine_reg0   <= 36'sb11111111010011100110110101100111111;
        end
        4289: begin
            cosine_reg0 <= 36'sb111101101000100011100111011111000000;
            sine_reg0   <= 36'sb11111111010011001001001011011100110;
        end
        4290: begin
            cosine_reg0 <= 36'sb111101100111110001011111010110001101;
            sine_reg0   <= 36'sb11111111010010101011010111011011110;
        end
        4291: begin
            cosine_reg0 <= 36'sb111101100110111111010111010011010001;
            sine_reg0   <= 36'sb11111111010010001101011001100100111;
        end
        4292: begin
            cosine_reg0 <= 36'sb111101100110001101001111010110001110;
            sine_reg0   <= 36'sb11111111010001101111010001111000000;
        end
        4293: begin
            cosine_reg0 <= 36'sb111101100101011011000111011111000111;
            sine_reg0   <= 36'sb11111111010001010001000000010101010;
        end
        4294: begin
            cosine_reg0 <= 36'sb111101100100101000111111101101111101;
            sine_reg0   <= 36'sb11111111010000110010100100111100110;
        end
        4295: begin
            cosine_reg0 <= 36'sb111101100011110110111000000010110011;
            sine_reg0   <= 36'sb11111111010000010011111111101110011;
        end
        4296: begin
            cosine_reg0 <= 36'sb111101100011000100110000011101101010;
            sine_reg0   <= 36'sb11111111001111110101010000101010001;
        end
        4297: begin
            cosine_reg0 <= 36'sb111101100010010010101000111110100100;
            sine_reg0   <= 36'sb11111111001111010110010111110000001;
        end
        4298: begin
            cosine_reg0 <= 36'sb111101100001100000100001100101100011;
            sine_reg0   <= 36'sb11111111001110110111010101000000011;
        end
        4299: begin
            cosine_reg0 <= 36'sb111101100000101110011010010010101010;
            sine_reg0   <= 36'sb11111111001110011000001000011010110;
        end
        4300: begin
            cosine_reg0 <= 36'sb111101011111111100010011000101111001;
            sine_reg0   <= 36'sb11111111001101111000110001111111100;
        end
        4301: begin
            cosine_reg0 <= 36'sb111101011111001010001011111111010011;
            sine_reg0   <= 36'sb11111111001101011001010001101110100;
        end
        4302: begin
            cosine_reg0 <= 36'sb111101011110011000000100111110111010;
            sine_reg0   <= 36'sb11111111001100111001100111100111110;
        end
        4303: begin
            cosine_reg0 <= 36'sb111101011101100101111110000100110000;
            sine_reg0   <= 36'sb11111111001100011001110011101011011;
        end
        4304: begin
            cosine_reg0 <= 36'sb111101011100110011110111010000110111;
            sine_reg0   <= 36'sb11111111001011111001110101111001011;
        end
        4305: begin
            cosine_reg0 <= 36'sb111101011100000001110000100011010000;
            sine_reg0   <= 36'sb11111111001011011001101110010001101;
        end
        4306: begin
            cosine_reg0 <= 36'sb111101011011001111101001111011111110;
            sine_reg0   <= 36'sb11111111001010111001011100110100010;
        end
        4307: begin
            cosine_reg0 <= 36'sb111101011010011101100011011011000010;
            sine_reg0   <= 36'sb11111111001010011001000001100001011;
        end
        4308: begin
            cosine_reg0 <= 36'sb111101011001101011011101000000011111;
            sine_reg0   <= 36'sb11111111001001111000011100011000110;
        end
        4309: begin
            cosine_reg0 <= 36'sb111101011000111001010110101100010110;
            sine_reg0   <= 36'sb11111111001001010111101101011010110;
        end
        4310: begin
            cosine_reg0 <= 36'sb111101011000000111010000011110101010;
            sine_reg0   <= 36'sb11111111001000110110110100100111000;
        end
        4311: begin
            cosine_reg0 <= 36'sb111101010111010101001010010111011100;
            sine_reg0   <= 36'sb11111111001000010101110001111101111;
        end
        4312: begin
            cosine_reg0 <= 36'sb111101010110100011000100010110101110;
            sine_reg0   <= 36'sb11111111000111110100100101011111001;
        end
        4313: begin
            cosine_reg0 <= 36'sb111101010101110000111110011100100010;
            sine_reg0   <= 36'sb11111111000111010011001111001011000;
        end
        4314: begin
            cosine_reg0 <= 36'sb111101010100111110111000101000111010;
            sine_reg0   <= 36'sb11111111000110110001101111000001011;
        end
        4315: begin
            cosine_reg0 <= 36'sb111101010100001100110010111011111000;
            sine_reg0   <= 36'sb11111111000110010000000101000010010;
        end
        4316: begin
            cosine_reg0 <= 36'sb111101010011011010101101010101011110;
            sine_reg0   <= 36'sb11111111000101101110010001001101110;
        end
        4317: begin
            cosine_reg0 <= 36'sb111101010010101000100111110101101110;
            sine_reg0   <= 36'sb11111111000101001100010011100011111;
        end
        4318: begin
            cosine_reg0 <= 36'sb111101010001110110100010011100101001;
            sine_reg0   <= 36'sb11111111000100101010001100000100100;
        end
        4319: begin
            cosine_reg0 <= 36'sb111101010001000100011101001010010010;
            sine_reg0   <= 36'sb11111111000100000111111010101111111;
        end
        4320: begin
            cosine_reg0 <= 36'sb111101010000010010010111111110101011;
            sine_reg0   <= 36'sb11111111000011100101011111100101110;
        end
        4321: begin
            cosine_reg0 <= 36'sb111101001111100000010010111001110110;
            sine_reg0   <= 36'sb11111111000011000010111010100110100;
        end
        4322: begin
            cosine_reg0 <= 36'sb111101001110101110001101111011110100;
            sine_reg0   <= 36'sb11111111000010100000001011110001110;
        end
        4323: begin
            cosine_reg0 <= 36'sb111101001101111100001001000100100111;
            sine_reg0   <= 36'sb11111111000001111101010011000111111;
        end
        4324: begin
            cosine_reg0 <= 36'sb111101001101001010000100010100010010;
            sine_reg0   <= 36'sb11111111000001011010010000101000101;
        end
        4325: begin
            cosine_reg0 <= 36'sb111101001100010111111111101010110101;
            sine_reg0   <= 36'sb11111111000000110111000100010100001;
        end
        4326: begin
            cosine_reg0 <= 36'sb111101001011100101111011001000010101;
            sine_reg0   <= 36'sb11111111000000010011101110001010100;
        end
        4327: begin
            cosine_reg0 <= 36'sb111101001010110011110110101100110001;
            sine_reg0   <= 36'sb11111110111111110000001110001011101;
        end
        4328: begin
            cosine_reg0 <= 36'sb111101001010000001110010011000001100;
            sine_reg0   <= 36'sb11111110111111001100100100010111101;
        end
        4329: begin
            cosine_reg0 <= 36'sb111101001001001111101110001010101001;
            sine_reg0   <= 36'sb11111110111110101000110000101110011;
        end
        4330: begin
            cosine_reg0 <= 36'sb111101001000011101101010000100001000;
            sine_reg0   <= 36'sb11111110111110000100110011010000001;
        end
        4331: begin
            cosine_reg0 <= 36'sb111101000111101011100110000100101100;
            sine_reg0   <= 36'sb11111110111101100000101011111100101;
        end
        4332: begin
            cosine_reg0 <= 36'sb111101000110111001100010001100010111;
            sine_reg0   <= 36'sb11111110111100111100011010110100001;
        end
        4333: begin
            cosine_reg0 <= 36'sb111101000110000111011110011011001011;
            sine_reg0   <= 36'sb11111110111100010111111111110110100;
        end
        4334: begin
            cosine_reg0 <= 36'sb111101000101010101011010110001001001;
            sine_reg0   <= 36'sb11111110111011110011011011000011110;
        end
        4335: begin
            cosine_reg0 <= 36'sb111101000100100011010111001110010100;
            sine_reg0   <= 36'sb11111110111011001110101100011100001;
        end
        4336: begin
            cosine_reg0 <= 36'sb111101000011110001010011110010101101;
            sine_reg0   <= 36'sb11111110111010101001110011111111011;
        end
        4337: begin
            cosine_reg0 <= 36'sb111101000010111111010000011110010111;
            sine_reg0   <= 36'sb11111110111010000100110001101101110;
        end
        4338: begin
            cosine_reg0 <= 36'sb111101000010001101001101010001010011;
            sine_reg0   <= 36'sb11111110111001011111100101100111001;
        end
        4339: begin
            cosine_reg0 <= 36'sb111101000001011011001010001011100100;
            sine_reg0   <= 36'sb11111110111000111010001111101011101;
        end
        4340: begin
            cosine_reg0 <= 36'sb111101000000101001000111001101001010;
            sine_reg0   <= 36'sb11111110111000010100101111111011001;
        end
        4341: begin
            cosine_reg0 <= 36'sb111100111111110111000100010110001001;
            sine_reg0   <= 36'sb11111110110111101111000110010101110;
        end
        4342: begin
            cosine_reg0 <= 36'sb111100111111000101000001100110100010;
            sine_reg0   <= 36'sb11111110110111001001010010111011100;
        end
        4343: begin
            cosine_reg0 <= 36'sb111100111110010010111110111110010111;
            sine_reg0   <= 36'sb11111110110110100011010101101100011;
        end
        4344: begin
            cosine_reg0 <= 36'sb111100111101100000111100011101101010;
            sine_reg0   <= 36'sb11111110110101111101001110101000100;
        end
        4345: begin
            cosine_reg0 <= 36'sb111100111100101110111010000100011101;
            sine_reg0   <= 36'sb11111110110101010110111101101111110;
        end
        4346: begin
            cosine_reg0 <= 36'sb111100111011111100110111110010110001;
            sine_reg0   <= 36'sb11111110110100110000100011000010011;
        end
        4347: begin
            cosine_reg0 <= 36'sb111100111011001010110101101000101010;
            sine_reg0   <= 36'sb11111110110100001001111110100000001;
        end
        4348: begin
            cosine_reg0 <= 36'sb111100111010011000110011100110001000;
            sine_reg0   <= 36'sb11111110110011100011010000001001001;
        end
        4349: begin
            cosine_reg0 <= 36'sb111100111001100110110001101011001101;
            sine_reg0   <= 36'sb11111110110010111100010111111101100;
        end
        4350: begin
            cosine_reg0 <= 36'sb111100111000110100101111110111111100;
            sine_reg0   <= 36'sb11111110110010010101010101111101001;
        end
        4351: begin
            cosine_reg0 <= 36'sb111100111000000010101110001100010111;
            sine_reg0   <= 36'sb11111110110001101110001010001000001;
        end
        4352: begin
            cosine_reg0 <= 36'sb111100110111010000101100101000011111;
            sine_reg0   <= 36'sb11111110110001000110110100011110011;
        end
        4353: begin
            cosine_reg0 <= 36'sb111100110110011110101011001100010110;
            sine_reg0   <= 36'sb11111110110000011111010101000000001;
        end
        4354: begin
            cosine_reg0 <= 36'sb111100110101101100101001110111111110;
            sine_reg0   <= 36'sb11111110101111110111101011101101010;
        end
        4355: begin
            cosine_reg0 <= 36'sb111100110100111010101000101011011010;
            sine_reg0   <= 36'sb11111110101111001111111000100101111;
        end
        4356: begin
            cosine_reg0 <= 36'sb111100110100001000100111100110101011;
            sine_reg0   <= 36'sb11111110101110100111111011101001111;
        end
        4357: begin
            cosine_reg0 <= 36'sb111100110011010110100110101001110010;
            sine_reg0   <= 36'sb11111110101101111111110100111001011;
        end
        4358: begin
            cosine_reg0 <= 36'sb111100110010100100100101110100110011;
            sine_reg0   <= 36'sb11111110101101010111100100010100100;
        end
        4359: begin
            cosine_reg0 <= 36'sb111100110001110010100101000111101111;
            sine_reg0   <= 36'sb11111110101100101111001001111011000;
        end
        4360: begin
            cosine_reg0 <= 36'sb111100110001000000100100100010100111;
            sine_reg0   <= 36'sb11111110101100000110100101101101001;
        end
        4361: begin
            cosine_reg0 <= 36'sb111100110000001110100100000101011110;
            sine_reg0   <= 36'sb11111110101011011101110111101010110;
        end
        4362: begin
            cosine_reg0 <= 36'sb111100101111011100100011110000010110;
            sine_reg0   <= 36'sb11111110101010110100111111110100001;
        end
        4363: begin
            cosine_reg0 <= 36'sb111100101110101010100011100011010000;
            sine_reg0   <= 36'sb11111110101010001011111110001001000;
        end
        4364: begin
            cosine_reg0 <= 36'sb111100101101111000100011011110001111;
            sine_reg0   <= 36'sb11111110101001100010110010101001101;
        end
        4365: begin
            cosine_reg0 <= 36'sb111100101101000110100011100001010100;
            sine_reg0   <= 36'sb11111110101000111001011101010101111;
        end
        4366: begin
            cosine_reg0 <= 36'sb111100101100010100100011101100100010;
            sine_reg0   <= 36'sb11111110101000001111111110001101110;
        end
        4367: begin
            cosine_reg0 <= 36'sb111100101011100010100011111111111010;
            sine_reg0   <= 36'sb11111110100111100110010101010001100;
        end
        4368: begin
            cosine_reg0 <= 36'sb111100101010110000100100011011011110;
            sine_reg0   <= 36'sb11111110100110111100100010100001000;
        end
        4369: begin
            cosine_reg0 <= 36'sb111100101001111110100100111111010000;
            sine_reg0   <= 36'sb11111110100110010010100101111100001;
        end
        4370: begin
            cosine_reg0 <= 36'sb111100101001001100100101101011010010;
            sine_reg0   <= 36'sb11111110100101101000011111100011001;
        end
        4371: begin
            cosine_reg0 <= 36'sb111100101000011010100110011111100111;
            sine_reg0   <= 36'sb11111110100100111110001111010110000;
        end
        4372: begin
            cosine_reg0 <= 36'sb111100100111101000100111011100001111;
            sine_reg0   <= 36'sb11111110100100010011110101010100110;
        end
        4373: begin
            cosine_reg0 <= 36'sb111100100110110110101000100001001101;
            sine_reg0   <= 36'sb11111110100011101001010001011111011;
        end
        4374: begin
            cosine_reg0 <= 36'sb111100100110000100101001101110100011;
            sine_reg0   <= 36'sb11111110100010111110100011110101111;
        end
        4375: begin
            cosine_reg0 <= 36'sb111100100101010010101011000100010011;
            sine_reg0   <= 36'sb11111110100010010011101100011000010;
        end
        4376: begin
            cosine_reg0 <= 36'sb111100100100100000101100100010011110;
            sine_reg0   <= 36'sb11111110100001101000101011000110101;
        end
        4377: begin
            cosine_reg0 <= 36'sb111100100011101110101110001001000111;
            sine_reg0   <= 36'sb11111110100000111101100000000001000;
        end
        4378: begin
            cosine_reg0 <= 36'sb111100100010111100101111111000010000;
            sine_reg0   <= 36'sb11111110100000010010001011000111011;
        end
        4379: begin
            cosine_reg0 <= 36'sb111100100010001010110001101111111001;
            sine_reg0   <= 36'sb11111110011111100110101100011001110;
        end
        4380: begin
            cosine_reg0 <= 36'sb111100100001011000110011110000000111;
            sine_reg0   <= 36'sb11111110011110111011000011111000010;
        end
        4381: begin
            cosine_reg0 <= 36'sb111100100000100110110101111000111001;
            sine_reg0   <= 36'sb11111110011110001111010001100010111;
        end
        4382: begin
            cosine_reg0 <= 36'sb111100011111110100111000001010010011;
            sine_reg0   <= 36'sb11111110011101100011010101011001100;
        end
        4383: begin
            cosine_reg0 <= 36'sb111100011111000010111010100100010101;
            sine_reg0   <= 36'sb11111110011100110111001111011100011;
        end
        4384: begin
            cosine_reg0 <= 36'sb111100011110010000111101000111000011;
            sine_reg0   <= 36'sb11111110011100001010111111101011010;
        end
        4385: begin
            cosine_reg0 <= 36'sb111100011101011110111111110010011110;
            sine_reg0   <= 36'sb11111110011011011110100110000110100;
        end
        4386: begin
            cosine_reg0 <= 36'sb111100011100101101000010100110101000;
            sine_reg0   <= 36'sb11111110011010110010000010101101111;
        end
        4387: begin
            cosine_reg0 <= 36'sb111100011011111011000101100011100010;
            sine_reg0   <= 36'sb11111110011010000101010101100001100;
        end
        4388: begin
            cosine_reg0 <= 36'sb111100011011001001001000101001001111;
            sine_reg0   <= 36'sb11111110011001011000011110100001100;
        end
        4389: begin
            cosine_reg0 <= 36'sb111100011010010111001011110111110001;
            sine_reg0   <= 36'sb11111110011000101011011101101101101;
        end
        4390: begin
            cosine_reg0 <= 36'sb111100011001100101001111001111001010;
            sine_reg0   <= 36'sb11111110010111111110010011000110010;
        end
        4391: begin
            cosine_reg0 <= 36'sb111100011000110011010010101111011011;
            sine_reg0   <= 36'sb11111110010111010000111110101011001;
        end
        4392: begin
            cosine_reg0 <= 36'sb111100011000000001010110011000100111;
            sine_reg0   <= 36'sb11111110010110100011100000011100011;
        end
        4393: begin
            cosine_reg0 <= 36'sb111100010111001111011010001010101111;
            sine_reg0   <= 36'sb11111110010101110101111000011010001;
        end
        4394: begin
            cosine_reg0 <= 36'sb111100010110011101011110000101110101;
            sine_reg0   <= 36'sb11111110010101001000000110100100010;
        end
        4395: begin
            cosine_reg0 <= 36'sb111100010101101011100010001001111011;
            sine_reg0   <= 36'sb11111110010100011010001010111010111;
        end
        4396: begin
            cosine_reg0 <= 36'sb111100010100111001100110010111000100;
            sine_reg0   <= 36'sb11111110010011101100000101011110000;
        end
        4397: begin
            cosine_reg0 <= 36'sb111100010100000111101010101101010001;
            sine_reg0   <= 36'sb11111110010010111101110110001101101;
        end
        4398: begin
            cosine_reg0 <= 36'sb111100010011010101101111001100100011;
            sine_reg0   <= 36'sb11111110010010001111011101001001110;
        end
        4399: begin
            cosine_reg0 <= 36'sb111100010010100011110011110100111110;
            sine_reg0   <= 36'sb11111110010001100000111010010010100;
        end
        4400: begin
            cosine_reg0 <= 36'sb111100010001110001111000100110100011;
            sine_reg0   <= 36'sb11111110010000110010001101100111111;
        end
        4401: begin
            cosine_reg0 <= 36'sb111100010000111111111101100001010011;
            sine_reg0   <= 36'sb11111110010000000011010111001001111;
        end
        4402: begin
            cosine_reg0 <= 36'sb111100010000001110000010100101010001;
            sine_reg0   <= 36'sb11111110001111010100010110111000100;
        end
        4403: begin
            cosine_reg0 <= 36'sb111100001111011100000111110010011111;
            sine_reg0   <= 36'sb11111110001110100101001100110011110;
        end
        4404: begin
            cosine_reg0 <= 36'sb111100001110101010001101001000111110;
            sine_reg0   <= 36'sb11111110001101110101111000111011111;
        end
        4405: begin
            cosine_reg0 <= 36'sb111100001101111000010010101000110001;
            sine_reg0   <= 36'sb11111110001101000110011011010000101;
        end
        4406: begin
            cosine_reg0 <= 36'sb111100001101000110011000010001111001;
            sine_reg0   <= 36'sb11111110001100010110110011110010010;
        end
        4407: begin
            cosine_reg0 <= 36'sb111100001100010100011110000100011000;
            sine_reg0   <= 36'sb11111110001011100111000010100000101;
        end
        4408: begin
            cosine_reg0 <= 36'sb111100001011100010100100000000010001;
            sine_reg0   <= 36'sb11111110001010110111000111011011110;
        end
        4409: begin
            cosine_reg0 <= 36'sb111100001010110000101010000101100101;
            sine_reg0   <= 36'sb11111110001010000111000010100011111;
        end
        4410: begin
            cosine_reg0 <= 36'sb111100001001111110110000010100010110;
            sine_reg0   <= 36'sb11111110001001010110110011111000111;
        end
        4411: begin
            cosine_reg0 <= 36'sb111100001001001100110110101100100110;
            sine_reg0   <= 36'sb11111110001000100110011011011010110;
        end
        4412: begin
            cosine_reg0 <= 36'sb111100001000011010111101001110010111;
            sine_reg0   <= 36'sb11111110000111110101111001001001100;
        end
        4413: begin
            cosine_reg0 <= 36'sb111100000111101001000011111001101011;
            sine_reg0   <= 36'sb11111110000111000101001101000101011;
        end
        4414: begin
            cosine_reg0 <= 36'sb111100000110110111001010101110100011;
            sine_reg0   <= 36'sb11111110000110010100010111001110001;
        end
        4415: begin
            cosine_reg0 <= 36'sb111100000110000101010001101101000011;
            sine_reg0   <= 36'sb11111110000101100011010111100100000;
        end
        4416: begin
            cosine_reg0 <= 36'sb111100000101010011011000110101001011;
            sine_reg0   <= 36'sb11111110000100110010001110000110111;
        end
        4417: begin
            cosine_reg0 <= 36'sb111100000100100001100000000110111101;
            sine_reg0   <= 36'sb11111110000100000000111010110111000;
        end
        4418: begin
            cosine_reg0 <= 36'sb111100000011101111100111100010011101;
            sine_reg0   <= 36'sb11111110000011001111011101110100001;
        end
        4419: begin
            cosine_reg0 <= 36'sb111100000010111101101111000111101010;
            sine_reg0   <= 36'sb11111110000010011101110110111110011;
        end
        4420: begin
            cosine_reg0 <= 36'sb111100000010001011110110110110101000;
            sine_reg0   <= 36'sb11111110000001101100000110010101111;
        end
        4421: begin
            cosine_reg0 <= 36'sb111100000001011001111110101111011000;
            sine_reg0   <= 36'sb11111110000000111010001011111010100;
        end
        4422: begin
            cosine_reg0 <= 36'sb111100000000101000000110110001111100;
            sine_reg0   <= 36'sb11111110000000001000000111101100100;
        end
        4423: begin
            cosine_reg0 <= 36'sb111011111111110110001110111110010111;
            sine_reg0   <= 36'sb11111101111111010101111001101011110;
        end
        4424: begin
            cosine_reg0 <= 36'sb111011111111000100010111010100101001;
            sine_reg0   <= 36'sb11111101111110100011100001111000010;
        end
        4425: begin
            cosine_reg0 <= 36'sb111011111110010010011111110100110110;
            sine_reg0   <= 36'sb11111101111101110001000000010010000;
        end
        4426: begin
            cosine_reg0 <= 36'sb111011111101100000101000011110111110;
            sine_reg0   <= 36'sb11111101111100111110010100111001010;
        end
        4427: begin
            cosine_reg0 <= 36'sb111011111100101110110001010011000100;
            sine_reg0   <= 36'sb11111101111100001011011111101101111;
        end
        4428: begin
            cosine_reg0 <= 36'sb111011111011111100111010010001001010;
            sine_reg0   <= 36'sb11111101111011011000100000110000000;
        end
        4429: begin
            cosine_reg0 <= 36'sb111011111011001011000011011001010001;
            sine_reg0   <= 36'sb11111101111010100101010111111111100;
        end
        4430: begin
            cosine_reg0 <= 36'sb111011111010011001001100101011011100;
            sine_reg0   <= 36'sb11111101111001110010000101011100011;
        end
        4431: begin
            cosine_reg0 <= 36'sb111011111001100111010110000111101101;
            sine_reg0   <= 36'sb11111101111000111110101001000111000;
        end
        4432: begin
            cosine_reg0 <= 36'sb111011111000110101011111101110000100;
            sine_reg0   <= 36'sb11111101111000001011000010111111000;
        end
        4433: begin
            cosine_reg0 <= 36'sb111011111000000011101001011110100110;
            sine_reg0   <= 36'sb11111101110111010111010011000100101;
        end
        4434: begin
            cosine_reg0 <= 36'sb111011110111010001110011011001010010;
            sine_reg0   <= 36'sb11111101110110100011011001010111111;
        end
        4435: begin
            cosine_reg0 <= 36'sb111011110110011111111101011110001100;
            sine_reg0   <= 36'sb11111101110101101111010101111000110;
        end
        4436: begin
            cosine_reg0 <= 36'sb111011110101101110000111101101010101;
            sine_reg0   <= 36'sb11111101110100111011001000100111011;
        end
        4437: begin
            cosine_reg0 <= 36'sb111011110100111100010010000110101110;
            sine_reg0   <= 36'sb11111101110100000110110001100011101;
        end
        4438: begin
            cosine_reg0 <= 36'sb111011110100001010011100101010011011;
            sine_reg0   <= 36'sb11111101110011010010010000101101110;
        end
        4439: begin
            cosine_reg0 <= 36'sb111011110011011000100111011000011101;
            sine_reg0   <= 36'sb11111101110010011101100110000101100;
        end
        4440: begin
            cosine_reg0 <= 36'sb111011110010100110110010010000110101;
            sine_reg0   <= 36'sb11111101110001101000110001101011001;
        end
        4441: begin
            cosine_reg0 <= 36'sb111011110001110100111101010011100110;
            sine_reg0   <= 36'sb11111101110000110011110011011110100;
        end
        4442: begin
            cosine_reg0 <= 36'sb111011110001000011001000100000110010;
            sine_reg0   <= 36'sb11111101101111111110101011011111110;
        end
        4443: begin
            cosine_reg0 <= 36'sb111011110000010001010011111000011010;
            sine_reg0   <= 36'sb11111101101111001001011001101111000;
        end
        4444: begin
            cosine_reg0 <= 36'sb111011101111011111011111011010100001;
            sine_reg0   <= 36'sb11111101101110010011111110001100001;
        end
        4445: begin
            cosine_reg0 <= 36'sb111011101110101101101011000111001000;
            sine_reg0   <= 36'sb11111101101101011110011000110111010;
        end
        4446: begin
            cosine_reg0 <= 36'sb111011101101111011110110111110010001;
            sine_reg0   <= 36'sb11111101101100101000101001110000010;
        end
        4447: begin
            cosine_reg0 <= 36'sb111011101101001010000010111111111111;
            sine_reg0   <= 36'sb11111101101011110010110000110111011;
        end
        4448: begin
            cosine_reg0 <= 36'sb111011101100011000001111001100010010;
            sine_reg0   <= 36'sb11111101101010111100101110001100100;
        end
        4449: begin
            cosine_reg0 <= 36'sb111011101011100110011011100011001110;
            sine_reg0   <= 36'sb11111101101010000110100001101111111;
        end
        4450: begin
            cosine_reg0 <= 36'sb111011101010110100101000000100110100;
            sine_reg0   <= 36'sb11111101101001010000001011100001010;
        end
        4451: begin
            cosine_reg0 <= 36'sb111011101010000010110100110001000110;
            sine_reg0   <= 36'sb11111101101000011001101011100000110;
        end
        4452: begin
            cosine_reg0 <= 36'sb111011101001010001000001101000000101;
            sine_reg0   <= 36'sb11111101100111100011000001101110100;
        end
        4453: begin
            cosine_reg0 <= 36'sb111011101000011111001110101001110101;
            sine_reg0   <= 36'sb11111101100110101100001110001010011;
        end
        4454: begin
            cosine_reg0 <= 36'sb111011100111101101011011110110010110;
            sine_reg0   <= 36'sb11111101100101110101010000110100101;
        end
        4455: begin
            cosine_reg0 <= 36'sb111011100110111011101001001101101010;
            sine_reg0   <= 36'sb11111101100100111110001001101101001;
        end
        4456: begin
            cosine_reg0 <= 36'sb111011100110001001110110101111110100;
            sine_reg0   <= 36'sb11111101100100000110111000110011111;
        end
        4457: begin
            cosine_reg0 <= 36'sb111011100101011000000100011100110110;
            sine_reg0   <= 36'sb11111101100011001111011110001001001;
        end
        4458: begin
            cosine_reg0 <= 36'sb111011100100100110010010010100110001;
            sine_reg0   <= 36'sb11111101100010010111111001101100101;
        end
        4459: begin
            cosine_reg0 <= 36'sb111011100011110100100000010111100111;
            sine_reg0   <= 36'sb11111101100001100000001011011110101;
        end
        4460: begin
            cosine_reg0 <= 36'sb111011100011000010101110100101011010;
            sine_reg0   <= 36'sb11111101100000101000010011011111001;
        end
        4461: begin
            cosine_reg0 <= 36'sb111011100010010000111100111110001100;
            sine_reg0   <= 36'sb11111101011111110000010001101110000;
        end
        4462: begin
            cosine_reg0 <= 36'sb111011100001011111001011100010000000;
            sine_reg0   <= 36'sb11111101011110111000000110001011100;
        end
        4463: begin
            cosine_reg0 <= 36'sb111011100000101101011010010000110110;
            sine_reg0   <= 36'sb11111101011101111111110000110111100;
        end
        4464: begin
            cosine_reg0 <= 36'sb111011011111111011101001001010110001;
            sine_reg0   <= 36'sb11111101011101000111010001110010001;
        end
        4465: begin
            cosine_reg0 <= 36'sb111011011111001001111000001111110011;
            sine_reg0   <= 36'sb11111101011100001110101000111011011;
        end
        4466: begin
            cosine_reg0 <= 36'sb111011011110011000000111011111111110;
            sine_reg0   <= 36'sb11111101011011010101110110010011010;
        end
        4467: begin
            cosine_reg0 <= 36'sb111011011101100110010110111011010011;
            sine_reg0   <= 36'sb11111101011010011100111001111001110;
        end
        4468: begin
            cosine_reg0 <= 36'sb111011011100110100100110100001110101;
            sine_reg0   <= 36'sb11111101011001100011110011101111001;
        end
        4469: begin
            cosine_reg0 <= 36'sb111011011100000010110110010011100110;
            sine_reg0   <= 36'sb11111101011000101010100011110011001;
        end
        4470: begin
            cosine_reg0 <= 36'sb111011011011010001000110010000100110;
            sine_reg0   <= 36'sb11111101010111110001001010000110000;
        end
        4471: begin
            cosine_reg0 <= 36'sb111011011010011111010110011000111001;
            sine_reg0   <= 36'sb11111101010110110111100110100111110;
        end
        4472: begin
            cosine_reg0 <= 36'sb111011011001101101100110101100100000;
            sine_reg0   <= 36'sb11111101010101111101111001011000010;
        end
        4473: begin
            cosine_reg0 <= 36'sb111011011000111011110111001011011110;
            sine_reg0   <= 36'sb11111101010101000100000010010111110;
        end
        4474: begin
            cosine_reg0 <= 36'sb111011011000001010000111110101110011;
            sine_reg0   <= 36'sb11111101010100001010000001100110001;
        end
        4475: begin
            cosine_reg0 <= 36'sb111011010111011000011000101011100010;
            sine_reg0   <= 36'sb11111101010011001111110111000011100;
        end
        4476: begin
            cosine_reg0 <= 36'sb111011010110100110101001101100101101;
            sine_reg0   <= 36'sb11111101010010010101100010101111111;
        end
        4477: begin
            cosine_reg0 <= 36'sb111011010101110100111010111001010110;
            sine_reg0   <= 36'sb11111101010001011011000100101011010;
        end
        4478: begin
            cosine_reg0 <= 36'sb111011010101000011001100010001011111;
            sine_reg0   <= 36'sb11111101010000100000011100110101110;
        end
        4479: begin
            cosine_reg0 <= 36'sb111011010100010001011101110101001001;
            sine_reg0   <= 36'sb11111101001111100101101011001111011;
        end
        4480: begin
            cosine_reg0 <= 36'sb111011010011011111101111100100010111;
            sine_reg0   <= 36'sb11111101001110101010101111111000001;
        end
        4481: begin
            cosine_reg0 <= 36'sb111011010010101110000001011111001011;
            sine_reg0   <= 36'sb11111101001101101111101010110000001;
        end
        4482: begin
            cosine_reg0 <= 36'sb111011010001111100010011100101100101;
            sine_reg0   <= 36'sb11111101001100110100011011110111010;
        end
        4483: begin
            cosine_reg0 <= 36'sb111011010001001010100101110111101001;
            sine_reg0   <= 36'sb11111101001011111001000011001101101;
        end
        4484: begin
            cosine_reg0 <= 36'sb111011010000011000111000010101011000;
            sine_reg0   <= 36'sb11111101001010111101100000110011011;
        end
        4485: begin
            cosine_reg0 <= 36'sb111011001111100111001010111110110101;
            sine_reg0   <= 36'sb11111101001010000001110100101000011;
        end
        4486: begin
            cosine_reg0 <= 36'sb111011001110110101011101110100000000;
            sine_reg0   <= 36'sb11111101001001000101111110101100110;
        end
        4487: begin
            cosine_reg0 <= 36'sb111011001110000011110000110100111101;
            sine_reg0   <= 36'sb11111101001000001001111111000000100;
        end
        4488: begin
            cosine_reg0 <= 36'sb111011001101010010000100000001101100;
            sine_reg0   <= 36'sb11111101000111001101110101100011110;
        end
        4489: begin
            cosine_reg0 <= 36'sb111011001100100000010111011010010000;
            sine_reg0   <= 36'sb11111101000110010001100010010110011;
        end
        4490: begin
            cosine_reg0 <= 36'sb111011001011101110101010111110101011;
            sine_reg0   <= 36'sb11111101000101010101000101011000100;
        end
        4491: begin
            cosine_reg0 <= 36'sb111011001010111100111110101110111110;
            sine_reg0   <= 36'sb11111101000100011000011110101010010;
        end
        4492: begin
            cosine_reg0 <= 36'sb111011001010001011010010101011001100;
            sine_reg0   <= 36'sb11111101000011011011101110001011101;
        end
        4493: begin
            cosine_reg0 <= 36'sb111011001001011001100110110011010110;
            sine_reg0   <= 36'sb11111101000010011110110011111100100;
        end
        4494: begin
            cosine_reg0 <= 36'sb111011001000100111111011000111011111;
            sine_reg0   <= 36'sb11111101000001100001101111111101001;
        end
        4495: begin
            cosine_reg0 <= 36'sb111011000111110110001111100111101000;
            sine_reg0   <= 36'sb11111101000000100100100010001101011;
        end
        4496: begin
            cosine_reg0 <= 36'sb111011000111000100100100010011110011;
            sine_reg0   <= 36'sb11111100111111100111001010101101010;
        end
        4497: begin
            cosine_reg0 <= 36'sb111011000110010010111001001100000011;
            sine_reg0   <= 36'sb11111100111110101001101001011101000;
        end
        4498: begin
            cosine_reg0 <= 36'sb111011000101100001001110010000011000;
            sine_reg0   <= 36'sb11111100111101101011111110011100101;
        end
        4499: begin
            cosine_reg0 <= 36'sb111011000100101111100011100000110101;
            sine_reg0   <= 36'sb11111100111100101110001001101100000;
        end
        4500: begin
            cosine_reg0 <= 36'sb111011000011111101111000111101011101;
            sine_reg0   <= 36'sb11111100111011110000001011001011010;
        end
        4501: begin
            cosine_reg0 <= 36'sb111011000011001100001110100110010000;
            sine_reg0   <= 36'sb11111100111010110010000010111010011;
        end
        4502: begin
            cosine_reg0 <= 36'sb111011000010011010100100011011010000;
            sine_reg0   <= 36'sb11111100111001110011110000111001100;
        end
        4503: begin
            cosine_reg0 <= 36'sb111011000001101000111010011100100001;
            sine_reg0   <= 36'sb11111100111000110101010101001000101;
        end
        4504: begin
            cosine_reg0 <= 36'sb111011000000110111010000101010000010;
            sine_reg0   <= 36'sb11111100110111110110101111100111110;
        end
        4505: begin
            cosine_reg0 <= 36'sb111011000000000101100111000011111000;
            sine_reg0   <= 36'sb11111100110110111000000000010110111;
        end
        4506: begin
            cosine_reg0 <= 36'sb111010111111010011111101101010000010;
            sine_reg0   <= 36'sb11111100110101111001000111010110010;
        end
        4507: begin
            cosine_reg0 <= 36'sb111010111110100010010100011100100100;
            sine_reg0   <= 36'sb11111100110100111010000100100101101;
        end
        4508: begin
            cosine_reg0 <= 36'sb111010111101110000101011011011011111;
            sine_reg0   <= 36'sb11111100110011111010111000000101010;
        end
        4509: begin
            cosine_reg0 <= 36'sb111010111100111111000010100110110101;
            sine_reg0   <= 36'sb11111100110010111011100001110101000;
        end
        4510: begin
            cosine_reg0 <= 36'sb111010111100001101011001111110101001;
            sine_reg0   <= 36'sb11111100110001111100000001110101001;
        end
        4511: begin
            cosine_reg0 <= 36'sb111010111011011011110001100010111011;
            sine_reg0   <= 36'sb11111100110000111100011000000101100;
        end
        4512: begin
            cosine_reg0 <= 36'sb111010111010101010001001010011101110;
            sine_reg0   <= 36'sb11111100101111111100100100100110001;
        end
        4513: begin
            cosine_reg0 <= 36'sb111010111001111000100001010001000011;
            sine_reg0   <= 36'sb11111100101110111100100111010111010;
        end
        4514: begin
            cosine_reg0 <= 36'sb111010111001000110111001011010111110;
            sine_reg0   <= 36'sb11111100101101111100100000011000101;
        end
        4515: begin
            cosine_reg0 <= 36'sb111010111000010101010001110001011110;
            sine_reg0   <= 36'sb11111100101100111100001111101010100;
        end
        4516: begin
            cosine_reg0 <= 36'sb111010110111100011101010010100101000;
            sine_reg0   <= 36'sb11111100101011111011110101001100111;
        end
        4517: begin
            cosine_reg0 <= 36'sb111010110110110010000011000100011100;
            sine_reg0   <= 36'sb11111100101010111011010000111111111;
        end
        4518: begin
            cosine_reg0 <= 36'sb111010110110000000011100000000111100;
            sine_reg0   <= 36'sb11111100101001111010100011000011010;
        end
        4519: begin
            cosine_reg0 <= 36'sb111010110101001110110101001010001010;
            sine_reg0   <= 36'sb11111100101000111001101011010111011;
        end
        4520: begin
            cosine_reg0 <= 36'sb111010110100011101001110100000001001;
            sine_reg0   <= 36'sb11111100100111111000101001111100000;
        end
        4521: begin
            cosine_reg0 <= 36'sb111010110011101011101000000010111001;
            sine_reg0   <= 36'sb11111100100110110111011110110001011;
        end
        4522: begin
            cosine_reg0 <= 36'sb111010110010111010000001110010011110;
            sine_reg0   <= 36'sb11111100100101110110001001110111100;
        end
        4523: begin
            cosine_reg0 <= 36'sb111010110010001000011011101110111000;
            sine_reg0   <= 36'sb11111100100100110100101011001110011;
        end
        4524: begin
            cosine_reg0 <= 36'sb111010110001010110110101111000001010;
            sine_reg0   <= 36'sb11111100100011110011000010110110000;
        end
        4525: begin
            cosine_reg0 <= 36'sb111010110000100101010000001110010110;
            sine_reg0   <= 36'sb11111100100010110001010000101110100;
        end
        4526: begin
            cosine_reg0 <= 36'sb111010101111110011101010110001011101;
            sine_reg0   <= 36'sb11111100100001101111010100110111111;
        end
        4527: begin
            cosine_reg0 <= 36'sb111010101111000010000101100001100010;
            sine_reg0   <= 36'sb11111100100000101101001111010010001;
        end
        4528: begin
            cosine_reg0 <= 36'sb111010101110010000100000011110100111;
            sine_reg0   <= 36'sb11111100011111101010111111111101011;
        end
        4529: begin
            cosine_reg0 <= 36'sb111010101101011110111011101000101100;
            sine_reg0   <= 36'sb11111100011110101000100110111001100;
        end
        4530: begin
            cosine_reg0 <= 36'sb111010101100101101010110111111110101;
            sine_reg0   <= 36'sb11111100011101100110000100000110110;
        end
        4531: begin
            cosine_reg0 <= 36'sb111010101011111011110010100100000100;
            sine_reg0   <= 36'sb11111100011100100011010111100101001;
        end
        4532: begin
            cosine_reg0 <= 36'sb111010101011001010001110010101011001;
            sine_reg0   <= 36'sb11111100011011100000100001010100100;
        end
        4533: begin
            cosine_reg0 <= 36'sb111010101010011000101010010011110111;
            sine_reg0   <= 36'sb11111100011010011101100001010101001;
        end
        4534: begin
            cosine_reg0 <= 36'sb111010101001100111000110011111100000;
            sine_reg0   <= 36'sb11111100011001011010010111100110111;
        end
        4535: begin
            cosine_reg0 <= 36'sb111010101000110101100010111000010110;
            sine_reg0   <= 36'sb11111100011000010111000100001001111;
        end
        4536: begin
            cosine_reg0 <= 36'sb111010101000000011111111011110011011;
            sine_reg0   <= 36'sb11111100010111010011100110111110010;
        end
        4537: begin
            cosine_reg0 <= 36'sb111010100111010010011100010001110000;
            sine_reg0   <= 36'sb11111100010110010000000000000011111;
        end
        4538: begin
            cosine_reg0 <= 36'sb111010100110100000111001010010011000;
            sine_reg0   <= 36'sb11111100010101001100001111011010110;
        end
        4539: begin
            cosine_reg0 <= 36'sb111010100101101111010110100000010100;
            sine_reg0   <= 36'sb11111100010100001000010101000011001;
        end
        4540: begin
            cosine_reg0 <= 36'sb111010100100111101110011111011100111;
            sine_reg0   <= 36'sb11111100010011000100010000111101000;
        end
        4541: begin
            cosine_reg0 <= 36'sb111010100100001100010001100100010010;
            sine_reg0   <= 36'sb11111100010010000000000011001000010;
        end
        4542: begin
            cosine_reg0 <= 36'sb111010100011011010101111011010010111;
            sine_reg0   <= 36'sb11111100010000111011101011100101001;
        end
        4543: begin
            cosine_reg0 <= 36'sb111010100010101001001101011101111000;
            sine_reg0   <= 36'sb11111100001111110111001010010011100;
        end
        4544: begin
            cosine_reg0 <= 36'sb111010100001110111101011101110110111;
            sine_reg0   <= 36'sb11111100001110110010011111010011011;
        end
        4545: begin
            cosine_reg0 <= 36'sb111010100001000110001010001101010111;
            sine_reg0   <= 36'sb11111100001101101101101010100101000;
        end
        4546: begin
            cosine_reg0 <= 36'sb111010100000010100101000111001011000;
            sine_reg0   <= 36'sb11111100001100101000101100001000011;
        end
        4547: begin
            cosine_reg0 <= 36'sb111010011111100011000111110010111100;
            sine_reg0   <= 36'sb11111100001011100011100011111101011;
        end
        4548: begin
            cosine_reg0 <= 36'sb111010011110110001100110111010000111;
            sine_reg0   <= 36'sb11111100001010011110010010000100001;
        end
        4549: begin
            cosine_reg0 <= 36'sb111010011110000000000110001110111000;
            sine_reg0   <= 36'sb11111100001001011000110110011100110;
        end
        4550: begin
            cosine_reg0 <= 36'sb111010011101001110100101110001010100;
            sine_reg0   <= 36'sb11111100001000010011010001000111010;
        end
        4551: begin
            cosine_reg0 <= 36'sb111010011100011101000101100001011010;
            sine_reg0   <= 36'sb11111100000111001101100010000011101;
        end
        4552: begin
            cosine_reg0 <= 36'sb111010011011101011100101011111001110;
            sine_reg0   <= 36'sb11111100000110000111101001010001111;
        end
        4553: begin
            cosine_reg0 <= 36'sb111010011010111010000101101010110001;
            sine_reg0   <= 36'sb11111100000101000001100110110010001;
        end
        4554: begin
            cosine_reg0 <= 36'sb111010011010001000100110000100000110;
            sine_reg0   <= 36'sb11111100000011111011011010100100100;
        end
        4555: begin
            cosine_reg0 <= 36'sb111010011001010111000110101011001101;
            sine_reg0   <= 36'sb11111100000010110101000100101000111;
        end
        4556: begin
            cosine_reg0 <= 36'sb111010011000100101100111100000001001;
            sine_reg0   <= 36'sb11111100000001101110100100111111010;
        end
        4557: begin
            cosine_reg0 <= 36'sb111010010111110100001000100010111100;
            sine_reg0   <= 36'sb11111100000000100111111011100111111;
        end
        4558: begin
            cosine_reg0 <= 36'sb111010010111000010101001110011101000;
            sine_reg0   <= 36'sb11111011111111100001001000100010110;
        end
        4559: begin
            cosine_reg0 <= 36'sb111010010110010001001011010010001110;
            sine_reg0   <= 36'sb11111011111110011010001011101111110;
        end
        4560: begin
            cosine_reg0 <= 36'sb111010010101011111101100111110110001;
            sine_reg0   <= 36'sb11111011111101010011000101001111001;
        end
        4561: begin
            cosine_reg0 <= 36'sb111010010100101110001110111001010010;
            sine_reg0   <= 36'sb11111011111100001011110101000000110;
        end
        4562: begin
            cosine_reg0 <= 36'sb111010010011111100110001000001110100;
            sine_reg0   <= 36'sb11111011111011000100011011000100110;
        end
        4563: begin
            cosine_reg0 <= 36'sb111010010011001011010011011000011000;
            sine_reg0   <= 36'sb11111011111001111100110111011011001;
        end
        4564: begin
            cosine_reg0 <= 36'sb111010010010011001110101111101000000;
            sine_reg0   <= 36'sb11111011111000110101001010000100000;
        end
        4565: begin
            cosine_reg0 <= 36'sb111010010001101000011000101111101110;
            sine_reg0   <= 36'sb11111011110111101101010010111111010;
        end
        4566: begin
            cosine_reg0 <= 36'sb111010010000110110111011110000100100;
            sine_reg0   <= 36'sb11111011110110100101010010001101001;
        end
        4567: begin
            cosine_reg0 <= 36'sb111010010000000101011110111111100100;
            sine_reg0   <= 36'sb11111011110101011101000111101101101;
        end
        4568: begin
            cosine_reg0 <= 36'sb111010001111010100000010011100110000;
            sine_reg0   <= 36'sb11111011110100010100110011100000110;
        end
        4569: begin
            cosine_reg0 <= 36'sb111010001110100010100110001000001001;
            sine_reg0   <= 36'sb11111011110011001100010101100110011;
        end
        4570: begin
            cosine_reg0 <= 36'sb111010001101110001001010000001110010;
            sine_reg0   <= 36'sb11111011110010000011101101111110111;
        end
        4571: begin
            cosine_reg0 <= 36'sb111010001100111111101110001001101101;
            sine_reg0   <= 36'sb11111011110000111010111100101010001;
        end
        4572: begin
            cosine_reg0 <= 36'sb111010001100001110010010011111111011;
            sine_reg0   <= 36'sb11111011101111110010000001101000001;
        end
        4573: begin
            cosine_reg0 <= 36'sb111010001011011100110111000100011110;
            sine_reg0   <= 36'sb11111011101110101000111100111000111;
        end
        4574: begin
            cosine_reg0 <= 36'sb111010001010101011011011110111011001;
            sine_reg0   <= 36'sb11111011101101011111101110011100101;
        end
        4575: begin
            cosine_reg0 <= 36'sb111010001001111010000000111000101100;
            sine_reg0   <= 36'sb11111011101100010110010110010011010;
        end
        4576: begin
            cosine_reg0 <= 36'sb111010001001001000100110001000011011;
            sine_reg0   <= 36'sb11111011101011001100110100011100111;
        end
        4577: begin
            cosine_reg0 <= 36'sb111010001000010111001011100110100111;
            sine_reg0   <= 36'sb11111011101010000011001000111001100;
        end
        4578: begin
            cosine_reg0 <= 36'sb111010000111100101110001010011010001;
            sine_reg0   <= 36'sb11111011101000111001010011101001010;
        end
        4579: begin
            cosine_reg0 <= 36'sb111010000110110100010111001110011101;
            sine_reg0   <= 36'sb11111011100111101111010100101100000;
        end
        4580: begin
            cosine_reg0 <= 36'sb111010000110000010111101011000001011;
            sine_reg0   <= 36'sb11111011100110100101001100000010000;
        end
        4581: begin
            cosine_reg0 <= 36'sb111010000101010001100011110000011101;
            sine_reg0   <= 36'sb11111011100101011010111001101011001;
        end
        4582: begin
            cosine_reg0 <= 36'sb111010000100100000001010010111010110;
            sine_reg0   <= 36'sb11111011100100010000011101100111100;
        end
        4583: begin
            cosine_reg0 <= 36'sb111010000011101110110001001100110111;
            sine_reg0   <= 36'sb11111011100011000101110111110111010;
        end
        4584: begin
            cosine_reg0 <= 36'sb111010000010111101011000010001000011;
            sine_reg0   <= 36'sb11111011100001111011001000011010010;
        end
        4585: begin
            cosine_reg0 <= 36'sb111010000010001011111111100011111011;
            sine_reg0   <= 36'sb11111011100000110000001111010000101;
        end
        4586: begin
            cosine_reg0 <= 36'sb111010000001011010100111000101100001;
            sine_reg0   <= 36'sb11111011011111100101001100011010011;
        end
        4587: begin
            cosine_reg0 <= 36'sb111010000000101001001110110101110111;
            sine_reg0   <= 36'sb11111011011110011001111111110111101;
        end
        4588: begin
            cosine_reg0 <= 36'sb111001111111110111110110110100111110;
            sine_reg0   <= 36'sb11111011011101001110101001101000100;
        end
        4589: begin
            cosine_reg0 <= 36'sb111001111111000110011111000010111010;
            sine_reg0   <= 36'sb11111011011100000011001001101100110;
        end
        4590: begin
            cosine_reg0 <= 36'sb111001111110010101000111011111101011;
            sine_reg0   <= 36'sb11111011011010110111100000000100110;
        end
        4591: begin
            cosine_reg0 <= 36'sb111001111101100011110000001011010100;
            sine_reg0   <= 36'sb11111011011001101011101100110000010;
        end
        4592: begin
            cosine_reg0 <= 36'sb111001111100110010011001000101110110;
            sine_reg0   <= 36'sb11111011011000011111101111101111100;
        end
        4593: begin
            cosine_reg0 <= 36'sb111001111100000001000010001111010100;
            sine_reg0   <= 36'sb11111011010111010011101001000010101;
        end
        4594: begin
            cosine_reg0 <= 36'sb111001111011001111101011100111101111;
            sine_reg0   <= 36'sb11111011010110000111011000101001011;
        end
        4595: begin
            cosine_reg0 <= 36'sb111001111010011110010101001111001010;
            sine_reg0   <= 36'sb11111011010100111010111110100100000;
        end
        4596: begin
            cosine_reg0 <= 36'sb111001111001101100111111000101100101;
            sine_reg0   <= 36'sb11111011010011101110011010110010100;
        end
        4597: begin
            cosine_reg0 <= 36'sb111001111000111011101001001011000011;
            sine_reg0   <= 36'sb11111011010010100001101101010100111;
        end
        4598: begin
            cosine_reg0 <= 36'sb111001111000001010010011011111100111;
            sine_reg0   <= 36'sb11111011010001010100110110001011010;
        end
        4599: begin
            cosine_reg0 <= 36'sb111001110111011000111110000011010001;
            sine_reg0   <= 36'sb11111011010000000111110101010101101;
        end
        4600: begin
            cosine_reg0 <= 36'sb111001110110100111101000110110000100;
            sine_reg0   <= 36'sb11111011001110111010101010110100001;
        end
        4601: begin
            cosine_reg0 <= 36'sb111001110101110110010011111000000001;
            sine_reg0   <= 36'sb11111011001101101101010110100110110;
        end
        4602: begin
            cosine_reg0 <= 36'sb111001110101000100111111001001001100;
            sine_reg0   <= 36'sb11111011001100011111111000101101011;
        end
        4603: begin
            cosine_reg0 <= 36'sb111001110100010011101010101001100100;
            sine_reg0   <= 36'sb11111011001011010010010001001000011;
        end
        4604: begin
            cosine_reg0 <= 36'sb111001110011100010010110011001001101;
            sine_reg0   <= 36'sb11111011001010000100011111110111100;
        end
        4605: begin
            cosine_reg0 <= 36'sb111001110010110001000010011000001000;
            sine_reg0   <= 36'sb11111011001000110110100100111011000;
        end
        4606: begin
            cosine_reg0 <= 36'sb111001110001111111101110100110010111;
            sine_reg0   <= 36'sb11111011000111101000100000010010110;
        end
        4607: begin
            cosine_reg0 <= 36'sb111001110001001110011011000011111100;
            sine_reg0   <= 36'sb11111011000110011010010001111111000;
        end
        4608: begin
            cosine_reg0 <= 36'sb111001110000011101000111110000111010;
            sine_reg0   <= 36'sb11111011000101001011111001111111101;
        end
        4609: begin
            cosine_reg0 <= 36'sb111001101111101011110100101101010001;
            sine_reg0   <= 36'sb11111011000011111101011000010100110;
        end
        4610: begin
            cosine_reg0 <= 36'sb111001101110111010100001111001000011;
            sine_reg0   <= 36'sb11111011000010101110101100111110011;
        end
        4611: begin
            cosine_reg0 <= 36'sb111001101110001001001111010100010100;
            sine_reg0   <= 36'sb11111011000001011111110111111100101;
        end
        4612: begin
            cosine_reg0 <= 36'sb111001101101010111111100111111000100;
            sine_reg0   <= 36'sb11111011000000010000111001001111011;
        end
        4613: begin
            cosine_reg0 <= 36'sb111001101100100110101010111001010101;
            sine_reg0   <= 36'sb11111010111111000001110000110110111;
        end
        4614: begin
            cosine_reg0 <= 36'sb111001101011110101011001000011001010;
            sine_reg0   <= 36'sb11111010111101110010011110110011001;
        end
        4615: begin
            cosine_reg0 <= 36'sb111001101011000100000111011100100100;
            sine_reg0   <= 36'sb11111010111100100011000011000100001;
        end
        4616: begin
            cosine_reg0 <= 36'sb111001101010010010110110000101100101;
            sine_reg0   <= 36'sb11111010111011010011011101101010000;
        end
        4617: begin
            cosine_reg0 <= 36'sb111001101001100001100100111110001111;
            sine_reg0   <= 36'sb11111010111010000011101110100100101;
        end
        4618: begin
            cosine_reg0 <= 36'sb111001101000110000010100000110100100;
            sine_reg0   <= 36'sb11111010111000110011110101110100010;
        end
        4619: begin
            cosine_reg0 <= 36'sb111001100111111111000011011110100110;
            sine_reg0   <= 36'sb11111010110111100011110011011000110;
        end
        4620: begin
            cosine_reg0 <= 36'sb111001100111001101110011000110010111;
            sine_reg0   <= 36'sb11111010110110010011100111010010011;
        end
        4621: begin
            cosine_reg0 <= 36'sb111001100110011100100010111101111000;
            sine_reg0   <= 36'sb11111010110101000011010001100001000;
        end
        4622: begin
            cosine_reg0 <= 36'sb111001100101101011010011000101001100;
            sine_reg0   <= 36'sb11111010110011110010110010000100110;
        end
        4623: begin
            cosine_reg0 <= 36'sb111001100100111010000011011100010100;
            sine_reg0   <= 36'sb11111010110010100010001000111101101;
        end
        4624: begin
            cosine_reg0 <= 36'sb111001100100001000110100000011010010;
            sine_reg0   <= 36'sb11111010110001010001010110001011101;
        end
        4625: begin
            cosine_reg0 <= 36'sb111001100011010111100100111010001001;
            sine_reg0   <= 36'sb11111010110000000000011001101111000;
        end
        4626: begin
            cosine_reg0 <= 36'sb111001100010100110010110000000111010;
            sine_reg0   <= 36'sb11111010101110101111010011100111101;
        end
        4627: begin
            cosine_reg0 <= 36'sb111001100001110101000111010111100111;
            sine_reg0   <= 36'sb11111010101101011110000011110101101;
        end
        4628: begin
            cosine_reg0 <= 36'sb111001100001000011111000111110010010;
            sine_reg0   <= 36'sb11111010101100001100101010011000111;
        end
        4629: begin
            cosine_reg0 <= 36'sb111001100000010010101010110100111101;
            sine_reg0   <= 36'sb11111010101010111011000111010001110;
        end
        4630: begin
            cosine_reg0 <= 36'sb111001011111100001011100111011101001;
            sine_reg0   <= 36'sb11111010101001101001011010100000000;
        end
        4631: begin
            cosine_reg0 <= 36'sb111001011110110000001111010010011001;
            sine_reg0   <= 36'sb11111010101000010111100100000011111;
        end
        4632: begin
            cosine_reg0 <= 36'sb111001011101111111000001111001001111;
            sine_reg0   <= 36'sb11111010100111000101100011111101011;
        end
        4633: begin
            cosine_reg0 <= 36'sb111001011101001101110100110000001100;
            sine_reg0   <= 36'sb11111010100101110011011010001100100;
        end
        4634: begin
            cosine_reg0 <= 36'sb111001011100011100100111110111010010;
            sine_reg0   <= 36'sb11111010100100100001000110110001010;
        end
        4635: begin
            cosine_reg0 <= 36'sb111001011011101011011011001110100011;
            sine_reg0   <= 36'sb11111010100011001110101001101011110;
        end
        4636: begin
            cosine_reg0 <= 36'sb111001011010111010001110110110000010;
            sine_reg0   <= 36'sb11111010100001111100000010111100000;
        end
        4637: begin
            cosine_reg0 <= 36'sb111001011010001001000010101101110000;
            sine_reg0   <= 36'sb11111010100000101001010010100010010;
        end
        4638: begin
            cosine_reg0 <= 36'sb111001011001010111110110110101101110;
            sine_reg0   <= 36'sb11111010011111010110011000011110010;
        end
        4639: begin
            cosine_reg0 <= 36'sb111001011000100110101011001101111111;
            sine_reg0   <= 36'sb11111010011110000011010100110000010;
        end
        4640: begin
            cosine_reg0 <= 36'sb111001010111110101011111110110100101;
            sine_reg0   <= 36'sb11111010011100110000000111011000010;
        end
        4641: begin
            cosine_reg0 <= 36'sb111001010111000100010100101111100010;
            sine_reg0   <= 36'sb11111010011011011100110000010110010;
        end
        4642: begin
            cosine_reg0 <= 36'sb111001010110010011001001111000110111;
            sine_reg0   <= 36'sb11111010011010001001001111101010011;
        end
        4643: begin
            cosine_reg0 <= 36'sb111001010101100001111111010010100110;
            sine_reg0   <= 36'sb11111010011000110101100101010100101;
        end
        4644: begin
            cosine_reg0 <= 36'sb111001010100110000110100111100110010;
            sine_reg0   <= 36'sb11111010010111100001110001010101000;
        end
        4645: begin
            cosine_reg0 <= 36'sb111001010011111111101010110111011100;
            sine_reg0   <= 36'sb11111010010110001101110011101011110;
        end
        4646: begin
            cosine_reg0 <= 36'sb111001010011001110100001000010100101;
            sine_reg0   <= 36'sb11111010010100111001101100011000110;
        end
        4647: begin
            cosine_reg0 <= 36'sb111001010010011101010111011110010001;
            sine_reg0   <= 36'sb11111010010011100101011011011100000;
        end
        4648: begin
            cosine_reg0 <= 36'sb111001010001101100001110001010100001;
            sine_reg0   <= 36'sb11111010010010010001000000110101110;
        end
        4649: begin
            cosine_reg0 <= 36'sb111001010000111011000101000111010110;
            sine_reg0   <= 36'sb11111010010000111100011100100110000;
        end
        4650: begin
            cosine_reg0 <= 36'sb111001010000001001111100010100110011;
            sine_reg0   <= 36'sb11111010001111100111101110101100101;
        end
        4651: begin
            cosine_reg0 <= 36'sb111001001111011000110011110010111010;
            sine_reg0   <= 36'sb11111010001110010010110111001001110;
        end
        4652: begin
            cosine_reg0 <= 36'sb111001001110100111101011100001101100;
            sine_reg0   <= 36'sb11111010001100111101110101111101101;
        end
        4653: begin
            cosine_reg0 <= 36'sb111001001101110110100011100001001011;
            sine_reg0   <= 36'sb11111010001011101000101011001000001;
        end
        4654: begin
            cosine_reg0 <= 36'sb111001001101000101011011110001011010;
            sine_reg0   <= 36'sb11111010001010010011010110101001010;
        end
        4655: begin
            cosine_reg0 <= 36'sb111001001100010100010100010010011010;
            sine_reg0   <= 36'sb11111010001000111101111000100001001;
        end
        4656: begin
            cosine_reg0 <= 36'sb111001001011100011001101000100001100;
            sine_reg0   <= 36'sb11111010000111101000010000101111111;
        end
        4657: begin
            cosine_reg0 <= 36'sb111001001010110010000110000110110100;
            sine_reg0   <= 36'sb11111010000110010010011111010101011;
        end
        4658: begin
            cosine_reg0 <= 36'sb111001001010000000111111011010010010;
            sine_reg0   <= 36'sb11111010000100111100100100010001111;
        end
        4659: begin
            cosine_reg0 <= 36'sb111001001001001111111000111110101001;
            sine_reg0   <= 36'sb11111010000011100110011111100101011;
        end
        4660: begin
            cosine_reg0 <= 36'sb111001001000011110110010110011111011;
            sine_reg0   <= 36'sb11111010000010010000010001001111110;
        end
        4661: begin
            cosine_reg0 <= 36'sb111001000111101101101100111010001001;
            sine_reg0   <= 36'sb11111010000000111001111001010001011;
        end
        4662: begin
            cosine_reg0 <= 36'sb111001000110111100100111010001010110;
            sine_reg0   <= 36'sb11111001111111100011010111101010000;
        end
        4663: begin
            cosine_reg0 <= 36'sb111001000110001011100001111001100010;
            sine_reg0   <= 36'sb11111001111110001100101100011001110;
        end
        4664: begin
            cosine_reg0 <= 36'sb111001000101011010011100110010110001;
            sine_reg0   <= 36'sb11111001111100110101110111100000110;
        end
        4665: begin
            cosine_reg0 <= 36'sb111001000100101001010111111101000100;
            sine_reg0   <= 36'sb11111001111011011110111000111111000;
        end
        4666: begin
            cosine_reg0 <= 36'sb111001000011111000010011011000011101;
            sine_reg0   <= 36'sb11111001111010000111110000110100101;
        end
        4667: begin
            cosine_reg0 <= 36'sb111001000011000111001111000100111110;
            sine_reg0   <= 36'sb11111001111000110000011111000001101;
        end
        4668: begin
            cosine_reg0 <= 36'sb111001000010010110001011000010101000;
            sine_reg0   <= 36'sb11111001110111011001000011100110000;
        end
        4669: begin
            cosine_reg0 <= 36'sb111001000001100101000111010001011110;
            sine_reg0   <= 36'sb11111001110110000001011110100001111;
        end
        4670: begin
            cosine_reg0 <= 36'sb111001000000110100000011110001100001;
            sine_reg0   <= 36'sb11111001110100101001101111110101011;
        end
        4671: begin
            cosine_reg0 <= 36'sb111001000000000011000000100010110100;
            sine_reg0   <= 36'sb11111001110011010001110111100000011;
        end
        4672: begin
            cosine_reg0 <= 36'sb111000111111010001111101100101011000;
            sine_reg0   <= 36'sb11111001110001111001110101100011000;
        end
        4673: begin
            cosine_reg0 <= 36'sb111000111110100000111010111001010000;
            sine_reg0   <= 36'sb11111001110000100001101001111101011;
        end
        4674: begin
            cosine_reg0 <= 36'sb111000111101101111111000011110011100;
            sine_reg0   <= 36'sb11111001101111001001010100101111100;
        end
        4675: begin
            cosine_reg0 <= 36'sb111000111100111110110110010100111111;
            sine_reg0   <= 36'sb11111001101101110000110101111001011;
        end
        4676: begin
            cosine_reg0 <= 36'sb111000111100001101110100011100111011;
            sine_reg0   <= 36'sb11111001101100011000001101011011001;
        end
        4677: begin
            cosine_reg0 <= 36'sb111000111011011100110010110110010010;
            sine_reg0   <= 36'sb11111001101010111111011011010100110;
        end
        4678: begin
            cosine_reg0 <= 36'sb111000111010101011110001100001000110;
            sine_reg0   <= 36'sb11111001101001100110011111100110011;
        end
        4679: begin
            cosine_reg0 <= 36'sb111000111001111010110000011101011000;
            sine_reg0   <= 36'sb11111001101000001101011010010000000;
        end
        4680: begin
            cosine_reg0 <= 36'sb111000111001001001101111101011001010;
            sine_reg0   <= 36'sb11111001100110110100001011010001110;
        end
        4681: begin
            cosine_reg0 <= 36'sb111000111000011000101111001010011111;
            sine_reg0   <= 36'sb11111001100101011010110010101011100;
        end
        4682: begin
            cosine_reg0 <= 36'sb111000110111100111101110111011011000;
            sine_reg0   <= 36'sb11111001100100000001010000011101100;
        end
        4683: begin
            cosine_reg0 <= 36'sb111000110110110110101110111101110111;
            sine_reg0   <= 36'sb11111001100010100111100100100111110;
        end
        4684: begin
            cosine_reg0 <= 36'sb111000110110000101101111010001111110;
            sine_reg0   <= 36'sb11111001100001001101101111001010010;
        end
        4685: begin
            cosine_reg0 <= 36'sb111000110101010100101111110111101111;
            sine_reg0   <= 36'sb11111001011111110011110000000101001;
        end
        4686: begin
            cosine_reg0 <= 36'sb111000110100100011110000101111001011;
            sine_reg0   <= 36'sb11111001011110011001100111011000010;
        end
        4687: begin
            cosine_reg0 <= 36'sb111000110011110010110001111000010101;
            sine_reg0   <= 36'sb11111001011100111111010101000100000;
        end
        4688: begin
            cosine_reg0 <= 36'sb111000110011000001110011010011001111;
            sine_reg0   <= 36'sb11111001011011100100111001001000001;
        end
        4689: begin
            cosine_reg0 <= 36'sb111000110010010000110100111111111010;
            sine_reg0   <= 36'sb11111001011010001010010011100100111;
        end
        4690: begin
            cosine_reg0 <= 36'sb111000110001011111110110111110011000;
            sine_reg0   <= 36'sb11111001011000101111100100011010010;
        end
        4691: begin
            cosine_reg0 <= 36'sb111000110000101110111001001110101100;
            sine_reg0   <= 36'sb11111001010111010100101011101000010;
        end
        4692: begin
            cosine_reg0 <= 36'sb111000101111111101111011110000110111;
            sine_reg0   <= 36'sb11111001010101111001101001001110111;
        end
        4693: begin
            cosine_reg0 <= 36'sb111000101111001100111110100100111010;
            sine_reg0   <= 36'sb11111001010100011110011101001110011;
        end
        4694: begin
            cosine_reg0 <= 36'sb111000101110011100000001101010111001;
            sine_reg0   <= 36'sb11111001010011000011000111100110110;
        end
        4695: begin
            cosine_reg0 <= 36'sb111000101101101011000101000010110100;
            sine_reg0   <= 36'sb11111001010001100111101000010111111;
        end
        4696: begin
            cosine_reg0 <= 36'sb111000101100111010001000101100101101;
            sine_reg0   <= 36'sb11111001010000001011111111100010001;
        end
        4697: begin
            cosine_reg0 <= 36'sb111000101100001001001100101000101000;
            sine_reg0   <= 36'sb11111001001110110000001101000101010;
        end
        4698: begin
            cosine_reg0 <= 36'sb111000101011011000010000110110100100;
            sine_reg0   <= 36'sb11111001001101010100010001000001011;
        end
        4699: begin
            cosine_reg0 <= 36'sb111000101010100111010101010110100101;
            sine_reg0   <= 36'sb11111001001011111000001011010110101;
        end
        4700: begin
            cosine_reg0 <= 36'sb111000101001110110011010001000101100;
            sine_reg0   <= 36'sb11111001001010011011111100000101001;
        end
        4701: begin
            cosine_reg0 <= 36'sb111000101001000101011111001100111011;
            sine_reg0   <= 36'sb11111001001000111111100011001100110;
        end
        4702: begin
            cosine_reg0 <= 36'sb111000101000010100100100100011010100;
            sine_reg0   <= 36'sb11111001000111100011000000101101101;
        end
        4703: begin
            cosine_reg0 <= 36'sb111000100111100011101010001011111001;
            sine_reg0   <= 36'sb11111001000110000110010100101000000;
        end
        4704: begin
            cosine_reg0 <= 36'sb111000100110110010110000000110101100;
            sine_reg0   <= 36'sb11111001000100101001011110111011101;
        end
        4705: begin
            cosine_reg0 <= 36'sb111000100110000001110110010011101110;
            sine_reg0   <= 36'sb11111001000011001100011111101000101;
        end
        4706: begin
            cosine_reg0 <= 36'sb111000100101010000111100110011000010;
            sine_reg0   <= 36'sb11111001000001101111010110101111010;
        end
        4707: begin
            cosine_reg0 <= 36'sb111000100100100000000011100100101001;
            sine_reg0   <= 36'sb11111001000000010010000100001111011;
        end
        4708: begin
            cosine_reg0 <= 36'sb111000100011101111001010101000100101;
            sine_reg0   <= 36'sb11111000111110110100101000001001000;
        end
        4709: begin
            cosine_reg0 <= 36'sb111000100010111110010001111110111000;
            sine_reg0   <= 36'sb11111000111101010111000010011100100;
        end
        4710: begin
            cosine_reg0 <= 36'sb111000100010001101011001100111100101;
            sine_reg0   <= 36'sb11111000111011111001010011001001100;
        end
        4711: begin
            cosine_reg0 <= 36'sb111000100001011100100001100010101100;
            sine_reg0   <= 36'sb11111000111010011011011010010000011;
        end
        4712: begin
            cosine_reg0 <= 36'sb111000100000101011101001110000010000;
            sine_reg0   <= 36'sb11111000111000111101010111110001001;
        end
        4713: begin
            cosine_reg0 <= 36'sb111000011111111010110010010000010011;
            sine_reg0   <= 36'sb11111000110111011111001011101011110;
        end
        4714: begin
            cosine_reg0 <= 36'sb111000011111001001111011000010110110;
            sine_reg0   <= 36'sb11111000110110000000110110000000010;
        end
        4715: begin
            cosine_reg0 <= 36'sb111000011110011001000100000111111100;
            sine_reg0   <= 36'sb11111000110100100010010110101110111;
        end
        4716: begin
            cosine_reg0 <= 36'sb111000011101101000001101011111100110;
            sine_reg0   <= 36'sb11111000110011000011101101110111100;
        end
        4717: begin
            cosine_reg0 <= 36'sb111000011100110111010111001001110110;
            sine_reg0   <= 36'sb11111000110001100100111011011010001;
        end
        4718: begin
            cosine_reg0 <= 36'sb111000011100000110100001000110101111;
            sine_reg0   <= 36'sb11111000110000000101111111010111000;
        end
        4719: begin
            cosine_reg0 <= 36'sb111000011011010101101011010110010001;
            sine_reg0   <= 36'sb11111000101110100110111001101110001;
        end
        4720: begin
            cosine_reg0 <= 36'sb111000011010100100110101111000011111;
            sine_reg0   <= 36'sb11111000101101000111101010011111101;
        end
        4721: begin
            cosine_reg0 <= 36'sb111000011001110100000000101101011011;
            sine_reg0   <= 36'sb11111000101011101000010001101011011;
        end
        4722: begin
            cosine_reg0 <= 36'sb111000011001000011001011110101000111;
            sine_reg0   <= 36'sb11111000101010001000101111010001100;
        end
        4723: begin
            cosine_reg0 <= 36'sb111000011000010010010111001111100100;
            sine_reg0   <= 36'sb11111000101000101001000011010010001;
        end
        4724: begin
            cosine_reg0 <= 36'sb111000010111100001100010111100110100;
            sine_reg0   <= 36'sb11111000100111001001001101101101010;
        end
        4725: begin
            cosine_reg0 <= 36'sb111000010110110000101110111100111010;
            sine_reg0   <= 36'sb11111000100101101001001110100011000;
        end
        4726: begin
            cosine_reg0 <= 36'sb111000010101111111111011001111110111;
            sine_reg0   <= 36'sb11111000100100001001000101110011011;
        end
        4727: begin
            cosine_reg0 <= 36'sb111000010101001111000111110101101101;
            sine_reg0   <= 36'sb11111000100010101000110011011110011;
        end
        4728: begin
            cosine_reg0 <= 36'sb111000010100011110010100101110011101;
            sine_reg0   <= 36'sb11111000100001001000010111100100001;
        end
        4729: begin
            cosine_reg0 <= 36'sb111000010011101101100001111010001011;
            sine_reg0   <= 36'sb11111000011111100111110010000100110;
        end
        4730: begin
            cosine_reg0 <= 36'sb111000010010111100101111011000110111;
            sine_reg0   <= 36'sb11111000011110000111000011000000010;
        end
        4731: begin
            cosine_reg0 <= 36'sb111000010010001011111101001010100100;
            sine_reg0   <= 36'sb11111000011100100110001010010110101;
        end
        4732: begin
            cosine_reg0 <= 36'sb111000010001011011001011001111010011;
            sine_reg0   <= 36'sb11111000011011000101001000001000000;
        end
        4733: begin
            cosine_reg0 <= 36'sb111000010000101010011001100111000111;
            sine_reg0   <= 36'sb11111000011001100011111100010100011;
        end
        4734: begin
            cosine_reg0 <= 36'sb111000001111111001101000010010000001;
            sine_reg0   <= 36'sb11111000011000000010100110111011111;
        end
        4735: begin
            cosine_reg0 <= 36'sb111000001111001000110111010000000010;
            sine_reg0   <= 36'sb11111000010110100001000111111110101;
        end
        4736: begin
            cosine_reg0 <= 36'sb111000001110011000000110100001001110;
            sine_reg0   <= 36'sb11111000010100111111011111011100100;
        end
        4737: begin
            cosine_reg0 <= 36'sb111000001101100111010110000101100110;
            sine_reg0   <= 36'sb11111000010011011101101101010101101;
        end
        4738: begin
            cosine_reg0 <= 36'sb111000001100110110100101111101001011;
            sine_reg0   <= 36'sb11111000010001111011110001101010001;
        end
        4739: begin
            cosine_reg0 <= 36'sb111000001100000101110110001000000000;
            sine_reg0   <= 36'sb11111000010000011001101100011010000;
        end
        4740: begin
            cosine_reg0 <= 36'sb111000001011010101000110100110000110;
            sine_reg0   <= 36'sb11111000001110110111011101100101011;
        end
        4741: begin
            cosine_reg0 <= 36'sb111000001010100100010111010111100000;
            sine_reg0   <= 36'sb11111000001101010101000101001100001;
        end
        4742: begin
            cosine_reg0 <= 36'sb111000001001110011101000011100001111;
            sine_reg0   <= 36'sb11111000001011110010100011001110101;
        end
        4743: begin
            cosine_reg0 <= 36'sb111000001001000010111001110100010101;
            sine_reg0   <= 36'sb11111000001010001111110111101100101;
        end
        4744: begin
            cosine_reg0 <= 36'sb111000001000010010001011011111110100;
            sine_reg0   <= 36'sb11111000001000101101000010100110011;
        end
        4745: begin
            cosine_reg0 <= 36'sb111000000111100001011101011110101110;
            sine_reg0   <= 36'sb11111000000111001010000011111011111;
        end
        4746: begin
            cosine_reg0 <= 36'sb111000000110110000101111110001000101;
            sine_reg0   <= 36'sb11111000000101100110111011101101001;
        end
        4747: begin
            cosine_reg0 <= 36'sb111000000110000000000010010110111010;
            sine_reg0   <= 36'sb11111000000100000011101001111010010;
        end
        4748: begin
            cosine_reg0 <= 36'sb111000000101001111010101010000010000;
            sine_reg0   <= 36'sb11111000000010100000001110100011011;
        end
        4749: begin
            cosine_reg0 <= 36'sb111000000100011110101000011101001001;
            sine_reg0   <= 36'sb11111000000000111100101001101000100;
        end
        4750: begin
            cosine_reg0 <= 36'sb111000000011101101111011111101100101;
            sine_reg0   <= 36'sb11110111111111011000111011001001101;
        end
        4751: begin
            cosine_reg0 <= 36'sb111000000010111101001111110001101000;
            sine_reg0   <= 36'sb11110111111101110101000011000110111;
        end
        4752: begin
            cosine_reg0 <= 36'sb111000000010001100100011111001010010;
            sine_reg0   <= 36'sb11110111111100010001000001100000010;
        end
        4753: begin
            cosine_reg0 <= 36'sb111000000001011011111000010100100111;
            sine_reg0   <= 36'sb11110111111010101100110110010101111;
        end
        4754: begin
            cosine_reg0 <= 36'sb111000000000101011001101000011100111;
            sine_reg0   <= 36'sb11110111111001001000100001100111110;
        end
        4755: begin
            cosine_reg0 <= 36'sb110111111111111010100010000110010101;
            sine_reg0   <= 36'sb11110111110111100100000011010110001;
        end
        4756: begin
            cosine_reg0 <= 36'sb110111111111001001110111011100110010;
            sine_reg0   <= 36'sb11110111110101111111011011100000110;
        end
        4757: begin
            cosine_reg0 <= 36'sb110111111110011001001101000111000001;
            sine_reg0   <= 36'sb11110111110100011010101010000111111;
        end
        4758: begin
            cosine_reg0 <= 36'sb110111111101101000100011000101000011;
            sine_reg0   <= 36'sb11110111110010110101101111001011101;
        end
        4759: begin
            cosine_reg0 <= 36'sb110111111100110111111001010110111011;
            sine_reg0   <= 36'sb11110111110001010000101010101011111;
        end
        4760: begin
            cosine_reg0 <= 36'sb110111111100000111001111111100101001;
            sine_reg0   <= 36'sb11110111101111101011011100101000110;
        end
        4761: begin
            cosine_reg0 <= 36'sb110111111011010110100110110110010000;
            sine_reg0   <= 36'sb11110111101110000110000101000010011;
        end
        4762: begin
            cosine_reg0 <= 36'sb110111111010100101111110000011110010;
            sine_reg0   <= 36'sb11110111101100100000100011111000111;
        end
        4763: begin
            cosine_reg0 <= 36'sb110111111001110101010101100101010001;
            sine_reg0   <= 36'sb11110111101010111010111001001100001;
        end
        4764: begin
            cosine_reg0 <= 36'sb110111111001000100101101011010101110;
            sine_reg0   <= 36'sb11110111101001010101000100111100010;
        end
        4765: begin
            cosine_reg0 <= 36'sb110111111000010100000101100100001011;
            sine_reg0   <= 36'sb11110111100111101111000111001001011;
        end
        4766: begin
            cosine_reg0 <= 36'sb110111110111100011011110000001101011;
            sine_reg0   <= 36'sb11110111100110001000111111110011100;
        end
        4767: begin
            cosine_reg0 <= 36'sb110111110110110010110110110011001111;
            sine_reg0   <= 36'sb11110111100100100010101110111010101;
        end
        4768: begin
            cosine_reg0 <= 36'sb110111110110000010001111111000111001;
            sine_reg0   <= 36'sb11110111100010111100010100011111000;
        end
        4769: begin
            cosine_reg0 <= 36'sb110111110101010001101001010010101011;
            sine_reg0   <= 36'sb11110111100001010101110000100000101;
        end
        4770: begin
            cosine_reg0 <= 36'sb110111110100100001000011000000100111;
            sine_reg0   <= 36'sb11110111011111101111000010111111011;
        end
        4771: begin
            cosine_reg0 <= 36'sb110111110011110000011101000010101110;
            sine_reg0   <= 36'sb11110111011110001000001011111011100;
        end
        4772: begin
            cosine_reg0 <= 36'sb110111110010111111110111011001000011;
            sine_reg0   <= 36'sb11110111011100100001001011010101001;
        end
        4773: begin
            cosine_reg0 <= 36'sb110111110010001111010010000011100111;
            sine_reg0   <= 36'sb11110111011010111010000001001100001;
        end
        4774: begin
            cosine_reg0 <= 36'sb110111110001011110101101000010011101;
            sine_reg0   <= 36'sb11110111011001010010101101100000101;
        end
        4775: begin
            cosine_reg0 <= 36'sb110111110000101110001000010101100101;
            sine_reg0   <= 36'sb11110111010111101011010000010010101;
        end
        4776: begin
            cosine_reg0 <= 36'sb110111101111111101100011111101000011;
            sine_reg0   <= 36'sb11110111010110000011101001100010011;
        end
        4777: begin
            cosine_reg0 <= 36'sb110111101111001100111111111000110111;
            sine_reg0   <= 36'sb11110111010100011011111001001111111;
        end
        4778: begin
            cosine_reg0 <= 36'sb110111101110011100011100001001000101;
            sine_reg0   <= 36'sb11110111010010110011111111011011000;
        end
        4779: begin
            cosine_reg0 <= 36'sb110111101101101011111000101101101100;
            sine_reg0   <= 36'sb11110111010001001011111100000100000;
        end
        4780: begin
            cosine_reg0 <= 36'sb110111101100111011010101100110110001;
            sine_reg0   <= 36'sb11110111001111100011101111001010111;
        end
        4781: begin
            cosine_reg0 <= 36'sb110111101100001010110010110100010100;
            sine_reg0   <= 36'sb11110111001101111011011000101111110;
        end
        4782: begin
            cosine_reg0 <= 36'sb110111101011011010010000010110010111;
            sine_reg0   <= 36'sb11110111001100010010111000110010101;
        end
        4783: begin
            cosine_reg0 <= 36'sb110111101010101001101110001100111100;
            sine_reg0   <= 36'sb11110111001010101010001111010011101;
        end
        4784: begin
            cosine_reg0 <= 36'sb110111101001111001001100011000000101;
            sine_reg0   <= 36'sb11110111001001000001011100010010110;
        end
        4785: begin
            cosine_reg0 <= 36'sb110111101001001000101010110111110100;
            sine_reg0   <= 36'sb11110111000111011000011111110000000;
        end
        4786: begin
            cosine_reg0 <= 36'sb110111101000011000001001101100001010;
            sine_reg0   <= 36'sb11110111000101101111011001101011101;
        end
        4787: begin
            cosine_reg0 <= 36'sb110111100111100111101000110101001011;
            sine_reg0   <= 36'sb11110111000100000110001010000101100;
        end
        4788: begin
            cosine_reg0 <= 36'sb110111100110110111001000010010110110;
            sine_reg0   <= 36'sb11110111000010011100110000111101110;
        end
        4789: begin
            cosine_reg0 <= 36'sb110111100110000110101000000101001111;
            sine_reg0   <= 36'sb11110111000000110011001110010100100;
        end
        4790: begin
            cosine_reg0 <= 36'sb110111100101010110001000001100011000;
            sine_reg0   <= 36'sb11110110111111001001100010001001110;
        end
        4791: begin
            cosine_reg0 <= 36'sb110111100100100101101000101000010001;
            sine_reg0   <= 36'sb11110110111101011111101100011101101;
        end
        4792: begin
            cosine_reg0 <= 36'sb110111100011110101001001011000111101;
            sine_reg0   <= 36'sb11110110111011110101101101010000001;
        end
        4793: begin
            cosine_reg0 <= 36'sb110111100011000100101010011110011110;
            sine_reg0   <= 36'sb11110110111010001011100100100001011;
        end
        4794: begin
            cosine_reg0 <= 36'sb110111100010010100001011111000110110;
            sine_reg0   <= 36'sb11110110111000100001010010010001011;
        end
        4795: begin
            cosine_reg0 <= 36'sb110111100001100011101101101000000111;
            sine_reg0   <= 36'sb11110110110110110110110110100000001;
        end
        4796: begin
            cosine_reg0 <= 36'sb110111100000110011001111101100010001;
            sine_reg0   <= 36'sb11110110110101001100010001001101111;
        end
        4797: begin
            cosine_reg0 <= 36'sb110111100000000010110010000101011000;
            sine_reg0   <= 36'sb11110110110011100001100010011010101;
        end
        4798: begin
            cosine_reg0 <= 36'sb110111011111010010010100110011011110;
            sine_reg0   <= 36'sb11110110110001110110101010000110011;
        end
        4799: begin
            cosine_reg0 <= 36'sb110111011110100001110111110110100011;
            sine_reg0   <= 36'sb11110110110000001011101000010001001;
        end
        4800: begin
            cosine_reg0 <= 36'sb110111011101110001011011001110101010;
            sine_reg0   <= 36'sb11110110101110100000011100111011001;
        end
        4801: begin
            cosine_reg0 <= 36'sb110111011101000000111110111011110101;
            sine_reg0   <= 36'sb11110110101100110101001000000100011;
        end
        4802: begin
            cosine_reg0 <= 36'sb110111011100010000100010111110000101;
            sine_reg0   <= 36'sb11110110101011001001101001101100111;
        end
        4803: begin
            cosine_reg0 <= 36'sb110111011011100000000111010101011101;
            sine_reg0   <= 36'sb11110110101001011110000001110100110;
        end
        4804: begin
            cosine_reg0 <= 36'sb110111011010101111101100000001111111;
            sine_reg0   <= 36'sb11110110100111110010010000011100000;
        end
        4805: begin
            cosine_reg0 <= 36'sb110111011001111111010001000011101100;
            sine_reg0   <= 36'sb11110110100110000110010101100010110;
        end
        4806: begin
            cosine_reg0 <= 36'sb110111011001001110110110011010100101;
            sine_reg0   <= 36'sb11110110100100011010010001001001001;
        end
        4807: begin
            cosine_reg0 <= 36'sb110111011000011110011100000110101110;
            sine_reg0   <= 36'sb11110110100010101110000011001111000;
        end
        4808: begin
            cosine_reg0 <= 36'sb110111010111101110000010001000000111;
            sine_reg0   <= 36'sb11110110100001000001101011110100101;
        end
        4809: begin
            cosine_reg0 <= 36'sb110111010110111101101000011110110100;
            sine_reg0   <= 36'sb11110110011111010101001010111010000;
        end
        4810: begin
            cosine_reg0 <= 36'sb110111010110001101001111001010110100;
            sine_reg0   <= 36'sb11110110011101101000100000011111010;
        end
        4811: begin
            cosine_reg0 <= 36'sb110111010101011100110110001100001100;
            sine_reg0   <= 36'sb11110110011011111011101100100100010;
        end
        4812: begin
            cosine_reg0 <= 36'sb110111010100101100011101100010111011;
            sine_reg0   <= 36'sb11110110011010001110101111001001010;
        end
        4813: begin
            cosine_reg0 <= 36'sb110111010011111100000101001111000101;
            sine_reg0   <= 36'sb11110110011000100001101000001110010;
        end
        4814: begin
            cosine_reg0 <= 36'sb110111010011001011101101010000101011;
            sine_reg0   <= 36'sb11110110010110110100010111110011011;
        end
        4815: begin
            cosine_reg0 <= 36'sb110111010010011011010101100111101110;
            sine_reg0   <= 36'sb11110110010101000110111101111000101;
        end
        4816: begin
            cosine_reg0 <= 36'sb110111010001101010111110010100010001;
            sine_reg0   <= 36'sb11110110010011011001011010011110000;
        end
        4817: begin
            cosine_reg0 <= 36'sb110111010000111010100111010110010110;
            sine_reg0   <= 36'sb11110110010001101011101101100011110;
        end
        4818: begin
            cosine_reg0 <= 36'sb110111010000001010010000101101111111;
            sine_reg0   <= 36'sb11110110001111111101110111001001110;
        end
        4819: begin
            cosine_reg0 <= 36'sb110111001111011001111010011011001101;
            sine_reg0   <= 36'sb11110110001110001111110111010000001;
        end
        4820: begin
            cosine_reg0 <= 36'sb110111001110101001100100011110000010;
            sine_reg0   <= 36'sb11110110001100100001101101110111001;
        end
        4821: begin
            cosine_reg0 <= 36'sb110111001101111001001110110110100000;
            sine_reg0   <= 36'sb11110110001010110011011010111110100;
        end
        4822: begin
            cosine_reg0 <= 36'sb110111001101001000111001100100101001;
            sine_reg0   <= 36'sb11110110001001000100111110100110100;
        end
        4823: begin
            cosine_reg0 <= 36'sb110111001100011000100100101000011111;
            sine_reg0   <= 36'sb11110110000111010110011000101111010;
        end
        4824: begin
            cosine_reg0 <= 36'sb110111001011101000010000000010000011;
            sine_reg0   <= 36'sb11110110000101100111101001011000110;
        end
        4825: begin
            cosine_reg0 <= 36'sb110111001010110111111011110001011000;
            sine_reg0   <= 36'sb11110110000011111000110000100011000;
        end
        4826: begin
            cosine_reg0 <= 36'sb110111001010000111100111110110100000;
            sine_reg0   <= 36'sb11110110000010001001101110001110001;
        end
        4827: begin
            cosine_reg0 <= 36'sb110111001001010111010100010001011011;
            sine_reg0   <= 36'sb11110110000000011010100010011010001;
        end
        4828: begin
            cosine_reg0 <= 36'sb110111001000100111000001000010001101;
            sine_reg0   <= 36'sb11110101111110101011001101000111010;
        end
        4829: begin
            cosine_reg0 <= 36'sb110111000111110110101110001000110111;
            sine_reg0   <= 36'sb11110101111100111011101110010101011;
        end
        4830: begin
            cosine_reg0 <= 36'sb110111000111000110011011100101011010;
            sine_reg0   <= 36'sb11110101111011001100000110000100101;
        end
        4831: begin
            cosine_reg0 <= 36'sb110111000110010110001001010111111010;
            sine_reg0   <= 36'sb11110101111001011100010100010101001;
        end
        4832: begin
            cosine_reg0 <= 36'sb110111000101100101110111100000010111;
            sine_reg0   <= 36'sb11110101110111101100011001000110111;
        end
        4833: begin
            cosine_reg0 <= 36'sb110111000100110101100101111110110011;
            sine_reg0   <= 36'sb11110101110101111100010100011010000;
        end
        4834: begin
            cosine_reg0 <= 36'sb110111000100000101010100110011010001;
            sine_reg0   <= 36'sb11110101110100001100000110001110011;
        end
        4835: begin
            cosine_reg0 <= 36'sb110111000011010101000011111101110001;
            sine_reg0   <= 36'sb11110101110010011011101110100100011;
        end
        4836: begin
            cosine_reg0 <= 36'sb110111000010100100110011011110010111;
            sine_reg0   <= 36'sb11110101110000101011001101011011111;
        end
        4837: begin
            cosine_reg0 <= 36'sb110111000001110100100011010101000100;
            sine_reg0   <= 36'sb11110101101110111010100010110101000;
        end
        4838: begin
            cosine_reg0 <= 36'sb110111000001000100010011100001111001;
            sine_reg0   <= 36'sb11110101101101001001101110101111111;
        end
        4839: begin
            cosine_reg0 <= 36'sb110111000000010100000100000100111001;
            sine_reg0   <= 36'sb11110101101011011000110001001100011;
        end
        4840: begin
            cosine_reg0 <= 36'sb110110111111100011110100111110000101;
            sine_reg0   <= 36'sb11110101101001100111101010001010110;
        end
        4841: begin
            cosine_reg0 <= 36'sb110110111110110011100110001101100000;
            sine_reg0   <= 36'sb11110101100111110110011001101011000;
        end
        4842: begin
            cosine_reg0 <= 36'sb110110111110000011010111110011001011;
            sine_reg0   <= 36'sb11110101100110000100111111101101001;
        end
        4843: begin
            cosine_reg0 <= 36'sb110110111101010011001001101111001000;
            sine_reg0   <= 36'sb11110101100100010011011100010001011;
        end
        4844: begin
            cosine_reg0 <= 36'sb110110111100100010111100000001011001;
            sine_reg0   <= 36'sb11110101100010100001101111010111101;
        end
        4845: begin
            cosine_reg0 <= 36'sb110110111011110010101110101001111111;
            sine_reg0   <= 36'sb11110101100000101111111001000000001;
        end
        4846: begin
            cosine_reg0 <= 36'sb110110111011000010100001101000111101;
            sine_reg0   <= 36'sb11110101011110111101111001001010111;
        end
        4847: begin
            cosine_reg0 <= 36'sb110110111010010010010100111110010101;
            sine_reg0   <= 36'sb11110101011101001011101111110111110;
        end
        4848: begin
            cosine_reg0 <= 36'sb110110111001100010001000101010001000;
            sine_reg0   <= 36'sb11110101011011011001011101000111001;
        end
        4849: begin
            cosine_reg0 <= 36'sb110110111000110001111100101100011000;
            sine_reg0   <= 36'sb11110101011001100111000000111000111;
        end
        4850: begin
            cosine_reg0 <= 36'sb110110111000000001110001000101000111;
            sine_reg0   <= 36'sb11110101010111110100011011001101001;
        end
        4851: begin
            cosine_reg0 <= 36'sb110110110111010001100101110100010111;
            sine_reg0   <= 36'sb11110101010110000001101100000100000;
        end
        4852: begin
            cosine_reg0 <= 36'sb110110110110100001011010111010001010;
            sine_reg0   <= 36'sb11110101010100001110110011011101100;
        end
        4853: begin
            cosine_reg0 <= 36'sb110110110101110001010000010110100001;
            sine_reg0   <= 36'sb11110101010010011011110001011001101;
        end
        4854: begin
            cosine_reg0 <= 36'sb110110110101000001000110001001011111;
            sine_reg0   <= 36'sb11110101010000101000100101111000101;
        end
        4855: begin
            cosine_reg0 <= 36'sb110110110100010000111100010011000101;
            sine_reg0   <= 36'sb11110101001110110101010000111010011;
        end
        4856: begin
            cosine_reg0 <= 36'sb110110110011100000110010110011010110;
            sine_reg0   <= 36'sb11110101001101000001110010011111001;
        end
        4857: begin
            cosine_reg0 <= 36'sb110110110010110000101001101010010010;
            sine_reg0   <= 36'sb11110101001011001110001010100110110;
        end
        4858: begin
            cosine_reg0 <= 36'sb110110110010000000100000110111111100;
            sine_reg0   <= 36'sb11110101001001011010011001010001100;
        end
        4859: begin
            cosine_reg0 <= 36'sb110110110001010000011000011100010110;
            sine_reg0   <= 36'sb11110101000111100110011110011111011;
        end
        4860: begin
            cosine_reg0 <= 36'sb110110110000100000010000010111100010;
            sine_reg0   <= 36'sb11110101000101110010011010010000100;
        end
        4861: begin
            cosine_reg0 <= 36'sb110110101111110000001000101001100001;
            sine_reg0   <= 36'sb11110101000011111110001100100100110;
        end
        4862: begin
            cosine_reg0 <= 36'sb110110101111000000000001010010010101;
            sine_reg0   <= 36'sb11110101000010001001110101011100100;
        end
        4863: begin
            cosine_reg0 <= 36'sb110110101110001111111010010010000001;
            sine_reg0   <= 36'sb11110101000000010101010100110111100;
        end
        4864: begin
            cosine_reg0 <= 36'sb110110101101011111110011101000100110;
            sine_reg0   <= 36'sb11110100111110100000101010110110001;
        end
        4865: begin
            cosine_reg0 <= 36'sb110110101100101111101101010110000101;
            sine_reg0   <= 36'sb11110100111100101011110111011000001;
        end
        4866: begin
            cosine_reg0 <= 36'sb110110101011111111100111011010100001;
            sine_reg0   <= 36'sb11110100111010110110111010011101111;
        end
        4867: begin
            cosine_reg0 <= 36'sb110110101011001111100001110101111100;
            sine_reg0   <= 36'sb11110100111001000001110100000111010;
        end
        4868: begin
            cosine_reg0 <= 36'sb110110101010011111011100101000010111;
            sine_reg0   <= 36'sb11110100110111001100100100010100011;
        end
        4869: begin
            cosine_reg0 <= 36'sb110110101001101111010111110001110101;
            sine_reg0   <= 36'sb11110100110101010111001011000101011;
        end
        4870: begin
            cosine_reg0 <= 36'sb110110101000111111010011010010010110;
            sine_reg0   <= 36'sb11110100110011100001101000011010010;
        end
        4871: begin
            cosine_reg0 <= 36'sb110110101000001111001111001001111110;
            sine_reg0   <= 36'sb11110100110001101011111100010011000;
        end
        4872: begin
            cosine_reg0 <= 36'sb110110100111011111001011011000101110;
            sine_reg0   <= 36'sb11110100101111110110000110101111111;
        end
        4873: begin
            cosine_reg0 <= 36'sb110110100110101111000111111110100111;
            sine_reg0   <= 36'sb11110100101110000000000111110000111;
        end
        4874: begin
            cosine_reg0 <= 36'sb110110100101111111000100111011101100;
            sine_reg0   <= 36'sb11110100101100001001111111010110001;
        end
        4875: begin
            cosine_reg0 <= 36'sb110110100101001111000010001111111110;
            sine_reg0   <= 36'sb11110100101010010011101101011111100;
        end
        4876: begin
            cosine_reg0 <= 36'sb110110100100011110111111111011011111;
            sine_reg0   <= 36'sb11110100101000011101010010001101010;
        end
        4877: begin
            cosine_reg0 <= 36'sb110110100011101110111101111110010010;
            sine_reg0   <= 36'sb11110100100110100110101101011111011;
        end
        4878: begin
            cosine_reg0 <= 36'sb110110100010111110111100011000010111;
            sine_reg0   <= 36'sb11110100100100101111111111010110000;
        end
        4879: begin
            cosine_reg0 <= 36'sb110110100010001110111011001001110010;
            sine_reg0   <= 36'sb11110100100010111001000111110001001;
        end
        4880: begin
            cosine_reg0 <= 36'sb110110100001011110111010010010100011;
            sine_reg0   <= 36'sb11110100100001000010000110110000111;
        end
        4881: begin
            cosine_reg0 <= 36'sb110110100000101110111001110010101100;
            sine_reg0   <= 36'sb11110100011111001010111100010101010;
        end
        4882: begin
            cosine_reg0 <= 36'sb110110011111111110111001101010010000;
            sine_reg0   <= 36'sb11110100011101010011101000011110011;
        end
        4883: begin
            cosine_reg0 <= 36'sb110110011111001110111001111001010000;
            sine_reg0   <= 36'sb11110100011011011100001011001100011;
        end
        4884: begin
            cosine_reg0 <= 36'sb110110011110011110111010011111101111;
            sine_reg0   <= 36'sb11110100011001100100100100011111010;
        end
        4885: begin
            cosine_reg0 <= 36'sb110110011101101110111011011101101101;
            sine_reg0   <= 36'sb11110100010111101100110100010111001;
        end
        4886: begin
            cosine_reg0 <= 36'sb110110011100111110111100110011001101;
            sine_reg0   <= 36'sb11110100010101110100111010110100001;
        end
        4887: begin
            cosine_reg0 <= 36'sb110110011100001110111110100000010000;
            sine_reg0   <= 36'sb11110100010011111100110111110110001;
        end
        4888: begin
            cosine_reg0 <= 36'sb110110011011011111000000100100111001;
            sine_reg0   <= 36'sb11110100010010000100101011011101010;
        end
        4889: begin
            cosine_reg0 <= 36'sb110110011010101111000011000001001010;
            sine_reg0   <= 36'sb11110100010000001100010101101001110;
        end
        4890: begin
            cosine_reg0 <= 36'sb110110011001111111000101110101000011;
            sine_reg0   <= 36'sb11110100001110010011110110011011100;
        end
        4891: begin
            cosine_reg0 <= 36'sb110110011001001111001001000000101000;
            sine_reg0   <= 36'sb11110100001100011011001101110010110;
        end
        4892: begin
            cosine_reg0 <= 36'sb110110011000011111001100100011111001;
            sine_reg0   <= 36'sb11110100001010100010011011101111011;
        end
        4893: begin
            cosine_reg0 <= 36'sb110110010111101111010000011110111001;
            sine_reg0   <= 36'sb11110100001000101001100000010001101;
        end
        4894: begin
            cosine_reg0 <= 36'sb110110010110111111010100110001101010;
            sine_reg0   <= 36'sb11110100000110110000011011011001100;
        end
        4895: begin
            cosine_reg0 <= 36'sb110110010110001111011001011100001101;
            sine_reg0   <= 36'sb11110100000100110111001101000111000;
        end
        4896: begin
            cosine_reg0 <= 36'sb110110010101011111011110011110100100;
            sine_reg0   <= 36'sb11110100000010111101110101011010010;
        end
        4897: begin
            cosine_reg0 <= 36'sb110110010100101111100011111000110010;
            sine_reg0   <= 36'sb11110100000001000100010100010011011;
        end
        4898: begin
            cosine_reg0 <= 36'sb110110010011111111101001101010110111;
            sine_reg0   <= 36'sb11110011111111001010101001110010100;
        end
        4899: begin
            cosine_reg0 <= 36'sb110110010011001111101111110100110110;
            sine_reg0   <= 36'sb11110011111101010000110101110111100;
        end
        4900: begin
            cosine_reg0 <= 36'sb110110010010011111110110010110110001;
            sine_reg0   <= 36'sb11110011111011010110111000100010101;
        end
        4901: begin
            cosine_reg0 <= 36'sb110110010001101111111101010000101001;
            sine_reg0   <= 36'sb11110011111001011100110001110011111;
        end
        4902: begin
            cosine_reg0 <= 36'sb110110010001000000000100100010100001;
            sine_reg0   <= 36'sb11110011110111100010100001101011010;
        end
        4903: begin
            cosine_reg0 <= 36'sb110110010000010000001100001100011010;
            sine_reg0   <= 36'sb11110011110101101000001000001001000;
        end
        4904: begin
            cosine_reg0 <= 36'sb110110001111100000010100001110010110;
            sine_reg0   <= 36'sb11110011110011101101100101001101000;
        end
        4905: begin
            cosine_reg0 <= 36'sb110110001110110000011100101000010111;
            sine_reg0   <= 36'sb11110011110001110010111000110111100;
        end
        4906: begin
            cosine_reg0 <= 36'sb110110001110000000100101011010011110;
            sine_reg0   <= 36'sb11110011101111111000000011001000100;
        end
        4907: begin
            cosine_reg0 <= 36'sb110110001101010000101110100100101110;
            sine_reg0   <= 36'sb11110011101101111101000100000000001;
        end
        4908: begin
            cosine_reg0 <= 36'sb110110001100100000111000000111001001;
            sine_reg0   <= 36'sb11110011101100000001111011011110011;
        end
        4909: begin
            cosine_reg0 <= 36'sb110110001011110001000010000001110000;
            sine_reg0   <= 36'sb11110011101010000110101001100011010;
        end
        4910: begin
            cosine_reg0 <= 36'sb110110001011000001001100010100100100;
            sine_reg0   <= 36'sb11110011101000001011001110001111000;
        end
        4911: begin
            cosine_reg0 <= 36'sb110110001010010001010110111111101001;
            sine_reg0   <= 36'sb11110011100110001111101001100001101;
        end
        4912: begin
            cosine_reg0 <= 36'sb110110001001100001100010000011000000;
            sine_reg0   <= 36'sb11110011100100010011111011011011010;
        end
        4913: begin
            cosine_reg0 <= 36'sb110110001000110001101101011110101010;
            sine_reg0   <= 36'sb11110011100010011000000011111011110;
        end
        4914: begin
            cosine_reg0 <= 36'sb110110001000000001111001010010101010;
            sine_reg0   <= 36'sb11110011100000011100000011000011100;
        end
        4915: begin
            cosine_reg0 <= 36'sb110110000111010010000101011111000001;
            sine_reg0   <= 36'sb11110011011110011111111000110010011;
        end
        4916: begin
            cosine_reg0 <= 36'sb110110000110100010010010000011110001;
            sine_reg0   <= 36'sb11110011011100100011100101001000100;
        end
        4917: begin
            cosine_reg0 <= 36'sb110110000101110010011111000000111100;
            sine_reg0   <= 36'sb11110011011010100111001000000101111;
        end
        4918: begin
            cosine_reg0 <= 36'sb110110000101000010101100010110100100;
            sine_reg0   <= 36'sb11110011011000101010100001101010101;
        end
        4919: begin
            cosine_reg0 <= 36'sb110110000100010010111010000100101011;
            sine_reg0   <= 36'sb11110011010110101101110001110111000;
        end
        4920: begin
            cosine_reg0 <= 36'sb110110000011100011001000001011010010;
            sine_reg0   <= 36'sb11110011010100110000111000101010110;
        end
        4921: begin
            cosine_reg0 <= 36'sb110110000010110011010110101010011100;
            sine_reg0   <= 36'sb11110011010010110011110110000110010;
        end
        4922: begin
            cosine_reg0 <= 36'sb110110000010000011100101100010001010;
            sine_reg0   <= 36'sb11110011010000110110101010001001011;
        end
        4923: begin
            cosine_reg0 <= 36'sb110110000001010011110100110010011110;
            sine_reg0   <= 36'sb11110011001110111001010100110100011;
        end
        4924: begin
            cosine_reg0 <= 36'sb110110000000100100000100011011011010;
            sine_reg0   <= 36'sb11110011001100111011110110000111001;
        end
        4925: begin
            cosine_reg0 <= 36'sb110101111111110100010100011101000000;
            sine_reg0   <= 36'sb11110011001010111110001110000001110;
        end
        4926: begin
            cosine_reg0 <= 36'sb110101111111000100100100110111010001;
            sine_reg0   <= 36'sb11110011001001000000011100100100100;
        end
        4927: begin
            cosine_reg0 <= 36'sb110101111110010100110101101010001111;
            sine_reg0   <= 36'sb11110011000111000010100001101111010;
        end
        4928: begin
            cosine_reg0 <= 36'sb110101111101100101000110110101111101;
            sine_reg0   <= 36'sb11110011000101000100011101100010001;
        end
        4929: begin
            cosine_reg0 <= 36'sb110101111100110101011000011010011100;
            sine_reg0   <= 36'sb11110011000011000110001111111101010;
        end
        4930: begin
            cosine_reg0 <= 36'sb110101111100000101101010010111101110;
            sine_reg0   <= 36'sb11110011000001000111111001000000110;
        end
        4931: begin
            cosine_reg0 <= 36'sb110101111011010101111100101101110101;
            sine_reg0   <= 36'sb11110010111111001001011000101100101;
        end
        4932: begin
            cosine_reg0 <= 36'sb110101111010100110001111011100110011;
            sine_reg0   <= 36'sb11110010111101001010101111000000111;
        end
        4933: begin
            cosine_reg0 <= 36'sb110101111001110110100010100100101000;
            sine_reg0   <= 36'sb11110010111011001011111011111101101;
        end
        4934: begin
            cosine_reg0 <= 36'sb110101111001000110110110000101011001;
            sine_reg0   <= 36'sb11110010111001001100111111100011001;
        end
        4935: begin
            cosine_reg0 <= 36'sb110101111000010111001001111111000101;
            sine_reg0   <= 36'sb11110010110111001101111001110001001;
        end
        4936: begin
            cosine_reg0 <= 36'sb110101110111100111011110010001101111;
            sine_reg0   <= 36'sb11110010110101001110101010101000000;
        end
        4937: begin
            cosine_reg0 <= 36'sb110101110110110111110010111101011001;
            sine_reg0   <= 36'sb11110010110011001111010010000111110;
        end
        4938: begin
            cosine_reg0 <= 36'sb110101110110001000001000000010000101;
            sine_reg0   <= 36'sb11110010110001001111110000010000011;
        end
        4939: begin
            cosine_reg0 <= 36'sb110101110101011000011101011111110100;
            sine_reg0   <= 36'sb11110010101111010000000101000001111;
        end
        4940: begin
            cosine_reg0 <= 36'sb110101110100101000110011010110101001;
            sine_reg0   <= 36'sb11110010101101010000010000011100101;
        end
        4941: begin
            cosine_reg0 <= 36'sb110101110011111001001001100110100101;
            sine_reg0   <= 36'sb11110010101011010000010010100000011;
        end
        4942: begin
            cosine_reg0 <= 36'sb110101110011001001100000001111101001;
            sine_reg0   <= 36'sb11110010101001010000001011001101011;
        end
        4943: begin
            cosine_reg0 <= 36'sb110101110010011001110111010001111001;
            sine_reg0   <= 36'sb11110010100111001111111010100011110;
        end
        4944: begin
            cosine_reg0 <= 36'sb110101110001101010001110101101010101;
            sine_reg0   <= 36'sb11110010100101001111100000100011100;
        end
        4945: begin
            cosine_reg0 <= 36'sb110101110000111010100110100010000000;
            sine_reg0   <= 36'sb11110010100011001110111101001100101;
        end
        4946: begin
            cosine_reg0 <= 36'sb110101110000001010111110101111111011;
            sine_reg0   <= 36'sb11110010100001001110010000011111010;
        end
        4947: begin
            cosine_reg0 <= 36'sb110101101111011011010111010111001001;
            sine_reg0   <= 36'sb11110010011111001101011010011011101;
        end
        4948: begin
            cosine_reg0 <= 36'sb110101101110101011110000010111101010;
            sine_reg0   <= 36'sb11110010011101001100011011000001101;
        end
        4949: begin
            cosine_reg0 <= 36'sb110101101101111100001001110001100010;
            sine_reg0   <= 36'sb11110010011011001011010010010001011;
        end
        4950: begin
            cosine_reg0 <= 36'sb110101101101001100100011100100110001;
            sine_reg0   <= 36'sb11110010011001001010000000001010111;
        end
        4951: begin
            cosine_reg0 <= 36'sb110101101100011100111101110001011001;
            sine_reg0   <= 36'sb11110010010111001000100100101110011;
        end
        4952: begin
            cosine_reg0 <= 36'sb110101101011101101011000010111011101;
            sine_reg0   <= 36'sb11110010010101000110111111111100000;
        end
        4953: begin
            cosine_reg0 <= 36'sb110101101010111101110011010110111110;
            sine_reg0   <= 36'sb11110010010011000101010001110011100;
        end
        4954: begin
            cosine_reg0 <= 36'sb110101101010001110001110101111111110;
            sine_reg0   <= 36'sb11110010010001000011011010010101010;
        end
        4955: begin
            cosine_reg0 <= 36'sb110101101001011110101010100010011111;
            sine_reg0   <= 36'sb11110010001111000001011001100001010;
        end
        4956: begin
            cosine_reg0 <= 36'sb110101101000101111000110101110100011;
            sine_reg0   <= 36'sb11110010001100111111001111010111100;
        end
        4957: begin
            cosine_reg0 <= 36'sb110101100111111111100011010100001011;
            sine_reg0   <= 36'sb11110010001010111100111011111000001;
        end
        4958: begin
            cosine_reg0 <= 36'sb110101100111010000000000010011011010;
            sine_reg0   <= 36'sb11110010001000111010011111000011010;
        end
        4959: begin
            cosine_reg0 <= 36'sb110101100110100000011101101100010000;
            sine_reg0   <= 36'sb11110010000110110111111000111001000;
        end
        4960: begin
            cosine_reg0 <= 36'sb110101100101110000111011011110110001;
            sine_reg0   <= 36'sb11110010000100110101001001011001010;
        end
        4961: begin
            cosine_reg0 <= 36'sb110101100101000001011001101010111110;
            sine_reg0   <= 36'sb11110010000010110010010000100100010;
        end
        4962: begin
            cosine_reg0 <= 36'sb110101100100010001111000010000111000;
            sine_reg0   <= 36'sb11110010000000101111001110011010000;
        end
        4963: begin
            cosine_reg0 <= 36'sb110101100011100010010111010000100010;
            sine_reg0   <= 36'sb11110001111110101100000010111010101;
        end
        4964: begin
            cosine_reg0 <= 36'sb110101100010110010110110101001111110;
            sine_reg0   <= 36'sb11110001111100101000101110000110010;
        end
        4965: begin
            cosine_reg0 <= 36'sb110101100010000011010110011101001100;
            sine_reg0   <= 36'sb11110001111010100101001111111100111;
        end
        4966: begin
            cosine_reg0 <= 36'sb110101100001010011110110101010010000;
            sine_reg0   <= 36'sb11110001111000100001101000011110100;
        end
        4967: begin
            cosine_reg0 <= 36'sb110101100000100100010111010001001010;
            sine_reg0   <= 36'sb11110001110110011101110111101011011;
        end
        4968: begin
            cosine_reg0 <= 36'sb110101011111110100111000010001111101;
            sine_reg0   <= 36'sb11110001110100011001111101100011101;
        end
        4969: begin
            cosine_reg0 <= 36'sb110101011111000101011001101100101011;
            sine_reg0   <= 36'sb11110001110010010101111010000111000;
        end
        4970: begin
            cosine_reg0 <= 36'sb110101011110010101111011100001010101;
            sine_reg0   <= 36'sb11110001110000010001101101010101111;
        end
        4971: begin
            cosine_reg0 <= 36'sb110101011101100110011101101111111101;
            sine_reg0   <= 36'sb11110001101110001101010111010000010;
        end
        4972: begin
            cosine_reg0 <= 36'sb110101011100110111000000011000100101;
            sine_reg0   <= 36'sb11110001101100001000110111110110010;
        end
        4973: begin
            cosine_reg0 <= 36'sb110101011100000111100011011011001111;
            sine_reg0   <= 36'sb11110001101010000100001111000111111;
        end
        4974: begin
            cosine_reg0 <= 36'sb110101011011011000000110110111111101;
            sine_reg0   <= 36'sb11110001100111111111011101000101010;
        end
        4975: begin
            cosine_reg0 <= 36'sb110101011010101000101010101110110000;
            sine_reg0   <= 36'sb11110001100101111010100001101110011;
        end
        4976: begin
            cosine_reg0 <= 36'sb110101011001111001001110111111101010;
            sine_reg0   <= 36'sb11110001100011110101011101000011011;
        end
        4977: begin
            cosine_reg0 <= 36'sb110101011001001001110011101010101110;
            sine_reg0   <= 36'sb11110001100001110000001111000100011;
        end
        4978: begin
            cosine_reg0 <= 36'sb110101011000011010011000101111111101;
            sine_reg0   <= 36'sb11110001011111101010110111110001100;
        end
        4979: begin
            cosine_reg0 <= 36'sb110101010111101010111110001111011000;
            sine_reg0   <= 36'sb11110001011101100101010111001010110;
        end
        4980: begin
            cosine_reg0 <= 36'sb110101010110111011100100001001000010;
            sine_reg0   <= 36'sb11110001011011011111101101010000001;
        end
        4981: begin
            cosine_reg0 <= 36'sb110101010110001100001010011100111101;
            sine_reg0   <= 36'sb11110001011001011001111010000001111;
        end
        4982: begin
            cosine_reg0 <= 36'sb110101010101011100110001001011001010;
            sine_reg0   <= 36'sb11110001010111010011111101100000000;
        end
        4983: begin
            cosine_reg0 <= 36'sb110101010100101101011000010011101011;
            sine_reg0   <= 36'sb11110001010101001101110111101010101;
        end
        4984: begin
            cosine_reg0 <= 36'sb110101010011111101111111110110100010;
            sine_reg0   <= 36'sb11110001010011000111101000100001101;
        end
        4985: begin
            cosine_reg0 <= 36'sb110101010011001110100111110011110001;
            sine_reg0   <= 36'sb11110001010001000001010000000101011;
        end
        4986: begin
            cosine_reg0 <= 36'sb110101010010011111010000001011011001;
            sine_reg0   <= 36'sb11110001001110111010101110010101110;
        end
        4987: begin
            cosine_reg0 <= 36'sb110101010001101111111000111101011101;
            sine_reg0   <= 36'sb11110001001100110100000011010011000;
        end
        4988: begin
            cosine_reg0 <= 36'sb110101010001000000100010001001111110;
            sine_reg0   <= 36'sb11110001001010101101001110111101001;
        end
        4989: begin
            cosine_reg0 <= 36'sb110101010000010001001011110000111110;
            sine_reg0   <= 36'sb11110001001000100110010001010100001;
        end
        4990: begin
            cosine_reg0 <= 36'sb110101001111100001110101110010011111;
            sine_reg0   <= 36'sb11110001000110011111001010011000001;
        end
        4991: begin
            cosine_reg0 <= 36'sb110101001110110010100000001110100011;
            sine_reg0   <= 36'sb11110001000100010111111010001001010;
        end
        4992: begin
            cosine_reg0 <= 36'sb110101001110000011001011000101001011;
            sine_reg0   <= 36'sb11110001000010010000100000100111101;
        end
        4993: begin
            cosine_reg0 <= 36'sb110101001101010011110110010110011010;
            sine_reg0   <= 36'sb11110001000000001000111101110011001;
        end
        4994: begin
            cosine_reg0 <= 36'sb110101001100100100100010000010010001;
            sine_reg0   <= 36'sb11110000111110000001010001101100001;
        end
        4995: begin
            cosine_reg0 <= 36'sb110101001011110101001110001000110010;
            sine_reg0   <= 36'sb11110000111011111001011100010010100;
        end
        4996: begin
            cosine_reg0 <= 36'sb110101001011000101111010101001111110;
            sine_reg0   <= 36'sb11110000111001110001011101100110011;
        end
        4997: begin
            cosine_reg0 <= 36'sb110101001010010110100111100101111001;
            sine_reg0   <= 36'sb11110000110111101001010101100111111;
        end
        4998: begin
            cosine_reg0 <= 36'sb110101001001100111010100111100100011;
            sine_reg0   <= 36'sb11110000110101100001000100010111001;
        end
        4999: begin
            cosine_reg0 <= 36'sb110101001000111000000010101101111110;
            sine_reg0   <= 36'sb11110000110011011000101001110100000;
        end
        5000: begin
            cosine_reg0 <= 36'sb110101001000001000110000111010001101;
            sine_reg0   <= 36'sb11110000110001010000000101111110110;
        end
        5001: begin
            cosine_reg0 <= 36'sb110101000111011001011111100001010000;
            sine_reg0   <= 36'sb11110000101111000111011000110111100;
        end
        5002: begin
            cosine_reg0 <= 36'sb110101000110101010001110100011001010;
            sine_reg0   <= 36'sb11110000101100111110100010011110001;
        end
        5003: begin
            cosine_reg0 <= 36'sb110101000101111010111101111111111101;
            sine_reg0   <= 36'sb11110000101010110101100010110011000;
        end
        5004: begin
            cosine_reg0 <= 36'sb110101000101001011101101110111101010;
            sine_reg0   <= 36'sb11110000101000101100011001110101111;
        end
        5005: begin
            cosine_reg0 <= 36'sb110101000100011100011110001010010100;
            sine_reg0   <= 36'sb11110000100110100011000111100111001;
        end
        5006: begin
            cosine_reg0 <= 36'sb110101000011101101001110110111111100;
            sine_reg0   <= 36'sb11110000100100011001101100000110110;
        end
        5007: begin
            cosine_reg0 <= 36'sb110101000010111110000000000000100011;
            sine_reg0   <= 36'sb11110000100010010000000111010100110;
        end
        5008: begin
            cosine_reg0 <= 36'sb110101000010001110110001100100001101;
            sine_reg0   <= 36'sb11110000100000000110011001010001001;
        end
        5009: begin
            cosine_reg0 <= 36'sb110101000001011111100011100010111001;
            sine_reg0   <= 36'sb11110000011101111100100001111100010;
        end
        5010: begin
            cosine_reg0 <= 36'sb110101000000110000010101111100101100;
            sine_reg0   <= 36'sb11110000011011110010100001010110000;
        end
        5011: begin
            cosine_reg0 <= 36'sb110101000000000001001000110001100101;
            sine_reg0   <= 36'sb11110000011001101000010111011110100;
        end
        5012: begin
            cosine_reg0 <= 36'sb110100111111010001111100000001100111;
            sine_reg0   <= 36'sb11110000010111011110000100010101110;
        end
        5013: begin
            cosine_reg0 <= 36'sb110100111110100010101111101100110100;
            sine_reg0   <= 36'sb11110000010101010011100111111100000;
        end
        5014: begin
            cosine_reg0 <= 36'sb110100111101110011100011110011001110;
            sine_reg0   <= 36'sb11110000010011001001000010010001010;
        end
        5015: begin
            cosine_reg0 <= 36'sb110100111101000100011000010100110111;
            sine_reg0   <= 36'sb11110000010000111110010011010101101;
        end
        5016: begin
            cosine_reg0 <= 36'sb110100111100010101001101010001101111;
            sine_reg0   <= 36'sb11110000001110110011011011001001001;
        end
        5017: begin
            cosine_reg0 <= 36'sb110100111011100110000010101001111010;
            sine_reg0   <= 36'sb11110000001100101000011001101011111;
        end
        5018: begin
            cosine_reg0 <= 36'sb110100111010110110111000011101011001;
            sine_reg0   <= 36'sb11110000001010011101001110111110000;
        end
        5019: begin
            cosine_reg0 <= 36'sb110100111010000111101110101100001101;
            sine_reg0   <= 36'sb11110000001000010001111010111111100;
        end
        5020: begin
            cosine_reg0 <= 36'sb110100111001011000100101010110011001;
            sine_reg0   <= 36'sb11110000000110000110011101110000100;
        end
        5021: begin
            cosine_reg0 <= 36'sb110100111000101001011100011011111110;
            sine_reg0   <= 36'sb11110000000011111010110111010001001;
        end
        5022: begin
            cosine_reg0 <= 36'sb110100110111111010010011111100111111;
            sine_reg0   <= 36'sb11110000000001101111000111100001011;
        end
        5023: begin
            cosine_reg0 <= 36'sb110100110111001011001011111001011100;
            sine_reg0   <= 36'sb11101111111111100011001110100001011;
        end
        5024: begin
            cosine_reg0 <= 36'sb110100110110011100000100010001011000;
            sine_reg0   <= 36'sb11101111111101010111001100010001010;
        end
        5025: begin
            cosine_reg0 <= 36'sb110100110101101100111101000100110101;
            sine_reg0   <= 36'sb11101111111011001011000000110001001;
        end
        5026: begin
            cosine_reg0 <= 36'sb110100110100111101110110010011110101;
            sine_reg0   <= 36'sb11101111111000111110101100000000111;
        end
        5027: begin
            cosine_reg0 <= 36'sb110100110100001110101111111110011001;
            sine_reg0   <= 36'sb11101111110110110010001110000000111;
        end
        5028: begin
            cosine_reg0 <= 36'sb110100110011011111101010000100100010;
            sine_reg0   <= 36'sb11101111110100100101100110110000111;
        end
        5029: begin
            cosine_reg0 <= 36'sb110100110010110000100100100110010100;
            sine_reg0   <= 36'sb11101111110010011000110110010001010;
        end
        5030: begin
            cosine_reg0 <= 36'sb110100110010000001011111100011101111;
            sine_reg0   <= 36'sb11101111110000001011111100100010000;
        end
        5031: begin
            cosine_reg0 <= 36'sb110100110001010010011010111100110110;
            sine_reg0   <= 36'sb11101111101101111110111001100011001;
        end
        5032: begin
            cosine_reg0 <= 36'sb110100110000100011010110110001101011;
            sine_reg0   <= 36'sb11101111101011110001101101010100110;
        end
        5033: begin
            cosine_reg0 <= 36'sb110100101111110100010011000010001110;
            sine_reg0   <= 36'sb11101111101001100100010111110111000;
        end
        5034: begin
            cosine_reg0 <= 36'sb110100101111000101001111101110100011;
            sine_reg0   <= 36'sb11101111100111010110111001001010000;
        end
        5035: begin
            cosine_reg0 <= 36'sb110100101110010110001100110110101010;
            sine_reg0   <= 36'sb11101111100101001001010001001101101;
        end
        5036: begin
            cosine_reg0 <= 36'sb110100101101100111001010011010100110;
            sine_reg0   <= 36'sb11101111100010111011100000000010010;
        end
        5037: begin
            cosine_reg0 <= 36'sb110100101100111000001000011010011000;
            sine_reg0   <= 36'sb11101111100000101101100101100111110;
        end
        5038: begin
            cosine_reg0 <= 36'sb110100101100001001000110110110000010;
            sine_reg0   <= 36'sb11101111011110011111100001111110010;
        end
        5039: begin
            cosine_reg0 <= 36'sb110100101011011010000101101101100111;
            sine_reg0   <= 36'sb11101111011100010001010101000110000;
        end
        5040: begin
            cosine_reg0 <= 36'sb110100101010101011000101000001000111;
            sine_reg0   <= 36'sb11101111011010000010111110111110111;
        end
        5041: begin
            cosine_reg0 <= 36'sb110100101001111100000100110000100110;
            sine_reg0   <= 36'sb11101111010111110100011111101001000;
        end
        5042: begin
            cosine_reg0 <= 36'sb110100101001001101000100111100000011;
            sine_reg0   <= 36'sb11101111010101100101110111000100100;
        end
        5043: begin
            cosine_reg0 <= 36'sb110100101000011110000101100011100010;
            sine_reg0   <= 36'sb11101111010011010111000101010001100;
        end
        5044: begin
            cosine_reg0 <= 36'sb110100100111101111000110100111000100;
            sine_reg0   <= 36'sb11101111010001001000001010010000000;
        end
        5045: begin
            cosine_reg0 <= 36'sb110100100111000000001000000110101011;
            sine_reg0   <= 36'sb11101111001110111001000110000000001;
        end
        5046: begin
            cosine_reg0 <= 36'sb110100100110010001001010000010011000;
            sine_reg0   <= 36'sb11101111001100101001111000100010000;
        end
        5047: begin
            cosine_reg0 <= 36'sb110100100101100010001100011010001111;
            sine_reg0   <= 36'sb11101111001010011010100001110101110;
        end
        5048: begin
            cosine_reg0 <= 36'sb110100100100110011001111001110001111;
            sine_reg0   <= 36'sb11101111001000001011000001111011010;
        end
        5049: begin
            cosine_reg0 <= 36'sb110100100100000100010010011110011100;
            sine_reg0   <= 36'sb11101111000101111011011000110010111;
        end
        5050: begin
            cosine_reg0 <= 36'sb110100100011010101010110001010110110;
            sine_reg0   <= 36'sb11101111000011101011100110011100100;
        end
        5051: begin
            cosine_reg0 <= 36'sb110100100010100110011010010011100001;
            sine_reg0   <= 36'sb11101111000001011011101010111000010;
        end
        5052: begin
            cosine_reg0 <= 36'sb110100100001110111011110111000011101;
            sine_reg0   <= 36'sb11101110111111001011100110000110010;
        end
        5053: begin
            cosine_reg0 <= 36'sb110100100001001000100011111001101100;
            sine_reg0   <= 36'sb11101110111100111011011000000110100;
        end
        5054: begin
            cosine_reg0 <= 36'sb110100100000011001101001010111010001;
            sine_reg0   <= 36'sb11101110111010101011000000111001010;
        end
        5055: begin
            cosine_reg0 <= 36'sb110100011111101010101111010001001101;
            sine_reg0   <= 36'sb11101110111000011010100000011110100;
        end
        5056: begin
            cosine_reg0 <= 36'sb110100011110111011110101100111100001;
            sine_reg0   <= 36'sb11101110110110001001110110110110010;
        end
        5057: begin
            cosine_reg0 <= 36'sb110100011110001100111100011010010000;
            sine_reg0   <= 36'sb11101110110011111001000100000000110;
        end
        5058: begin
            cosine_reg0 <= 36'sb110100011101011110000011101001011100;
            sine_reg0   <= 36'sb11101110110001101000000111111110000;
        end
        5059: begin
            cosine_reg0 <= 36'sb110100011100101111001011010101000110;
            sine_reg0   <= 36'sb11101110101111010111000010101110001;
        end
        5060: begin
            cosine_reg0 <= 36'sb110100011100000000010011011101001111;
            sine_reg0   <= 36'sb11101110101101000101110100010001001;
        end
        5061: begin
            cosine_reg0 <= 36'sb110100011011010001011100000001111011;
            sine_reg0   <= 36'sb11101110101010110100011100100111001;
        end
        5062: begin
            cosine_reg0 <= 36'sb110100011010100010100101000011001011;
            sine_reg0   <= 36'sb11101110101000100010111011110000010;
        end
        5063: begin
            cosine_reg0 <= 36'sb110100011001110011101110100000111111;
            sine_reg0   <= 36'sb11101110100110010001010001101100101;
        end
        5064: begin
            cosine_reg0 <= 36'sb110100011001000100111000011011011100;
            sine_reg0   <= 36'sb11101110100011111111011110011100010;
        end
        5065: begin
            cosine_reg0 <= 36'sb110100011000010110000010110010100001;
            sine_reg0   <= 36'sb11101110100001101101100001111111010;
        end
        5066: begin
            cosine_reg0 <= 36'sb110100010111100111001101100110010001;
            sine_reg0   <= 36'sb11101110011111011011011100010101101;
        end
        5067: begin
            cosine_reg0 <= 36'sb110100010110111000011000110110101110;
            sine_reg0   <= 36'sb11101110011101001001001101011111101;
        end
        5068: begin
            cosine_reg0 <= 36'sb110100010110001001100100100011111001;
            sine_reg0   <= 36'sb11101110011010110110110101011101010;
        end
        5069: begin
            cosine_reg0 <= 36'sb110100010101011010110000101101110101;
            sine_reg0   <= 36'sb11101110011000100100010100001110101;
        end
        5070: begin
            cosine_reg0 <= 36'sb110100010100101011111101010100100011;
            sine_reg0   <= 36'sb11101110010110010001101001110011110;
        end
        5071: begin
            cosine_reg0 <= 36'sb110100010011111101001010011000000100;
            sine_reg0   <= 36'sb11101110010011111110110110001100111;
        end
        5072: begin
            cosine_reg0 <= 36'sb110100010011001110010111111000011100;
            sine_reg0   <= 36'sb11101110010001101011111001011001111;
        end
        5073: begin
            cosine_reg0 <= 36'sb110100010010011111100101110101101011;
            sine_reg0   <= 36'sb11101110001111011000110011011011000;
        end
        5074: begin
            cosine_reg0 <= 36'sb110100010001110000110100001111110011;
            sine_reg0   <= 36'sb11101110001101000101100100010000011;
        end
        5075: begin
            cosine_reg0 <= 36'sb110100010001000010000011000110110111;
            sine_reg0   <= 36'sb11101110001010110010001011111001111;
        end
        5076: begin
            cosine_reg0 <= 36'sb110100010000010011010010011010110111;
            sine_reg0   <= 36'sb11101110001000011110101010010111110;
        end
        5077: begin
            cosine_reg0 <= 36'sb110100001111100100100010001011110110;
            sine_reg0   <= 36'sb11101110000110001010111111101010001;
        end
        5078: begin
            cosine_reg0 <= 36'sb110100001110110101110010011001110110;
            sine_reg0   <= 36'sb11101110000011110111001011110001000;
        end
        5079: begin
            cosine_reg0 <= 36'sb110100001110000111000011000100111000;
            sine_reg0   <= 36'sb11101110000001100011001110101100011;
        end
        5080: begin
            cosine_reg0 <= 36'sb110100001101011000010100001100111110;
            sine_reg0   <= 36'sb11101101111111001111001000011100100;
        end
        5081: begin
            cosine_reg0 <= 36'sb110100001100101001100101110010001010;
            sine_reg0   <= 36'sb11101101111100111010111001000001100;
        end
        5082: begin
            cosine_reg0 <= 36'sb110100001011111010110111110100011110;
            sine_reg0   <= 36'sb11101101111010100110100000011011011;
        end
        5083: begin
            cosine_reg0 <= 36'sb110100001011001100001010010011111011;
            sine_reg0   <= 36'sb11101101111000010001111110101010001;
        end
        5084: begin
            cosine_reg0 <= 36'sb110100001010011101011101010000100100;
            sine_reg0   <= 36'sb11101101110101111101010011101110000;
        end
        5085: begin
            cosine_reg0 <= 36'sb110100001001101110110000101010011010;
            sine_reg0   <= 36'sb11101101110011101000011111100110111;
        end
        5086: begin
            cosine_reg0 <= 36'sb110100001001000000000100100001011111;
            sine_reg0   <= 36'sb11101101110001010011100010010101001;
        end
        5087: begin
            cosine_reg0 <= 36'sb110100001000010001011000110101110100;
            sine_reg0   <= 36'sb11101101101110111110011011111000110;
        end
        5088: begin
            cosine_reg0 <= 36'sb110100000111100010101101100111011101;
            sine_reg0   <= 36'sb11101101101100101001001100010001101;
        end
        5089: begin
            cosine_reg0 <= 36'sb110100000110110100000010110110011001;
            sine_reg0   <= 36'sb11101101101010010011110011100000001;
        end
        5090: begin
            cosine_reg0 <= 36'sb110100000110000101011000100010101100;
            sine_reg0   <= 36'sb11101101100111111110010001100100001;
        end
        5091: begin
            cosine_reg0 <= 36'sb110100000101010110101110101100010111;
            sine_reg0   <= 36'sb11101101100101101000100110011101111;
        end
        5092: begin
            cosine_reg0 <= 36'sb110100000100101000000101010011011011;
            sine_reg0   <= 36'sb11101101100011010010110010001101100;
        end
        5093: begin
            cosine_reg0 <= 36'sb110100000011111001011100010111111011;
            sine_reg0   <= 36'sb11101101100000111100110100110010111;
        end
        5094: begin
            cosine_reg0 <= 36'sb110100000011001010110011111001111000;
            sine_reg0   <= 36'sb11101101011110100110101110001110001;
        end
        5095: begin
            cosine_reg0 <= 36'sb110100000010011100001011111001010101;
            sine_reg0   <= 36'sb11101101011100010000011110011111101;
        end
        5096: begin
            cosine_reg0 <= 36'sb110100000001101101100100010110010010;
            sine_reg0   <= 36'sb11101101011001111010000101100111001;
        end
        5097: begin
            cosine_reg0 <= 36'sb110100000000111110111101010000110010;
            sine_reg0   <= 36'sb11101101010111100011100011100100111;
        end
        5098: begin
            cosine_reg0 <= 36'sb110100000000010000010110101000110111;
            sine_reg0   <= 36'sb11101101010101001100111000011000111;
        end
        5099: begin
            cosine_reg0 <= 36'sb110011111111100001110000011110100010;
            sine_reg0   <= 36'sb11101101010010110110000100000011011;
        end
        5100: begin
            cosine_reg0 <= 36'sb110011111110110011001010110001110101;
            sine_reg0   <= 36'sb11101101010000011111000110100100011;
        end
        5101: begin
            cosine_reg0 <= 36'sb110011111110000100100101100010110010;
            sine_reg0   <= 36'sb11101101001110000111111111111011111;
        end
        5102: begin
            cosine_reg0 <= 36'sb110011111101010110000000110001011011;
            sine_reg0   <= 36'sb11101101001011110000110000001010001;
        end
        5103: begin
            cosine_reg0 <= 36'sb110011111100100111011100011101110001;
            sine_reg0   <= 36'sb11101101001001011001010111001111010;
        end
        5104: begin
            cosine_reg0 <= 36'sb110011111011111000111000100111110111;
            sine_reg0   <= 36'sb11101101000111000001110101001011001;
        end
        5105: begin
            cosine_reg0 <= 36'sb110011111011001010010101001111101101;
            sine_reg0   <= 36'sb11101101000100101010001001111101111;
        end
        5106: begin
            cosine_reg0 <= 36'sb110011111010011011110010010101010111;
            sine_reg0   <= 36'sb11101101000010010010010101100111111;
        end
        5107: begin
            cosine_reg0 <= 36'sb110011111001101101001111111000110101;
            sine_reg0   <= 36'sb11101100111111111010011000001000111;
        end
        5108: begin
            cosine_reg0 <= 36'sb110011111000111110101101111010001010;
            sine_reg0   <= 36'sb11101100111101100010010001100001001;
        end
        5109: begin
            cosine_reg0 <= 36'sb110011111000010000001100011001010111;
            sine_reg0   <= 36'sb11101100111011001010000001110000101;
        end
        5110: begin
            cosine_reg0 <= 36'sb110011110111100001101011010110011110;
            sine_reg0   <= 36'sb11101100111000110001101000110111101;
        end
        5111: begin
            cosine_reg0 <= 36'sb110011110110110011001010110001100001;
            sine_reg0   <= 36'sb11101100110110011001000110110110001;
        end
        5112: begin
            cosine_reg0 <= 36'sb110011110110000100101010101010100010;
            sine_reg0   <= 36'sb11101100110100000000011011101100010;
        end
        5113: begin
            cosine_reg0 <= 36'sb110011110101010110001011000001100010;
            sine_reg0   <= 36'sb11101100110001100111100111011010000;
        end
        5114: begin
            cosine_reg0 <= 36'sb110011110100100111101011110110100011;
            sine_reg0   <= 36'sb11101100101111001110101001111111101;
        end
        5115: begin
            cosine_reg0 <= 36'sb110011110011111001001101001001101000;
            sine_reg0   <= 36'sb11101100101100110101100011011101000;
        end
        5116: begin
            cosine_reg0 <= 36'sb110011110011001010101110111010110001;
            sine_reg0   <= 36'sb11101100101010011100010011110010011;
        end
        5117: begin
            cosine_reg0 <= 36'sb110011110010011100010001001010000001;
            sine_reg0   <= 36'sb11101100101000000010111010111111111;
        end
        5118: begin
            cosine_reg0 <= 36'sb110011110001101101110011110111011001;
            sine_reg0   <= 36'sb11101100100101101001011001000101100;
        end
        5119: begin
            cosine_reg0 <= 36'sb110011110000111111010111000010111100;
            sine_reg0   <= 36'sb11101100100011001111101110000011010;
        end
        5120: begin
            cosine_reg0 <= 36'sb110011110000010000111010101100101011;
            sine_reg0   <= 36'sb11101100100000110101111001111001100;
        end
        5121: begin
            cosine_reg0 <= 36'sb110011101111100010011110110100100111;
            sine_reg0   <= 36'sb11101100011110011011111100101000001;
        end
        5122: begin
            cosine_reg0 <= 36'sb110011101110110100000011011010110011;
            sine_reg0   <= 36'sb11101100011100000001110110001111010;
        end
        5123: begin
            cosine_reg0 <= 36'sb110011101110000101101000011111010000;
            sine_reg0   <= 36'sb11101100011001100111100110101110111;
        end
        5124: begin
            cosine_reg0 <= 36'sb110011101101010111001110000010000001;
            sine_reg0   <= 36'sb11101100010111001101001110000111011;
        end
        5125: begin
            cosine_reg0 <= 36'sb110011101100101000110100000011000110;
            sine_reg0   <= 36'sb11101100010100110010101100011000101;
        end
        5126: begin
            cosine_reg0 <= 36'sb110011101011111010011010100010100010;
            sine_reg0   <= 36'sb11101100010010011000000001100010110;
        end
        5127: begin
            cosine_reg0 <= 36'sb110011101011001100000001100000010111;
            sine_reg0   <= 36'sb11101100001111111101001101100101111;
        end
        5128: begin
            cosine_reg0 <= 36'sb110011101010011101101000111100100110;
            sine_reg0   <= 36'sb11101100001101100010010000100010000;
        end
        5129: begin
            cosine_reg0 <= 36'sb110011101001101111010000110111010001;
            sine_reg0   <= 36'sb11101100001011000111001010010111011;
        end
        5130: begin
            cosine_reg0 <= 36'sb110011101001000000111001010000011010;
            sine_reg0   <= 36'sb11101100001000101011111011000110000;
        end
        5131: begin
            cosine_reg0 <= 36'sb110011101000010010100010001000000010;
            sine_reg0   <= 36'sb11101100000110010000100010101110000;
        end
        5132: begin
            cosine_reg0 <= 36'sb110011100111100100001011011110001100;
            sine_reg0   <= 36'sb11101100000011110101000001001111100;
        end
        5133: begin
            cosine_reg0 <= 36'sb110011100110110101110101010010111010;
            sine_reg0   <= 36'sb11101100000001011001010110101010100;
        end
        5134: begin
            cosine_reg0 <= 36'sb110011100110000111011111100110001100;
            sine_reg0   <= 36'sb11101011111110111101100010111111001;
        end
        5135: begin
            cosine_reg0 <= 36'sb110011100101011001001010011000000101;
            sine_reg0   <= 36'sb11101011111100100001100110001101100;
        end
        5136: begin
            cosine_reg0 <= 36'sb110011100100101010110101101000100111;
            sine_reg0   <= 36'sb11101011111010000101100000010101101;
        end
        5137: begin
            cosine_reg0 <= 36'sb110011100011111100100001010111110100;
            sine_reg0   <= 36'sb11101011110111101001010001010111110;
        end
        5138: begin
            cosine_reg0 <= 36'sb110011100011001110001101100101101100;
            sine_reg0   <= 36'sb11101011110101001100111001010011111;
        end
        5139: begin
            cosine_reg0 <= 36'sb110011100010011111111010010010010010;
            sine_reg0   <= 36'sb11101011110010110000011000001010001;
        end
        5140: begin
            cosine_reg0 <= 36'sb110011100001110001100111011101101001;
            sine_reg0   <= 36'sb11101011110000010011101101111010101;
        end
        5141: begin
            cosine_reg0 <= 36'sb110011100001000011010101000111110000;
            sine_reg0   <= 36'sb11101011101101110110111010100101011;
        end
        5142: begin
            cosine_reg0 <= 36'sb110011100000010101000011010000101011;
            sine_reg0   <= 36'sb11101011101011011001111110001010100;
        end
        5143: begin
            cosine_reg0 <= 36'sb110011011111100110110001111000011011;
            sine_reg0   <= 36'sb11101011101000111100111000101010000;
        end
        5144: begin
            cosine_reg0 <= 36'sb110011011110111000100000111111000010;
            sine_reg0   <= 36'sb11101011100110011111101010000100010;
        end
        5145: begin
            cosine_reg0 <= 36'sb110011011110001010010000100100100010;
            sine_reg0   <= 36'sb11101011100100000010010010011001001;
        end
        5146: begin
            cosine_reg0 <= 36'sb110011011101011100000000101000111100;
            sine_reg0   <= 36'sb11101011100001100100110001101000110;
        end
        5147: begin
            cosine_reg0 <= 36'sb110011011100101101110001001100010011;
            sine_reg0   <= 36'sb11101011011111000111000111110011010;
        end
        5148: begin
            cosine_reg0 <= 36'sb110011011011111111100010001110100111;
            sine_reg0   <= 36'sb11101011011100101001010100111000110;
        end
        5149: begin
            cosine_reg0 <= 36'sb110011011011010001010011101111111011;
            sine_reg0   <= 36'sb11101011011010001011011000111001010;
        end
        5150: begin
            cosine_reg0 <= 36'sb110011011010100011000101110000010001;
            sine_reg0   <= 36'sb11101011010111101101010011110101000;
        end
        5151: begin
            cosine_reg0 <= 36'sb110011011001110100111000001111101010;
            sine_reg0   <= 36'sb11101011010101001111000101101011111;
        end
        5152: begin
            cosine_reg0 <= 36'sb110011011001000110101011001110001001;
            sine_reg0   <= 36'sb11101011010010110000101110011110010;
        end
        5153: begin
            cosine_reg0 <= 36'sb110011011000011000011110101011101110;
            sine_reg0   <= 36'sb11101011010000010010001110001011111;
        end
        5154: begin
            cosine_reg0 <= 36'sb110011010111101010010010101000011100;
            sine_reg0   <= 36'sb11101011001101110011100100110101001;
        end
        5155: begin
            cosine_reg0 <= 36'sb110011010110111100000111000100010101;
            sine_reg0   <= 36'sb11101011001011010100110010011010000;
        end
        5156: begin
            cosine_reg0 <= 36'sb110011010110001101111011111111011001;
            sine_reg0   <= 36'sb11101011001000110101110110111010101;
        end
        5157: begin
            cosine_reg0 <= 36'sb110011010101011111110001011001101100;
            sine_reg0   <= 36'sb11101011000110010110110010010111000;
        end
        5158: begin
            cosine_reg0 <= 36'sb110011010100110001100111010011001111;
            sine_reg0   <= 36'sb11101011000011110111100100101111011;
        end
        5159: begin
            cosine_reg0 <= 36'sb110011010100000011011101101100000011;
            sine_reg0   <= 36'sb11101011000001011000001110000011110;
        end
        5160: begin
            cosine_reg0 <= 36'sb110011010011010101010100100100001011;
            sine_reg0   <= 36'sb11101010111110111000101110010100001;
        end
        5161: begin
            cosine_reg0 <= 36'sb110011010010100111001011111011101000;
            sine_reg0   <= 36'sb11101010111100011001000101100000110;
        end
        5162: begin
            cosine_reg0 <= 36'sb110011010001111001000011110010011100;
            sine_reg0   <= 36'sb11101010111001111001010011101001110;
        end
        5163: begin
            cosine_reg0 <= 36'sb110011010001001010111100001000101000;
            sine_reg0   <= 36'sb11101010110111011001011000101111001;
        end
        5164: begin
            cosine_reg0 <= 36'sb110011010000011100110100111110001111;
            sine_reg0   <= 36'sb11101010110100111001010100110001000;
        end
        5165: begin
            cosine_reg0 <= 36'sb110011001111101110101110010011010011;
            sine_reg0   <= 36'sb11101010110010011001000111101111011;
        end
        5166: begin
            cosine_reg0 <= 36'sb110011001111000000101000000111110100;
            sine_reg0   <= 36'sb11101010101111111000110001101010100;
        end
        5167: begin
            cosine_reg0 <= 36'sb110011001110010010100010011011110101;
            sine_reg0   <= 36'sb11101010101101011000010010100010011;
        end
        5168: begin
            cosine_reg0 <= 36'sb110011001101100100011101001111011000;
            sine_reg0   <= 36'sb11101010101010110111101010010111001;
        end
        5169: begin
            cosine_reg0 <= 36'sb110011001100110110011000100010011110;
            sine_reg0   <= 36'sb11101010101000010110111001001000111;
        end
        5170: begin
            cosine_reg0 <= 36'sb110011001100001000010100010101001010;
            sine_reg0   <= 36'sb11101010100101110101111110110111110;
        end
        5171: begin
            cosine_reg0 <= 36'sb110011001011011010010000100111011100;
            sine_reg0   <= 36'sb11101010100011010100111011100011110;
        end
        5172: begin
            cosine_reg0 <= 36'sb110011001010101100001101011001010111;
            sine_reg0   <= 36'sb11101010100000110011101111001101000;
        end
        5173: begin
            cosine_reg0 <= 36'sb110011001001111110001010101010111101;
            sine_reg0   <= 36'sb11101010011110010010011001110011101;
        end
        5174: begin
            cosine_reg0 <= 36'sb110011001001010000001000011100001111;
            sine_reg0   <= 36'sb11101010011011110000111011010111110;
        end
        5175: begin
            cosine_reg0 <= 36'sb110011001000100010000110101101001111;
            sine_reg0   <= 36'sb11101010011001001111010011111001011;
        end
        5176: begin
            cosine_reg0 <= 36'sb110011000111110100000101011101111111;
            sine_reg0   <= 36'sb11101010010110101101100011011000101;
        end
        5177: begin
            cosine_reg0 <= 36'sb110011000111000110000100101110100000;
            sine_reg0   <= 36'sb11101010010100001011101001110101110;
        end
        5178: begin
            cosine_reg0 <= 36'sb110011000110011000000100011110110101;
            sine_reg0   <= 36'sb11101010010001101001100111010000101;
        end
        5179: begin
            cosine_reg0 <= 36'sb110011000101101010000100101110111111;
            sine_reg0   <= 36'sb11101010001111000111011011101001100;
        end
        5180: begin
            cosine_reg0 <= 36'sb110011000100111100000101011110111111;
            sine_reg0   <= 36'sb11101010001100100101000111000000011;
        end
        5181: begin
            cosine_reg0 <= 36'sb110011000100001110000110101110111001;
            sine_reg0   <= 36'sb11101010001010000010101001010101011;
        end
        5182: begin
            cosine_reg0 <= 36'sb110011000011100000001000011110101101;
            sine_reg0   <= 36'sb11101010000111100000000010101000101;
        end
        5183: begin
            cosine_reg0 <= 36'sb110011000010110010001010101110011101;
            sine_reg0   <= 36'sb11101010000100111101010010111010010;
        end
        5184: begin
            cosine_reg0 <= 36'sb110011000010000100001101011110001011;
            sine_reg0   <= 36'sb11101010000010011010011010001010011;
        end
        5185: begin
            cosine_reg0 <= 36'sb110011000001010110010000101101111001;
            sine_reg0   <= 36'sb11101001111111110111011000011000111;
        end
        5186: begin
            cosine_reg0 <= 36'sb110011000000101000010100011101101001;
            sine_reg0   <= 36'sb11101001111101010100001101100110001;
        end
        5187: begin
            cosine_reg0 <= 36'sb110010111111111010011000101101011100;
            sine_reg0   <= 36'sb11101001111010110000111001110010001;
        end
        5188: begin
            cosine_reg0 <= 36'sb110010111111001100011101011101010100;
            sine_reg0   <= 36'sb11101001111000001101011100111100111;
        end
        5189: begin
            cosine_reg0 <= 36'sb110010111110011110100010101101010010;
            sine_reg0   <= 36'sb11101001110101101001110111000110101;
        end
        5190: begin
            cosine_reg0 <= 36'sb110010111101110000101000011101011010;
            sine_reg0   <= 36'sb11101001110011000110001000001111010;
        end
        5191: begin
            cosine_reg0 <= 36'sb110010111101000010101110101101101100;
            sine_reg0   <= 36'sb11101001110000100010010000010111001;
        end
        5192: begin
            cosine_reg0 <= 36'sb110010111100010100110101011110001010;
            sine_reg0   <= 36'sb11101001101101111110001111011110010;
        end
        5193: begin
            cosine_reg0 <= 36'sb110010111011100110111100101110110110;
            sine_reg0   <= 36'sb11101001101011011010000101100100101;
        end
        5194: begin
            cosine_reg0 <= 36'sb110010111010111001000100011111110001;
            sine_reg0   <= 36'sb11101001101000110101110010101010100;
        end
        5195: begin
            cosine_reg0 <= 36'sb110010111010001011001100110000111111;
            sine_reg0   <= 36'sb11101001100110010001010110101111111;
        end
        5196: begin
            cosine_reg0 <= 36'sb110010111001011101010101100010011111;
            sine_reg0   <= 36'sb11101001100011101100110001110100111;
        end
        5197: begin
            cosine_reg0 <= 36'sb110010111000101111011110110100010100;
            sine_reg0   <= 36'sb11101001100001001000000011111001100;
        end
        5198: begin
            cosine_reg0 <= 36'sb110010111000000001101000100110100001;
            sine_reg0   <= 36'sb11101001011110100011001100111110000;
        end
        5199: begin
            cosine_reg0 <= 36'sb110010110111010011110010111001000101;
            sine_reg0   <= 36'sb11101001011011111110001101000010100;
        end
        5200: begin
            cosine_reg0 <= 36'sb110010110110100101111101101100000101;
            sine_reg0   <= 36'sb11101001011001011001000100000110111;
        end
        5201: begin
            cosine_reg0 <= 36'sb110010110101111000001000111111100000;
            sine_reg0   <= 36'sb11101001010110110011110010001011100;
        end
        5202: begin
            cosine_reg0 <= 36'sb110010110101001010010100110011011001;
            sine_reg0   <= 36'sb11101001010100001110010111010000010;
        end
        5203: begin
            cosine_reg0 <= 36'sb110010110100011100100001000111110001;
            sine_reg0   <= 36'sb11101001010001101000110011010101011;
        end
        5204: begin
            cosine_reg0 <= 36'sb110010110011101110101101111100101100;
            sine_reg0   <= 36'sb11101001001111000011000110011010111;
        end
        5205: begin
            cosine_reg0 <= 36'sb110010110011000000111011010010001001;
            sine_reg0   <= 36'sb11101001001100011101010000100000111;
        end
        5206: begin
            cosine_reg0 <= 36'sb110010110010010011001001001000001011;
            sine_reg0   <= 36'sb11101001001001110111010001100111100;
        end
        5207: begin
            cosine_reg0 <= 36'sb110010110001100101010111011110110100;
            sine_reg0   <= 36'sb11101001000111010001001001101110111;
        end
        5208: begin
            cosine_reg0 <= 36'sb110010110000110111100110010110000101;
            sine_reg0   <= 36'sb11101001000100101010111000110111001;
        end
        5209: begin
            cosine_reg0 <= 36'sb110010110000001001110101101110000000;
            sine_reg0   <= 36'sb11101001000010000100011111000000001;
        end
        5210: begin
            cosine_reg0 <= 36'sb110010101111011100000101100110101000;
            sine_reg0   <= 36'sb11101000111111011101111100001010010;
        end
        5211: begin
            cosine_reg0 <= 36'sb110010101110101110010101111111111101;
            sine_reg0   <= 36'sb11101000111100110111010000010101100;
        end
        5212: begin
            cosine_reg0 <= 36'sb110010101110000000100110111010000010;
            sine_reg0   <= 36'sb11101000111010010000011011100001111;
        end
        5213: begin
            cosine_reg0 <= 36'sb110010101101010010111000010100111000;
            sine_reg0   <= 36'sb11101000110111101001011101101111101;
        end
        5214: begin
            cosine_reg0 <= 36'sb110010101100100101001010010000100001;
            sine_reg0   <= 36'sb11101000110101000010010110111110111;
        end
        5215: begin
            cosine_reg0 <= 36'sb110010101011110111011100101100111110;
            sine_reg0   <= 36'sb11101000110010011011000111001111100;
        end
        5216: begin
            cosine_reg0 <= 36'sb110010101011001001101111101010010011;
            sine_reg0   <= 36'sb11101000101111110011101110100001111;
        end
        5217: begin
            cosine_reg0 <= 36'sb110010101010011100000011001000011111;
            sine_reg0   <= 36'sb11101000101101001100001100110101111;
        end
        5218: begin
            cosine_reg0 <= 36'sb110010101001101110010111000111100110;
            sine_reg0   <= 36'sb11101000101010100100100010001011110;
        end
        5219: begin
            cosine_reg0 <= 36'sb110010101001000000101011100111101001;
            sine_reg0   <= 36'sb11101000100111111100101110100011100;
        end
        5220: begin
            cosine_reg0 <= 36'sb110010101000010011000000101000101001;
            sine_reg0   <= 36'sb11101000100101010100110001111101010;
        end
        5221: begin
            cosine_reg0 <= 36'sb110010100111100101010110001010101000;
            sine_reg0   <= 36'sb11101000100010101100101100011001001;
        end
        5222: begin
            cosine_reg0 <= 36'sb110010100110110111101100001101101001;
            sine_reg0   <= 36'sb11101000100000000100011101110111011;
        end
        5223: begin
            cosine_reg0 <= 36'sb110010100110001010000010110001101101;
            sine_reg0   <= 36'sb11101000011101011100000110010111110;
        end
        5224: begin
            cosine_reg0 <= 36'sb110010100101011100011001110110110101;
            sine_reg0   <= 36'sb11101000011010110011100101111010110;
        end
        5225: begin
            cosine_reg0 <= 36'sb110010100100101110110001011101000011;
            sine_reg0   <= 36'sb11101000011000001010111100100000001;
        end
        5226: begin
            cosine_reg0 <= 36'sb110010100100000001001001100100011010;
            sine_reg0   <= 36'sb11101000010101100010001010001000001;
        end
        5227: begin
            cosine_reg0 <= 36'sb110010100011010011100010001100111011;
            sine_reg0   <= 36'sb11101000010010111001001110110011000;
        end
        5228: begin
            cosine_reg0 <= 36'sb110010100010100101111011010110100111;
            sine_reg0   <= 36'sb11101000010000010000001010100000101;
        end
        5229: begin
            cosine_reg0 <= 36'sb110010100001111000010101000001100001;
            sine_reg0   <= 36'sb11101000001101100110111101010001001;
        end
        5230: begin
            cosine_reg0 <= 36'sb110010100001001010101111001101101010;
            sine_reg0   <= 36'sb11101000001010111101100111000100110;
        end
        5231: begin
            cosine_reg0 <= 36'sb110010100000011101001001111011000100;
            sine_reg0   <= 36'sb11101000001000010100000111111011100;
        end
        5232: begin
            cosine_reg0 <= 36'sb110010011111101111100101001001110001;
            sine_reg0   <= 36'sb11101000000101101010011111110101100;
        end
        5233: begin
            cosine_reg0 <= 36'sb110010011111000010000000111001110010;
            sine_reg0   <= 36'sb11101000000011000000101110110010110;
        end
        5234: begin
            cosine_reg0 <= 36'sb110010011110010100011101001011001001;
            sine_reg0   <= 36'sb11101000000000010110110100110011101;
        end
        5235: begin
            cosine_reg0 <= 36'sb110010011101100110111001111101111000;
            sine_reg0   <= 36'sb11100111111101101100110001110111111;
        end
        5236: begin
            cosine_reg0 <= 36'sb110010011100111001010111010010000001;
            sine_reg0   <= 36'sb11100111111011000010100101111111111;
        end
        5237: begin
            cosine_reg0 <= 36'sb110010011100001011110101000111100110;
            sine_reg0   <= 36'sb11100111111000011000010001001011101;
        end
        5238: begin
            cosine_reg0 <= 36'sb110010011011011110010011011110101000;
            sine_reg0   <= 36'sb11100111110101101101110011011011001;
        end
        5239: begin
            cosine_reg0 <= 36'sb110010011010110000110010010111001000;
            sine_reg0   <= 36'sb11100111110011000011001100101110110;
        end
        5240: begin
            cosine_reg0 <= 36'sb110010011010000011010001110001001010;
            sine_reg0   <= 36'sb11100111110000011000011101000110011;
        end
        5241: begin
            cosine_reg0 <= 36'sb110010011001010101110001101100101110;
            sine_reg0   <= 36'sb11100111101101101101100100100010001;
        end
        5242: begin
            cosine_reg0 <= 36'sb110010011000101000010010001001110110;
            sine_reg0   <= 36'sb11100111101011000010100011000010001;
        end
        5243: begin
            cosine_reg0 <= 36'sb110010010111111010110011001000100101;
            sine_reg0   <= 36'sb11100111101000010111011000100110100;
        end
        5244: begin
            cosine_reg0 <= 36'sb110010010111001101010100101000111011;
            sine_reg0   <= 36'sb11100111100101101100000101001111100;
        end
        5245: begin
            cosine_reg0 <= 36'sb110010010110011111110110101010111011;
            sine_reg0   <= 36'sb11100111100011000000101000111100111;
        end
        5246: begin
            cosine_reg0 <= 36'sb110010010101110010011001001110100110;
            sine_reg0   <= 36'sb11100111100000010101000011101111000;
        end
        5247: begin
            cosine_reg0 <= 36'sb110010010101000100111100010011111101;
            sine_reg0   <= 36'sb11100111011101101001010101100110000;
        end
        5248: begin
            cosine_reg0 <= 36'sb110010010100010111011111111011000100;
            sine_reg0   <= 36'sb11100111011010111101011110100001110;
        end
        5249: begin
            cosine_reg0 <= 36'sb110010010011101010000100000011111100;
            sine_reg0   <= 36'sb11100111011000010001011110100010101;
        end
        5250: begin
            cosine_reg0 <= 36'sb110010010010111100101000101110100101;
            sine_reg0   <= 36'sb11100111010101100101010101101000100;
        end
        5251: begin
            cosine_reg0 <= 36'sb110010010010001111001101111011000011;
            sine_reg0   <= 36'sb11100111010010111001000011110011101;
        end
        5252: begin
            cosine_reg0 <= 36'sb110010010001100001110011101001010110;
            sine_reg0   <= 36'sb11100111010000001100101001000100000;
        end
        5253: begin
            cosine_reg0 <= 36'sb110010010000110100011001111001100001;
            sine_reg0   <= 36'sb11100111001101100000000101011001110;
        end
        5254: begin
            cosine_reg0 <= 36'sb110010010000000111000000101011100101;
            sine_reg0   <= 36'sb11100111001010110011011000110101001;
        end
        5255: begin
            cosine_reg0 <= 36'sb110010001111011001100111111111100101;
            sine_reg0   <= 36'sb11100111001000000110100011010110000;
        end
        5256: begin
            cosine_reg0 <= 36'sb110010001110101100001111110101100001;
            sine_reg0   <= 36'sb11100111000101011001100100111100110;
        end
        5257: begin
            cosine_reg0 <= 36'sb110010001101111110111000001101011011;
            sine_reg0   <= 36'sb11100111000010101100011101101001001;
        end
        5258: begin
            cosine_reg0 <= 36'sb110010001101010001100001000111010110;
            sine_reg0   <= 36'sb11100110111111111111001101011011100;
        end
        5259: begin
            cosine_reg0 <= 36'sb110010001100100100001010100011010011;
            sine_reg0   <= 36'sb11100110111101010001110100010100000;
        end
        5260: begin
            cosine_reg0 <= 36'sb110010001011110110110100100001010100;
            sine_reg0   <= 36'sb11100110111010100100010010010010100;
        end
        5261: begin
            cosine_reg0 <= 36'sb110010001011001001011111000001011010;
            sine_reg0   <= 36'sb11100110110111110110100111010111011;
        end
        5262: begin
            cosine_reg0 <= 36'sb110010001010011100001010000011101000;
            sine_reg0   <= 36'sb11100110110101001000110011100010100;
        end
        5263: begin
            cosine_reg0 <= 36'sb110010001001101110110101100111111110;
            sine_reg0   <= 36'sb11100110110010011010110110110100001;
        end
        5264: begin
            cosine_reg0 <= 36'sb110010001001000001100001101110100000;
            sine_reg0   <= 36'sb11100110101111101100110001001100010;
        end
        5265: begin
            cosine_reg0 <= 36'sb110010001000010100001110010111001110;
            sine_reg0   <= 36'sb11100110101100111110100010101011000;
        end
        5266: begin
            cosine_reg0 <= 36'sb110010000111100110111011100010001010;
            sine_reg0   <= 36'sb11100110101010010000001011010000101;
        end
        5267: begin
            cosine_reg0 <= 36'sb110010000110111001101001001111010110;
            sine_reg0   <= 36'sb11100110100111100001101010111101000;
        end
        5268: begin
            cosine_reg0 <= 36'sb110010000110001100010111011110110100;
            sine_reg0   <= 36'sb11100110100100110011000001110000100;
        end
        5269: begin
            cosine_reg0 <= 36'sb110010000101011111000110010000100110;
            sine_reg0   <= 36'sb11100110100010000100001111101011000;
        end
        5270: begin
            cosine_reg0 <= 36'sb110010000100110001110101100100101100;
            sine_reg0   <= 36'sb11100110011111010101010100101100101;
        end
        5271: begin
            cosine_reg0 <= 36'sb110010000100000100100101011011001010;
            sine_reg0   <= 36'sb11100110011100100110010000110101101;
        end
        5272: begin
            cosine_reg0 <= 36'sb110010000011010111010101110100000000;
            sine_reg0   <= 36'sb11100110011001110111000100000110000;
        end
        5273: begin
            cosine_reg0 <= 36'sb110010000010101010000110101111010001;
            sine_reg0   <= 36'sb11100110010111000111101110011101111;
        end
        5274: begin
            cosine_reg0 <= 36'sb110010000001111100111000001100111111;
            sine_reg0   <= 36'sb11100110010100011000001111111101010;
        end
        5275: begin
            cosine_reg0 <= 36'sb110010000001001111101010001101001010;
            sine_reg0   <= 36'sb11100110010001101000101000100100100;
        end
        5276: begin
            cosine_reg0 <= 36'sb110010000000100010011100101111110101;
            sine_reg0   <= 36'sb11100110001110111000111000010011100;
        end
        5277: begin
            cosine_reg0 <= 36'sb110001111111110101001111110101000001;
            sine_reg0   <= 36'sb11100110001100001000111111001010011;
        end
        5278: begin
            cosine_reg0 <= 36'sb110001111111001000000011011100110001;
            sine_reg0   <= 36'sb11100110001001011000111101001001011;
        end
        5279: begin
            cosine_reg0 <= 36'sb110001111110011010110111100111000101;
            sine_reg0   <= 36'sb11100110000110101000110010010000100;
        end
        5280: begin
            cosine_reg0 <= 36'sb110001111101101101101100010100000000;
            sine_reg0   <= 36'sb11100110000011111000011110011111110;
        end
        5281: begin
            cosine_reg0 <= 36'sb110001111101000000100001100011100100;
            sine_reg0   <= 36'sb11100110000001001000000001110111100;
        end
        5282: begin
            cosine_reg0 <= 36'sb110001111100010011010111010101110010;
            sine_reg0   <= 36'sb11100101111110010111011100010111101;
        end
        5283: begin
            cosine_reg0 <= 36'sb110001111011100110001101101010101011;
            sine_reg0   <= 36'sb11100101111011100110101110000000010;
        end
        5284: begin
            cosine_reg0 <= 36'sb110001111010111001000100100010010011;
            sine_reg0   <= 36'sb11100101111000110101110110110001101;
        end
        5285: begin
            cosine_reg0 <= 36'sb110001111010001011111011111100101010;
            sine_reg0   <= 36'sb11100101110110000100110110101011110;
        end
        5286: begin
            cosine_reg0 <= 36'sb110001111001011110110011111001110001;
            sine_reg0   <= 36'sb11100101110011010011101101101110111;
        end
        5287: begin
            cosine_reg0 <= 36'sb110001111000110001101100011001101100;
            sine_reg0   <= 36'sb11100101110000100010011011111010111;
        end
        5288: begin
            cosine_reg0 <= 36'sb110001111000000100100101011100011100;
            sine_reg0   <= 36'sb11100101101101110001000001001111111;
        end
        5289: begin
            cosine_reg0 <= 36'sb110001110111010111011111000010000001;
            sine_reg0   <= 36'sb11100101101010111111011101101110010;
        end
        5290: begin
            cosine_reg0 <= 36'sb110001110110101010011001001010011111;
            sine_reg0   <= 36'sb11100101101000001101110001010101111;
        end
        5291: begin
            cosine_reg0 <= 36'sb110001110101111101010011110101110111;
            sine_reg0   <= 36'sb11100101100101011011111100000110111;
        end
        5292: begin
            cosine_reg0 <= 36'sb110001110101010000001111000100001010;
            sine_reg0   <= 36'sb11100101100010101001111110000001011;
        end
        5293: begin
            cosine_reg0 <= 36'sb110001110100100011001010110101011011;
            sine_reg0   <= 36'sb11100101011111110111110111000101100;
        end
        5294: begin
            cosine_reg0 <= 36'sb110001110011110110000111001001101010;
            sine_reg0   <= 36'sb11100101011101000101100111010011100;
        end
        5295: begin
            cosine_reg0 <= 36'sb110001110011001001000100000000111011;
            sine_reg0   <= 36'sb11100101011010010011001110101011010;
        end
        5296: begin
            cosine_reg0 <= 36'sb110001110010011100000001011011001110;
            sine_reg0   <= 36'sb11100101010111100000101101001100111;
        end
        5297: begin
            cosine_reg0 <= 36'sb110001110001101110111111011000100101;
            sine_reg0   <= 36'sb11100101010100101110000010111000101;
        end
        5298: begin
            cosine_reg0 <= 36'sb110001110001000001111101111001000010;
            sine_reg0   <= 36'sb11100101010001111011001111101110101;
        end
        5299: begin
            cosine_reg0 <= 36'sb110001110000010100111100111100100111;
            sine_reg0   <= 36'sb11100101001111001000010011101110110;
        end
        5300: begin
            cosine_reg0 <= 36'sb110001101111100111111100100011010101;
            sine_reg0   <= 36'sb11100101001100010101001110111001011;
        end
        5301: begin
            cosine_reg0 <= 36'sb110001101110111010111100101101001111;
            sine_reg0   <= 36'sb11100101001001100010000001001110100;
        end
        5302: begin
            cosine_reg0 <= 36'sb110001101110001101111101011010010101;
            sine_reg0   <= 36'sb11100101000110101110101010101110001;
        end
        5303: begin
            cosine_reg0 <= 36'sb110001101101100000111110101010101010;
            sine_reg0   <= 36'sb11100101000011111011001011011000100;
        end
        5304: begin
            cosine_reg0 <= 36'sb110001101100110100000000011110010000;
            sine_reg0   <= 36'sb11100101000001000111100011001101110;
        end
        5305: begin
            cosine_reg0 <= 36'sb110001101100000111000010110101000111;
            sine_reg0   <= 36'sb11100100111110010011110010001101110;
        end
        5306: begin
            cosine_reg0 <= 36'sb110001101011011010000101101111010011;
            sine_reg0   <= 36'sb11100100111011011111111000011001000;
        end
        5307: begin
            cosine_reg0 <= 36'sb110001101010101101001001001100110100;
            sine_reg0   <= 36'sb11100100111000101011110101101111010;
        end
        5308: begin
            cosine_reg0 <= 36'sb110001101010000000001101001101101100;
            sine_reg0   <= 36'sb11100100110101110111101010010000110;
        end
        5309: begin
            cosine_reg0 <= 36'sb110001101001010011010001110001111110;
            sine_reg0   <= 36'sb11100100110011000011010101111101101;
        end
        5310: begin
            cosine_reg0 <= 36'sb110001101000100110010110111001101010;
            sine_reg0   <= 36'sb11100100110000001110111000110110000;
        end
        5311: begin
            cosine_reg0 <= 36'sb110001100111111001011100100100110011;
            sine_reg0   <= 36'sb11100100101101011010010010111001111;
        end
        5312: begin
            cosine_reg0 <= 36'sb110001100111001100100010110011011010;
            sine_reg0   <= 36'sb11100100101010100101100100001001100;
        end
        5313: begin
            cosine_reg0 <= 36'sb110001100110011111101001100101100001;
            sine_reg0   <= 36'sb11100100100111110000101100100100111;
        end
        5314: begin
            cosine_reg0 <= 36'sb110001100101110010110000111011001010;
            sine_reg0   <= 36'sb11100100100100111011101100001100010;
        end
        5315: begin
            cosine_reg0 <= 36'sb110001100101000101111000110100010110;
            sine_reg0   <= 36'sb11100100100010000110100010111111100;
        end
        5316: begin
            cosine_reg0 <= 36'sb110001100100011001000001010001001000;
            sine_reg0   <= 36'sb11100100011111010001010000111110111;
        end
        5317: begin
            cosine_reg0 <= 36'sb110001100011101100001010010001100000;
            sine_reg0   <= 36'sb11100100011100011011110110001010101;
        end
        5318: begin
            cosine_reg0 <= 36'sb110001100010111111010011110101100001;
            sine_reg0   <= 36'sb11100100011001100110010010100010100;
        end
        5319: begin
            cosine_reg0 <= 36'sb110001100010010010011101111101001101;
            sine_reg0   <= 36'sb11100100010110110000100110000111000;
        end
        5320: begin
            cosine_reg0 <= 36'sb110001100001100101101000101000100100;
            sine_reg0   <= 36'sb11100100010011111010110000111000000;
        end
        5321: begin
            cosine_reg0 <= 36'sb110001100000111000110011110111101010;
            sine_reg0   <= 36'sb11100100010001000100110010110101101;
        end
        5322: begin
            cosine_reg0 <= 36'sb110001100000001011111111101010011110;
            sine_reg0   <= 36'sb11100100001110001110101100000000000;
        end
        5323: begin
            cosine_reg0 <= 36'sb110001011111011111001100000001000101;
            sine_reg0   <= 36'sb11100100001011011000011100010111011;
        end
        5324: begin
            cosine_reg0 <= 36'sb110001011110110010011000111011011110;
            sine_reg0   <= 36'sb11100100001000100010000011111011101;
        end
        5325: begin
            cosine_reg0 <= 36'sb110001011110000101100110011001101100;
            sine_reg0   <= 36'sb11100100000101101011100010101101000;
        end
        5326: begin
            cosine_reg0 <= 36'sb110001011101011000110100011011110000;
            sine_reg0   <= 36'sb11100100000010110100111000101011101;
        end
        5327: begin
            cosine_reg0 <= 36'sb110001011100101100000011000001101101;
            sine_reg0   <= 36'sb11100011111111111110000101110111101;
        end
        5328: begin
            cosine_reg0 <= 36'sb110001011011111111010010001011100011;
            sine_reg0   <= 36'sb11100011111101000111001010010001000;
        end
        5329: begin
            cosine_reg0 <= 36'sb110001011011010010100001111001010101;
            sine_reg0   <= 36'sb11100011111010010000000101110111111;
        end
        5330: begin
            cosine_reg0 <= 36'sb110001011010100101110010001011000101;
            sine_reg0   <= 36'sb11100011110111011000111000101100100;
        end
        5331: begin
            cosine_reg0 <= 36'sb110001011001111001000011000000110100;
            sine_reg0   <= 36'sb11100011110100100001100010101110111;
        end
        5332: begin
            cosine_reg0 <= 36'sb110001011001001100010100011010100011;
            sine_reg0   <= 36'sb11100011110001101010000011111111000;
        end
        5333: begin
            cosine_reg0 <= 36'sb110001011000011111100110011000010101;
            sine_reg0   <= 36'sb11100011101110110010011100011101010;
        end
        5334: begin
            cosine_reg0 <= 36'sb110001010111110010111000111010001011;
            sine_reg0   <= 36'sb11100011101011111010101100001001100;
        end
        5335: begin
            cosine_reg0 <= 36'sb110001010111000110001100000000000111;
            sine_reg0   <= 36'sb11100011101001000010110011000100000;
        end
        5336: begin
            cosine_reg0 <= 36'sb110001010110011001011111101010001011;
            sine_reg0   <= 36'sb11100011100110001010110001001100111;
        end
        5337: begin
            cosine_reg0 <= 36'sb110001010101101100110011111000011001;
            sine_reg0   <= 36'sb11100011100011010010100110100100001;
        end
        5338: begin
            cosine_reg0 <= 36'sb110001010101000000001000101010110001;
            sine_reg0   <= 36'sb11100011100000011010010011001001111;
        end
        5339: begin
            cosine_reg0 <= 36'sb110001010100010011011110000001010111;
            sine_reg0   <= 36'sb11100011011101100001110110111110011;
        end
        5340: begin
            cosine_reg0 <= 36'sb110001010011100110110011111100001011;
            sine_reg0   <= 36'sb11100011011010101001010010000001100;
        end
        5341: begin
            cosine_reg0 <= 36'sb110001010010111010001010011011001111;
            sine_reg0   <= 36'sb11100011010111110000100100010011101;
        end
        5342: begin
            cosine_reg0 <= 36'sb110001010010001101100001011110100110;
            sine_reg0   <= 36'sb11100011010100110111101101110100101;
        end
        5343: begin
            cosine_reg0 <= 36'sb110001010001100000111001000110010000;
            sine_reg0   <= 36'sb11100011010001111110101110100100110;
        end
        5344: begin
            cosine_reg0 <= 36'sb110001010000110100010001010010010000;
            sine_reg0   <= 36'sb11100011001111000101100110100100001;
        end
        5345: begin
            cosine_reg0 <= 36'sb110001010000000111101010000010100111;
            sine_reg0   <= 36'sb11100011001100001100010101110010111;
        end
        5346: begin
            cosine_reg0 <= 36'sb110001001111011011000011010111010110;
            sine_reg0   <= 36'sb11100011001001010010111100010000111;
        end
        5347: begin
            cosine_reg0 <= 36'sb110001001110101110011101010000100001;
            sine_reg0   <= 36'sb11100011000110011001011001111110101;
        end
        5348: begin
            cosine_reg0 <= 36'sb110001001110000001110111101110001000;
            sine_reg0   <= 36'sb11100011000011011111101110111011111;
        end
        5349: begin
            cosine_reg0 <= 36'sb110001001101010101010010110000001101;
            sine_reg0   <= 36'sb11100011000000100101111011001001000;
        end
        5350: begin
            cosine_reg0 <= 36'sb110001001100101000101110010110110001;
            sine_reg0   <= 36'sb11100010111101101011111110100101111;
        end
        5351: begin
            cosine_reg0 <= 36'sb110001001011111100001010100001111000;
            sine_reg0   <= 36'sb11100010111010110001111001010010111;
        end
        5352: begin
            cosine_reg0 <= 36'sb110001001011001111100111010001100001;
            sine_reg0   <= 36'sb11100010110111110111101011001111111;
        end
        5353: begin
            cosine_reg0 <= 36'sb110001001010100011000100100101110000;
            sine_reg0   <= 36'sb11100010110100111101010100011101001;
        end
        5354: begin
            cosine_reg0 <= 36'sb110001001001110110100010011110100101;
            sine_reg0   <= 36'sb11100010110010000010110100111010101;
        end
        5355: begin
            cosine_reg0 <= 36'sb110001001001001010000000111100000010;
            sine_reg0   <= 36'sb11100010101111001000001100101000101;
        end
        5356: begin
            cosine_reg0 <= 36'sb110001001000011101011111111110001010;
            sine_reg0   <= 36'sb11100010101100001101011011100111010;
        end
        5357: begin
            cosine_reg0 <= 36'sb110001000111110000111111100100111110;
            sine_reg0   <= 36'sb11100010101001010010100001110110100;
        end
        5358: begin
            cosine_reg0 <= 36'sb110001000111000100011111110000011111;
            sine_reg0   <= 36'sb11100010100110010111011111010110100;
        end
        5359: begin
            cosine_reg0 <= 36'sb110001000110011000000000100000101111;
            sine_reg0   <= 36'sb11100010100011011100010100000111011;
        end
        5360: begin
            cosine_reg0 <= 36'sb110001000101101011100001110101110000;
            sine_reg0   <= 36'sb11100010100000100001000000001001010;
        end
        5361: begin
            cosine_reg0 <= 36'sb110001000100111111000011101111100100;
            sine_reg0   <= 36'sb11100010011101100101100011011100010;
        end
        5362: begin
            cosine_reg0 <= 36'sb110001000100010010100110001110001101;
            sine_reg0   <= 36'sb11100010011010101001111110000000100;
        end
        5363: begin
            cosine_reg0 <= 36'sb110001000011100110001001010001101011;
            sine_reg0   <= 36'sb11100010010111101110001111110110000;
        end
        5364: begin
            cosine_reg0 <= 36'sb110001000010111001101100111010000001;
            sine_reg0   <= 36'sb11100010010100110010011000111101001;
        end
        5365: begin
            cosine_reg0 <= 36'sb110001000010001101010001000111010001;
            sine_reg0   <= 36'sb11100010010001110110011001010101101;
        end
        5366: begin
            cosine_reg0 <= 36'sb110001000001100000110101111001011100;
            sine_reg0   <= 36'sb11100010001110111010010000111111111;
        end
        5367: begin
            cosine_reg0 <= 36'sb110001000000110100011011010000100101;
            sine_reg0   <= 36'sb11100010001011111101111111111100000;
        end
        5368: begin
            cosine_reg0 <= 36'sb110001000000001000000001001100101011;
            sine_reg0   <= 36'sb11100010001001000001100110001010000;
        end
        5369: begin
            cosine_reg0 <= 36'sb110000111111011011100111101101110010;
            sine_reg0   <= 36'sb11100010000110000101000011101001111;
        end
        5370: begin
            cosine_reg0 <= 36'sb110000111110101111001110110011111100;
            sine_reg0   <= 36'sb11100010000011001000011000011100000;
        end
        5371: begin
            cosine_reg0 <= 36'sb110000111110000010110110011111001001;
            sine_reg0   <= 36'sb11100010000000001011100100100000011;
        end
        5372: begin
            cosine_reg0 <= 36'sb110000111101010110011110101111011100;
            sine_reg0   <= 36'sb11100001111101001110100111110111001;
        end
        5373: begin
            cosine_reg0 <= 36'sb110000111100101010000111100100110101;
            sine_reg0   <= 36'sb11100001111010010001100010100000011;
        end
        5374: begin
            cosine_reg0 <= 36'sb110000111011111101110000111111011000;
            sine_reg0   <= 36'sb11100001110111010100010100011100001;
        end
        5375: begin
            cosine_reg0 <= 36'sb110000111011010001011010111111000110;
            sine_reg0   <= 36'sb11100001110100010110111101101010101;
        end
        5376: begin
            cosine_reg0 <= 36'sb110000111010100101000101100100000000;
            sine_reg0   <= 36'sb11100001110001011001011110001011111;
        end
        5377: begin
            cosine_reg0 <= 36'sb110000111001111000110000101110001000;
            sine_reg0   <= 36'sb11100001101110011011110110000000001;
        end
        5378: begin
            cosine_reg0 <= 36'sb110000111001001100011100011101011111;
            sine_reg0   <= 36'sb11100001101011011110000101000111011;
        end
        5379: begin
            cosine_reg0 <= 36'sb110000111000100000001000110010001001;
            sine_reg0   <= 36'sb11100001101000100000001011100001111;
        end
        5380: begin
            cosine_reg0 <= 36'sb110000110111110011110101101100000101;
            sine_reg0   <= 36'sb11100001100101100010001001001111101;
        end
        5381: begin
            cosine_reg0 <= 36'sb110000110111000111100011001011010110;
            sine_reg0   <= 36'sb11100001100010100011111110010000101;
        end
        5382: begin
            cosine_reg0 <= 36'sb110000110110011011010001001111111110;
            sine_reg0   <= 36'sb11100001011111100101101010100101010;
        end
        5383: begin
            cosine_reg0 <= 36'sb110000110101101110111111111001111111;
            sine_reg0   <= 36'sb11100001011100100111001110001101100;
        end
        5384: begin
            cosine_reg0 <= 36'sb110000110101000010101111001001011001;
            sine_reg0   <= 36'sb11100001011001101000101001001001100;
        end
        5385: begin
            cosine_reg0 <= 36'sb110000110100010110011110111110001111;
            sine_reg0   <= 36'sb11100001010110101001111011011001010;
        end
        5386: begin
            cosine_reg0 <= 36'sb110000110011101010001111011000100010;
            sine_reg0   <= 36'sb11100001010011101011000100111101000;
        end
        5387: begin
            cosine_reg0 <= 36'sb110000110010111110000000011000010101;
            sine_reg0   <= 36'sb11100001010000101100000101110100111;
        end
        5388: begin
            cosine_reg0 <= 36'sb110000110010010001110001111101101001;
            sine_reg0   <= 36'sb11100001001101101100111110000000111;
        end
        5389: begin
            cosine_reg0 <= 36'sb110000110001100101100100001000011111;
            sine_reg0   <= 36'sb11100001001010101101101101100001010;
        end
        5390: begin
            cosine_reg0 <= 36'sb110000110000111001010110111000111001;
            sine_reg0   <= 36'sb11100001000111101110010100010110000;
        end
        5391: begin
            cosine_reg0 <= 36'sb110000110000001101001010001110111001;
            sine_reg0   <= 36'sb11100001000100101110110010011111010;
        end
        5392: begin
            cosine_reg0 <= 36'sb110000101111100000111110001010100001;
            sine_reg0   <= 36'sb11100001000001101111000111111101001;
        end
        5393: begin
            cosine_reg0 <= 36'sb110000101110110100110010101011110011;
            sine_reg0   <= 36'sb11100000111110101111010100101111111;
        end
        5394: begin
            cosine_reg0 <= 36'sb110000101110001000100111110010101111;
            sine_reg0   <= 36'sb11100000111011101111011000110111100;
        end
        5395: begin
            cosine_reg0 <= 36'sb110000101101011100011101011111011001;
            sine_reg0   <= 36'sb11100000111000101111010100010100001;
        end
        5396: begin
            cosine_reg0 <= 36'sb110000101100110000010011110001110000;
            sine_reg0   <= 36'sb11100000110101101111000111000101110;
        end
        5397: begin
            cosine_reg0 <= 36'sb110000101100000100001010101001111000;
            sine_reg0   <= 36'sb11100000110010101110110001001100110;
        end
        5398: begin
            cosine_reg0 <= 36'sb110000101011011000000010000111110010;
            sine_reg0   <= 36'sb11100000101111101110010010101001000;
        end
        5399: begin
            cosine_reg0 <= 36'sb110000101010101011111010001011011111;
            sine_reg0   <= 36'sb11100000101100101101101011011010110;
        end
        5400: begin
            cosine_reg0 <= 36'sb110000101001111111110010110101000010;
            sine_reg0   <= 36'sb11100000101001101100111011100010001;
        end
        5401: begin
            cosine_reg0 <= 36'sb110000101001010011101100000100011100;
            sine_reg0   <= 36'sb11100000100110101100000010111111001;
        end
        5402: begin
            cosine_reg0 <= 36'sb110000101000100111100101111001101110;
            sine_reg0   <= 36'sb11100000100011101011000001110010000;
        end
        5403: begin
            cosine_reg0 <= 36'sb110000100111111011100000010100111011;
            sine_reg0   <= 36'sb11100000100000101001110111111010110;
        end
        5404: begin
            cosine_reg0 <= 36'sb110000100111001111011011010110000100;
            sine_reg0   <= 36'sb11100000011101101000100101011001100;
        end
        5405: begin
            cosine_reg0 <= 36'sb110000100110100011010110111101001011;
            sine_reg0   <= 36'sb11100000011010100111001010001110100;
        end
        5406: begin
            cosine_reg0 <= 36'sb110000100101110111010011001010010001;
            sine_reg0   <= 36'sb11100000010111100101100110011001110;
        end
        5407: begin
            cosine_reg0 <= 36'sb110000100101001011001111111101011000;
            sine_reg0   <= 36'sb11100000010100100011111001111011011;
        end
        5408: begin
            cosine_reg0 <= 36'sb110000100100011111001101010110100011;
            sine_reg0   <= 36'sb11100000010001100010000100110011100;
        end
        5409: begin
            cosine_reg0 <= 36'sb110000100011110011001011010101110001;
            sine_reg0   <= 36'sb11100000001110100000000111000010010;
        end
        5410: begin
            cosine_reg0 <= 36'sb110000100011000111001001111011000111;
            sine_reg0   <= 36'sb11100000001011011110000000100111110;
        end
        5411: begin
            cosine_reg0 <= 36'sb110000100010011011001001000110100100;
            sine_reg0   <= 36'sb11100000001000011011110001100100001;
        end
        5412: begin
            cosine_reg0 <= 36'sb110000100001101111001000111000001011;
            sine_reg0   <= 36'sb11100000000101011001011001110111100;
        end
        5413: begin
            cosine_reg0 <= 36'sb110000100001000011001001001111111101;
            sine_reg0   <= 36'sb11100000000010010110111001100001111;
        end
        5414: begin
            cosine_reg0 <= 36'sb110000100000010111001010001101111100;
            sine_reg0   <= 36'sb11011111111111010100010000100011100;
        end
        5415: begin
            cosine_reg0 <= 36'sb110000011111101011001011110010001010;
            sine_reg0   <= 36'sb11011111111100010001011110111100100;
        end
        5416: begin
            cosine_reg0 <= 36'sb110000011110111111001101111100101000;
            sine_reg0   <= 36'sb11011111111001001110100100101101000;
        end
        5417: begin
            cosine_reg0 <= 36'sb110000011110010011010000101101011001;
            sine_reg0   <= 36'sb11011111110110001011100001110100111;
        end
        5418: begin
            cosine_reg0 <= 36'sb110000011101100111010100000100011110;
            sine_reg0   <= 36'sb11011111110011001000010110010100101;
        end
        5419: begin
            cosine_reg0 <= 36'sb110000011100111011011000000001111000;
            sine_reg0   <= 36'sb11011111110000000101000010001100001;
        end
        5420: begin
            cosine_reg0 <= 36'sb110000011100001111011100100101101001;
            sine_reg0   <= 36'sb11011111101101000001100101011011100;
        end
        5421: begin
            cosine_reg0 <= 36'sb110000011011100011100001101111110011;
            sine_reg0   <= 36'sb11011111101001111110000000000010111;
        end
        5422: begin
            cosine_reg0 <= 36'sb110000011010110111100111100000011000;
            sine_reg0   <= 36'sb11011111100110111010010010000010011;
        end
        5423: begin
            cosine_reg0 <= 36'sb110000011010001011101101110111011001;
            sine_reg0   <= 36'sb11011111100011110110011011011010010;
        end
        5424: begin
            cosine_reg0 <= 36'sb110000011001011111110100110100111001;
            sine_reg0   <= 36'sb11011111100000110010011100001010100;
        end
        5425: begin
            cosine_reg0 <= 36'sb110000011000110011111100011000110111;
            sine_reg0   <= 36'sb11011111011101101110010100010011010;
        end
        5426: begin
            cosine_reg0 <= 36'sb110000011000001000000100100011011000;
            sine_reg0   <= 36'sb11011111011010101010000011110100101;
        end
        5427: begin
            cosine_reg0 <= 36'sb110000010111011100001101010100011011;
            sine_reg0   <= 36'sb11011111010111100101101010101110101;
        end
        5428: begin
            cosine_reg0 <= 36'sb110000010110110000010110101100000011;
            sine_reg0   <= 36'sb11011111010100100001001001000001101;
        end
        5429: begin
            cosine_reg0 <= 36'sb110000010110000100100000101010010010;
            sine_reg0   <= 36'sb11011111010001011100011110101101101;
        end
        5430: begin
            cosine_reg0 <= 36'sb110000010101011000101011001111001001;
            sine_reg0   <= 36'sb11011111001110010111101011110010101;
        end
        5431: begin
            cosine_reg0 <= 36'sb110000010100101100110110011010101001;
            sine_reg0   <= 36'sb11011111001011010010110000010000111;
        end
        5432: begin
            cosine_reg0 <= 36'sb110000010100000001000010001100110110;
            sine_reg0   <= 36'sb11011111001000001101101100001000011;
        end
        5433: begin
            cosine_reg0 <= 36'sb110000010011010101001110100101101111;
            sine_reg0   <= 36'sb11011111000101001000011111011001100;
        end
        5434: begin
            cosine_reg0 <= 36'sb110000010010101001011011100101010111;
            sine_reg0   <= 36'sb11011111000010000011001010000100001;
        end
        5435: begin
            cosine_reg0 <= 36'sb110000010001111101101001001011110000;
            sine_reg0   <= 36'sb11011110111110111101101100001000011;
        end
        5436: begin
            cosine_reg0 <= 36'sb110000010001010001110111011000111100;
            sine_reg0   <= 36'sb11011110111011111000000101100110100;
        end
        5437: begin
            cosine_reg0 <= 36'sb110000010000100110000110001100111011;
            sine_reg0   <= 36'sb11011110111000110010010110011110100;
        end
        5438: begin
            cosine_reg0 <= 36'sb110000001111111010010101100111110000;
            sine_reg0   <= 36'sb11011110110101101100011110110000101;
        end
        5439: begin
            cosine_reg0 <= 36'sb110000001111001110100101101001011100;
            sine_reg0   <= 36'sb11011110110010100110011110011100111;
        end
        5440: begin
            cosine_reg0 <= 36'sb110000001110100010110110010010000001;
            sine_reg0   <= 36'sb11011110101111100000010101100011011;
        end
        5441: begin
            cosine_reg0 <= 36'sb110000001101110111000111100001100001;
            sine_reg0   <= 36'sb11011110101100011010000100000100011;
        end
        5442: begin
            cosine_reg0 <= 36'sb110000001101001011011001010111111110;
            sine_reg0   <= 36'sb11011110101001010011101001111111110;
        end
        5443: begin
            cosine_reg0 <= 36'sb110000001100011111101011110101011001;
            sine_reg0   <= 36'sb11011110100110001101000111010101111;
        end
        5444: begin
            cosine_reg0 <= 36'sb110000001011110011111110111001110011;
            sine_reg0   <= 36'sb11011110100011000110011100000110110;
        end
        5445: begin
            cosine_reg0 <= 36'sb110000001011001000010010100101001111;
            sine_reg0   <= 36'sb11011110011111111111101000010010100;
        end
        5446: begin
            cosine_reg0 <= 36'sb110000001010011100100110110111101110;
            sine_reg0   <= 36'sb11011110011100111000101011111001010;
        end
        5447: begin
            cosine_reg0 <= 36'sb110000001001110000111011110001010010;
            sine_reg0   <= 36'sb11011110011001110001100110111011001;
        end
        5448: begin
            cosine_reg0 <= 36'sb110000001001000101010001010001111100;
            sine_reg0   <= 36'sb11011110010110101010011001011000010;
        end
        5449: begin
            cosine_reg0 <= 36'sb110000001000011001100111011001101110;
            sine_reg0   <= 36'sb11011110010011100011000011010000110;
        end
        5450: begin
            cosine_reg0 <= 36'sb110000000111101101111110001000101011;
            sine_reg0   <= 36'sb11011110010000011011100100100100110;
        end
        5451: begin
            cosine_reg0 <= 36'sb110000000111000010010101011110110011;
            sine_reg0   <= 36'sb11011110001101010011111101010100011;
        end
        5452: begin
            cosine_reg0 <= 36'sb110000000110010110101101011100001000;
            sine_reg0   <= 36'sb11011110001010001100001101011111101;
        end
        5453: begin
            cosine_reg0 <= 36'sb110000000101101011000110000000101100;
            sine_reg0   <= 36'sb11011110000111000100010101000110110;
        end
        5454: begin
            cosine_reg0 <= 36'sb110000000100111111011111001100100001;
            sine_reg0   <= 36'sb11011110000011111100010100001001111;
        end
        5455: begin
            cosine_reg0 <= 36'sb110000000100010011111000111111101000;
            sine_reg0   <= 36'sb11011110000000110100001010101001001;
        end
        5456: begin
            cosine_reg0 <= 36'sb110000000011101000010011011010000100;
            sine_reg0   <= 36'sb11011101111101101011111000100100100;
        end
        5457: begin
            cosine_reg0 <= 36'sb110000000010111100101110011011110100;
            sine_reg0   <= 36'sb11011101111010100011011101111100010;
        end
        5458: begin
            cosine_reg0 <= 36'sb110000000010010001001010000100111101;
            sine_reg0   <= 36'sb11011101110111011010111010110000011;
        end
        5459: begin
            cosine_reg0 <= 36'sb110000000001100101100110010101011110;
            sine_reg0   <= 36'sb11011101110100010010001111000001001;
        end
        5460: begin
            cosine_reg0 <= 36'sb110000000000111010000011001101011010;
            sine_reg0   <= 36'sb11011101110001001001011010101110101;
        end
        5461: begin
            cosine_reg0 <= 36'sb110000000000001110100000101100110010;
            sine_reg0   <= 36'sb11011101101110000000011101111000111;
        end
        5462: begin
            cosine_reg0 <= 36'sb101111111111100010111110110011101000;
            sine_reg0   <= 36'sb11011101101010110111011000100000000;
        end
        5463: begin
            cosine_reg0 <= 36'sb101111111110110111011101100001111110;
            sine_reg0   <= 36'sb11011101100111101110001010100100010;
        end
        5464: begin
            cosine_reg0 <= 36'sb101111111110001011111100110111110110;
            sine_reg0   <= 36'sb11011101100100100100110100000101101;
        end
        5465: begin
            cosine_reg0 <= 36'sb101111111101100000011100110101010000;
            sine_reg0   <= 36'sb11011101100001011011010101000100010;
        end
        5466: begin
            cosine_reg0 <= 36'sb101111111100110100111101011010001111;
            sine_reg0   <= 36'sb11011101011110010001101101100000011;
        end
        5467: begin
            cosine_reg0 <= 36'sb101111111100001001011110100110110101;
            sine_reg0   <= 36'sb11011101011011000111111101011010000;
        end
        5468: begin
            cosine_reg0 <= 36'sb101111111011011110000000011011000011;
            sine_reg0   <= 36'sb11011101010111111110000100110001011;
        end
        5469: begin
            cosine_reg0 <= 36'sb101111111010110010100010110110111011;
            sine_reg0   <= 36'sb11011101010100110100000011100110011;
        end
        5470: begin
            cosine_reg0 <= 36'sb101111111010000111000101111010011110;
            sine_reg0   <= 36'sb11011101010001101001111001111001011;
        end
        5471: begin
            cosine_reg0 <= 36'sb101111111001011011101001100101101110;
            sine_reg0   <= 36'sb11011101001110011111100111101010011;
        end
        5472: begin
            cosine_reg0 <= 36'sb101111111000110000001101111000101101;
            sine_reg0   <= 36'sb11011101001011010101001100111001101;
        end
        5473: begin
            cosine_reg0 <= 36'sb101111111000000100110010110011011101;
            sine_reg0   <= 36'sb11011101001000001010101001100111000;
        end
        5474: begin
            cosine_reg0 <= 36'sb101111110111011001011000010101111111;
            sine_reg0   <= 36'sb11011101000100111111111101110010110;
        end
        5475: begin
            cosine_reg0 <= 36'sb101111110110101101111110100000010101;
            sine_reg0   <= 36'sb11011101000001110101001001011101001;
        end
        5476: begin
            cosine_reg0 <= 36'sb101111110110000010100101010010100000;
            sine_reg0   <= 36'sb11011100111110101010001100100110001;
        end
        5477: begin
            cosine_reg0 <= 36'sb101111110101010111001100101100100010;
            sine_reg0   <= 36'sb11011100111011011111000111001101110;
        end
        5478: begin
            cosine_reg0 <= 36'sb101111110100101011110100101110011101;
            sine_reg0   <= 36'sb11011100111000010011111001010100011;
        end
        5479: begin
            cosine_reg0 <= 36'sb101111110100000000011101011000010011;
            sine_reg0   <= 36'sb11011100110101001000100010111010000;
        end
        5480: begin
            cosine_reg0 <= 36'sb101111110011010101000110101010000101;
            sine_reg0   <= 36'sb11011100110001111101000011111110101;
        end
        5481: begin
            cosine_reg0 <= 36'sb101111110010101001110000100011110101;
            sine_reg0   <= 36'sb11011100101110110001011100100010101;
        end
        5482: begin
            cosine_reg0 <= 36'sb101111110001111110011011000101100100;
            sine_reg0   <= 36'sb11011100101011100101101100100110000;
        end
        5483: begin
            cosine_reg0 <= 36'sb101111110001010011000110001111010101;
            sine_reg0   <= 36'sb11011100101000011001110100001000110;
        end
        5484: begin
            cosine_reg0 <= 36'sb101111110000100111110010000001001001;
            sine_reg0   <= 36'sb11011100100101001101110011001011010;
        end
        5485: begin
            cosine_reg0 <= 36'sb101111101111111100011110011011000001;
            sine_reg0   <= 36'sb11011100100010000001101001101101011;
        end
        5486: begin
            cosine_reg0 <= 36'sb101111101111010001001011011100111111;
            sine_reg0   <= 36'sb11011100011110110101010111101111011;
        end
        5487: begin
            cosine_reg0 <= 36'sb101111101110100101111001000111000101;
            sine_reg0   <= 36'sb11011100011011101000111101010001011;
        end
        5488: begin
            cosine_reg0 <= 36'sb101111101101111010100111011001010101;
            sine_reg0   <= 36'sb11011100011000011100011010010011100;
        end
        5489: begin
            cosine_reg0 <= 36'sb101111101101001111010110010011110000;
            sine_reg0   <= 36'sb11011100010101001111101110110101111;
        end
        5490: begin
            cosine_reg0 <= 36'sb101111101100100100000101110110011000;
            sine_reg0   <= 36'sb11011100010010000010111010111000101;
        end
        5491: begin
            cosine_reg0 <= 36'sb101111101011111000110110000001001110;
            sine_reg0   <= 36'sb11011100001110110101111110011011110;
        end
        5492: begin
            cosine_reg0 <= 36'sb101111101011001101100110110100010101;
            sine_reg0   <= 36'sb11011100001011101000111001011111100;
        end
        5493: begin
            cosine_reg0 <= 36'sb101111101010100010011000001111101110;
            sine_reg0   <= 36'sb11011100001000011011101100000100000;
        end
        5494: begin
            cosine_reg0 <= 36'sb101111101001110111001010010011011010;
            sine_reg0   <= 36'sb11011100000101001110010110001001011;
        end
        5495: begin
            cosine_reg0 <= 36'sb101111101001001011111100111111011100;
            sine_reg0   <= 36'sb11011100000010000000110111101111110;
        end
        5496: begin
            cosine_reg0 <= 36'sb101111101000100000110000010011110100;
            sine_reg0   <= 36'sb11011011111110110011010000110111001;
        end
        5497: begin
            cosine_reg0 <= 36'sb101111100111110101100100010000100101;
            sine_reg0   <= 36'sb11011011111011100101100001011111110;
        end
        5498: begin
            cosine_reg0 <= 36'sb101111100111001010011000110101110000;
            sine_reg0   <= 36'sb11011011111000010111101001101001110;
        end
        5499: begin
            cosine_reg0 <= 36'sb101111100110011111001110000011010111;
            sine_reg0   <= 36'sb11011011110101001001101001010101001;
        end
        5500: begin
            cosine_reg0 <= 36'sb101111100101110100000011111001011100;
            sine_reg0   <= 36'sb11011011110001111011100000100010010;
        end
        5501: begin
            cosine_reg0 <= 36'sb101111100101001000111010011000000000;
            sine_reg0   <= 36'sb11011011101110101101001111010000111;
        end
        5502: begin
            cosine_reg0 <= 36'sb101111100100011101110001011111000101;
            sine_reg0   <= 36'sb11011011101011011110110101100001100;
        end
        5503: begin
            cosine_reg0 <= 36'sb101111100011110010101001001110101100;
            sine_reg0   <= 36'sb11011011101000010000010011010100000;
        end
        5504: begin
            cosine_reg0 <= 36'sb101111100011000111100001100110111000;
            sine_reg0   <= 36'sb11011011100101000001101000101000101;
        end
        5505: begin
            cosine_reg0 <= 36'sb101111100010011100011010100111101001;
            sine_reg0   <= 36'sb11011011100001110010110101011111100;
        end
        5506: begin
            cosine_reg0 <= 36'sb101111100001110001010100010001000010;
            sine_reg0   <= 36'sb11011011011110100011111001111000110;
        end
        5507: begin
            cosine_reg0 <= 36'sb101111100001000110001110100011000100;
            sine_reg0   <= 36'sb11011011011011010100110101110100011;
        end
        5508: begin
            cosine_reg0 <= 36'sb101111100000011011001001011101110010;
            sine_reg0   <= 36'sb11011011011000000101101001010010101;
        end
        5509: begin
            cosine_reg0 <= 36'sb101111011111110000000101000001001011;
            sine_reg0   <= 36'sb11011011010100110110010100010011100;
        end
        5510: begin
            cosine_reg0 <= 36'sb101111011111000101000001001101010011;
            sine_reg0   <= 36'sb11011011010001100110110110110111010;
        end
        5511: begin
            cosine_reg0 <= 36'sb101111011110011001111110000010001011;
            sine_reg0   <= 36'sb11011011001110010111010000111110000;
        end
        5512: begin
            cosine_reg0 <= 36'sb101111011101101110111011011111110100;
            sine_reg0   <= 36'sb11011011001011000111100010100111111;
        end
        5513: begin
            cosine_reg0 <= 36'sb101111011101000011111001100110010000;
            sine_reg0   <= 36'sb11011011000111110111101011110100111;
        end
        5514: begin
            cosine_reg0 <= 36'sb101111011100011000111000010101100001;
            sine_reg0   <= 36'sb11011011000100100111101100100101010;
        end
        5515: begin
            cosine_reg0 <= 36'sb101111011011101101110111101101101001;
            sine_reg0   <= 36'sb11011011000001010111100100111001000;
        end
        5516: begin
            cosine_reg0 <= 36'sb101111011011000010110111101110101001;
            sine_reg0   <= 36'sb11011010111110000111010100110000100;
        end
        5517: begin
            cosine_reg0 <= 36'sb101111011010010111111000011000100010;
            sine_reg0   <= 36'sb11011010111010110110111100001011101;
        end
        5518: begin
            cosine_reg0 <= 36'sb101111011001101100111001101011010111;
            sine_reg0   <= 36'sb11011010110111100110011011001010100;
        end
        5519: begin
            cosine_reg0 <= 36'sb101111011001000001111011100111001010;
            sine_reg0   <= 36'sb11011010110100010101110001101101100;
        end
        5520: begin
            cosine_reg0 <= 36'sb101111011000010110111110001011111011;
            sine_reg0   <= 36'sb11011010110001000100111111110100100;
        end
        5521: begin
            cosine_reg0 <= 36'sb101111010111101100000001011001101100;
            sine_reg0   <= 36'sb11011010101101110100000101011111101;
        end
        5522: begin
            cosine_reg0 <= 36'sb101111010111000001000101010000011111;
            sine_reg0   <= 36'sb11011010101010100011000010101111010;
        end
        5523: begin
            cosine_reg0 <= 36'sb101111010110010110001001110000010111;
            sine_reg0   <= 36'sb11011010100111010001110111100011010;
        end
        5524: begin
            cosine_reg0 <= 36'sb101111010101101011001110111001010011;
            sine_reg0   <= 36'sb11011010100100000000100011111011111;
        end
        5525: begin
            cosine_reg0 <= 36'sb101111010101000000010100101011010111;
            sine_reg0   <= 36'sb11011010100000101111000111111001010;
        end
        5526: begin
            cosine_reg0 <= 36'sb101111010100010101011011000110100011;
            sine_reg0   <= 36'sb11011010011101011101100011011011011;
        end
        5527: begin
            cosine_reg0 <= 36'sb101111010011101010100010001010111010;
            sine_reg0   <= 36'sb11011010011010001011110110100010101;
        end
        5528: begin
            cosine_reg0 <= 36'sb101111010010111111101001111000011101;
            sine_reg0   <= 36'sb11011010010110111010000001001110111;
        end
        5529: begin
            cosine_reg0 <= 36'sb101111010010010100110010001111001101;
            sine_reg0   <= 36'sb11011010010011101000000011100000011;
        end
        5530: begin
            cosine_reg0 <= 36'sb101111010001101001111011001111001101;
            sine_reg0   <= 36'sb11011010010000010101111101010111001;
        end
        5531: begin
            cosine_reg0 <= 36'sb101111010000111111000100111000011101;
            sine_reg0   <= 36'sb11011010001101000011101110110011100;
        end
        5532: begin
            cosine_reg0 <= 36'sb101111010000010100001111001011000001;
            sine_reg0   <= 36'sb11011010001001110001010111110101011;
        end
        5533: begin
            cosine_reg0 <= 36'sb101111001111101001011010000110111000;
            sine_reg0   <= 36'sb11011010000110011110111000011101000;
        end
        5534: begin
            cosine_reg0 <= 36'sb101111001110111110100101101100000110;
            sine_reg0   <= 36'sb11011010000011001100010000101010100;
        end
        5535: begin
            cosine_reg0 <= 36'sb101111001110010011110001111010101011;
            sine_reg0   <= 36'sb11011001111111111001100000011110000;
        end
        5536: begin
            cosine_reg0 <= 36'sb101111001101101000111110110010101001;
            sine_reg0   <= 36'sb11011001111100100110100111110111100;
        end
        5537: begin
            cosine_reg0 <= 36'sb101111001100111110001100010100000010;
            sine_reg0   <= 36'sb11011001111001010011100110110111011;
        end
        5538: begin
            cosine_reg0 <= 36'sb101111001100010011011010011110111000;
            sine_reg0   <= 36'sb11011001110110000000011101011101101;
        end
        5539: begin
            cosine_reg0 <= 36'sb101111001011101000101001010011001100;
            sine_reg0   <= 36'sb11011001110010101101001011101010010;
        end
        5540: begin
            cosine_reg0 <= 36'sb101111001010111101111000110001000000;
            sine_reg0   <= 36'sb11011001101111011001110001011101100;
        end
        5541: begin
            cosine_reg0 <= 36'sb101111001010010011001000111000010101;
            sine_reg0   <= 36'sb11011001101100000110001110110111101;
        end
        5542: begin
            cosine_reg0 <= 36'sb101111001001101000011001101001001101;
            sine_reg0   <= 36'sb11011001101000110010100011111000100;
        end
        5543: begin
            cosine_reg0 <= 36'sb101111001000111101101011000011101010;
            sine_reg0   <= 36'sb11011001100101011110110000100000100;
        end
        5544: begin
            cosine_reg0 <= 36'sb101111001000010010111101000111101110;
            sine_reg0   <= 36'sb11011001100010001010110100101111100;
        end
        5545: begin
            cosine_reg0 <= 36'sb101111000111101000001111110101011001;
            sine_reg0   <= 36'sb11011001011110110110110000100101110;
        end
        5546: begin
            cosine_reg0 <= 36'sb101111000110111101100011001100101110;
            sine_reg0   <= 36'sb11011001011011100010100100000011100;
        end
        5547: begin
            cosine_reg0 <= 36'sb101111000110010010110111001101101111;
            sine_reg0   <= 36'sb11011001011000001110001111001000110;
        end
        5548: begin
            cosine_reg0 <= 36'sb101111000101101000001011111000011101;
            sine_reg0   <= 36'sb11011001010100111001110001110101100;
        end
        5549: begin
            cosine_reg0 <= 36'sb101111000100111101100001001100111001;
            sine_reg0   <= 36'sb11011001010001100101001100001010001;
        end
        5550: begin
            cosine_reg0 <= 36'sb101111000100010010110111001011000101;
            sine_reg0   <= 36'sb11011001001110010000011110000110101;
        end
        5551: begin
            cosine_reg0 <= 36'sb101111000011101000001101110011000100;
            sine_reg0   <= 36'sb11011001001010111011100111101011010;
        end
        5552: begin
            cosine_reg0 <= 36'sb101111000010111101100101000100110110;
            sine_reg0   <= 36'sb11011001000111100110101000110111111;
        end
        5553: begin
            cosine_reg0 <= 36'sb101111000010010010111101000000011101;
            sine_reg0   <= 36'sb11011001000100010001100001101100111;
        end
        5554: begin
            cosine_reg0 <= 36'sb101111000001101000010101100101111011;
            sine_reg0   <= 36'sb11011001000000111100010010001010010;
        end
        5555: begin
            cosine_reg0 <= 36'sb101111000000111101101110110101010010;
            sine_reg0   <= 36'sb11011000111101100110111010010000001;
        end
        5556: begin
            cosine_reg0 <= 36'sb101111000000010011001000101110100011;
            sine_reg0   <= 36'sb11011000111010010001011001111110110;
        end
        5557: begin
            cosine_reg0 <= 36'sb101110111111101000100011010001101111;
            sine_reg0   <= 36'sb11011000110110111011110001010110001;
        end
        5558: begin
            cosine_reg0 <= 36'sb101110111110111101111110011110111001;
            sine_reg0   <= 36'sb11011000110011100110000000010110011;
        end
        5559: begin
            cosine_reg0 <= 36'sb101110111110010011011010010110000011;
            sine_reg0   <= 36'sb11011000110000010000000110111111110;
        end
        5560: begin
            cosine_reg0 <= 36'sb101110111101101000110110110111001100;
            sine_reg0   <= 36'sb11011000101100111010000101010010010;
        end
        5561: begin
            cosine_reg0 <= 36'sb101110111100111110010100000010011001;
            sine_reg0   <= 36'sb11011000101001100011111011001110001;
        end
        5562: begin
            cosine_reg0 <= 36'sb101110111100010011110001110111101001;
            sine_reg0   <= 36'sb11011000100110001101101000110011011;
        end
        5563: begin
            cosine_reg0 <= 36'sb101110111011101001010000010110111111;
            sine_reg0   <= 36'sb11011000100010110111001110000010010;
        end
        5564: begin
            cosine_reg0 <= 36'sb101110111010111110101111100000011100;
            sine_reg0   <= 36'sb11011000011111100000101010111010110;
        end
        5565: begin
            cosine_reg0 <= 36'sb101110111010010100001111010100000010;
            sine_reg0   <= 36'sb11011000011100001001111111011101001;
        end
        5566: begin
            cosine_reg0 <= 36'sb101110111001101001101111110001110010;
            sine_reg0   <= 36'sb11011000011000110011001011101001100;
        end
        5567: begin
            cosine_reg0 <= 36'sb101110111000111111010000111001101111;
            sine_reg0   <= 36'sb11011000010101011100001111011111111;
        end
        5568: begin
            cosine_reg0 <= 36'sb101110111000010100110010101011111010;
            sine_reg0   <= 36'sb11011000010010000101001011000000100;
        end
        5569: begin
            cosine_reg0 <= 36'sb101110110111101010010101001000010100;
            sine_reg0   <= 36'sb11011000001110101101111110001011100;
        end
        5570: begin
            cosine_reg0 <= 36'sb101110110110111111111000001110111111;
            sine_reg0   <= 36'sb11011000001011010110101001000001000;
        end
        5571: begin
            cosine_reg0 <= 36'sb101110110110010101011011111111111101;
            sine_reg0   <= 36'sb11011000000111111111001011100001000;
        end
        5572: begin
            cosine_reg0 <= 36'sb101110110101101011000000011011001111;
            sine_reg0   <= 36'sb11011000000100100111100101101011110;
        end
        5573: begin
            cosine_reg0 <= 36'sb101110110101000000100101100000111000;
            sine_reg0   <= 36'sb11011000000001001111110111100001100;
        end
        5574: begin
            cosine_reg0 <= 36'sb101110110100010110001011010000111000;
            sine_reg0   <= 36'sb11010111111101111000000001000010001;
        end
        5575: begin
            cosine_reg0 <= 36'sb101110110011101011110001101011010001;
            sine_reg0   <= 36'sb11010111111010100000000010001101111;
        end
        5576: begin
            cosine_reg0 <= 36'sb101110110011000001011000110000000101;
            sine_reg0   <= 36'sb11010111110111000111111011000100111;
        end
        5577: begin
            cosine_reg0 <= 36'sb101110110010010111000000011111010110;
            sine_reg0   <= 36'sb11010111110011101111101011100111010;
        end
        5578: begin
            cosine_reg0 <= 36'sb101110110001101100101000111001000101;
            sine_reg0   <= 36'sb11010111110000010111010011110101010;
        end
        5579: begin
            cosine_reg0 <= 36'sb101110110001000010010001111101010011;
            sine_reg0   <= 36'sb11010111101100111110110011101110110;
        end
        5580: begin
            cosine_reg0 <= 36'sb101110110000010111111011101100000100;
            sine_reg0   <= 36'sb11010111101001100110001011010100001;
        end
        5581: begin
            cosine_reg0 <= 36'sb101110101111101101100110000101010111;
            sine_reg0   <= 36'sb11010111100110001101011010100101011;
        end
        5582: begin
            cosine_reg0 <= 36'sb101110101111000011010001001001001111;
            sine_reg0   <= 36'sb11010111100010110100100001100010101;
        end
        5583: begin
            cosine_reg0 <= 36'sb101110101110011000111100110111101101;
            sine_reg0   <= 36'sb11010111011111011011100000001100000;
        end
        5584: begin
            cosine_reg0 <= 36'sb101110101101101110101001010000110100;
            sine_reg0   <= 36'sb11010111011100000010010110100001110;
        end
        5585: begin
            cosine_reg0 <= 36'sb101110101101000100010110010100100100;
            sine_reg0   <= 36'sb11010111011000101001000100100100000;
        end
        5586: begin
            cosine_reg0 <= 36'sb101110101100011010000100000010111111;
            sine_reg0   <= 36'sb11010111010101001111101010010010101;
        end
        5587: begin
            cosine_reg0 <= 36'sb101110101011101111110010011100000111;
            sine_reg0   <= 36'sb11010111010001110110000111101110001;
        end
        5588: begin
            cosine_reg0 <= 36'sb101110101011000101100001011111111110;
            sine_reg0   <= 36'sb11010111001110011100011100110110010;
        end
        5589: begin
            cosine_reg0 <= 36'sb101110101010011011010001001110100100;
            sine_reg0   <= 36'sb11010111001011000010101001101011100;
        end
        5590: begin
            cosine_reg0 <= 36'sb101110101001110001000001100111111101;
            sine_reg0   <= 36'sb11010111000111101000101110001101110;
        end
        5591: begin
            cosine_reg0 <= 36'sb101110101001000110110010101100001001;
            sine_reg0   <= 36'sb11010111000100001110101010011101010;
        end
        5592: begin
            cosine_reg0 <= 36'sb101110101000011100100100011011001010;
            sine_reg0   <= 36'sb11010111000000110100011110011010001;
        end
        5593: begin
            cosine_reg0 <= 36'sb101110100111110010010110110101000001;
            sine_reg0   <= 36'sb11010110111101011010001010000100011;
        end
        5594: begin
            cosine_reg0 <= 36'sb101110100111001000001001111001110001;
            sine_reg0   <= 36'sb11010110111001111111101101011100010;
        end
        5595: begin
            cosine_reg0 <= 36'sb101110100110011101111101101001011011;
            sine_reg0   <= 36'sb11010110110110100101001000100010000;
        end
        5596: begin
            cosine_reg0 <= 36'sb101110100101110011110010000100000000;
            sine_reg0   <= 36'sb11010110110011001010011011010101100;
        end
        5597: begin
            cosine_reg0 <= 36'sb101110100101001001100111001001100010;
            sine_reg0   <= 36'sb11010110101111101111100101110111000;
        end
        5598: begin
            cosine_reg0 <= 36'sb101110100100011111011100111010000100;
            sine_reg0   <= 36'sb11010110101100010100101000000110101;
        end
        5599: begin
            cosine_reg0 <= 36'sb101110100011110101010011010101100101;
            sine_reg0   <= 36'sb11010110101000111001100010000100101;
        end
        5600: begin
            cosine_reg0 <= 36'sb101110100011001011001010011100001001;
            sine_reg0   <= 36'sb11010110100101011110010011110001000;
        end
        5601: begin
            cosine_reg0 <= 36'sb101110100010100001000010001101110000;
            sine_reg0   <= 36'sb11010110100010000010111101001011111;
        end
        5602: begin
            cosine_reg0 <= 36'sb101110100001110110111010101010011101;
            sine_reg0   <= 36'sb11010110011110100111011110010101011;
        end
        5603: begin
            cosine_reg0 <= 36'sb101110100001001100110011110010010000;
            sine_reg0   <= 36'sb11010110011011001011110111001101101;
        end
        5604: begin
            cosine_reg0 <= 36'sb101110100000100010101101100101001100;
            sine_reg0   <= 36'sb11010110010111110000000111110100111;
        end
        5605: begin
            cosine_reg0 <= 36'sb101110011111111000101000000011010010;
            sine_reg0   <= 36'sb11010110010100010100010000001011010;
        end
        5606: begin
            cosine_reg0 <= 36'sb101110011111001110100011001100100100;
            sine_reg0   <= 36'sb11010110010000111000010000010000110;
        end
        5607: begin
            cosine_reg0 <= 36'sb101110011110100100011111000001000100;
            sine_reg0   <= 36'sb11010110001101011100001000000101101;
        end
        5608: begin
            cosine_reg0 <= 36'sb101110011101111010011011100000110010;
            sine_reg0   <= 36'sb11010110001001111111110111101001111;
        end
        5609: begin
            cosine_reg0 <= 36'sb101110011101010000011000101011110001;
            sine_reg0   <= 36'sb11010110000110100011011110111101110;
        end
        5610: begin
            cosine_reg0 <= 36'sb101110011100100110010110100010000010;
            sine_reg0   <= 36'sb11010110000011000110111110000001011;
        end
        5611: begin
            cosine_reg0 <= 36'sb101110011011111100010101000011100111;
            sine_reg0   <= 36'sb11010101111111101010010100110100110;
        end
        5612: begin
            cosine_reg0 <= 36'sb101110011011010010010100010000100010;
            sine_reg0   <= 36'sb11010101111100001101100011011000010;
        end
        5613: begin
            cosine_reg0 <= 36'sb101110011010101000010100001000110100;
            sine_reg0   <= 36'sb11010101111000110000101001101011111;
        end
        5614: begin
            cosine_reg0 <= 36'sb101110011001111110010100101100011110;
            sine_reg0   <= 36'sb11010101110101010011100111101111101;
        end
        5615: begin
            cosine_reg0 <= 36'sb101110011001010100010101111011100011;
            sine_reg0   <= 36'sb11010101110001110110011101100011111;
        end
        5616: begin
            cosine_reg0 <= 36'sb101110011000101010010111110110000100;
            sine_reg0   <= 36'sb11010101101110011001001011001000101;
        end
        5617: begin
            cosine_reg0 <= 36'sb101110011000000000011010011100000010;
            sine_reg0   <= 36'sb11010101101010111011110000011110000;
        end
        5618: begin
            cosine_reg0 <= 36'sb101110010111010110011101101101100000;
            sine_reg0   <= 36'sb11010101100111011110001101100100001;
        end
        5619: begin
            cosine_reg0 <= 36'sb101110010110101100100001101010011110;
            sine_reg0   <= 36'sb11010101100100000000100010011011010;
        end
        5620: begin
            cosine_reg0 <= 36'sb101110010110000010100110010010111111;
            sine_reg0   <= 36'sb11010101100000100010101111000011100;
        end
        5621: begin
            cosine_reg0 <= 36'sb101110010101011000101011100111000100;
            sine_reg0   <= 36'sb11010101011101000100110011011100110;
        end
        5622: begin
            cosine_reg0 <= 36'sb101110010100101110110001100110101111;
            sine_reg0   <= 36'sb11010101011001100110101111100111100;
        end
        5623: begin
            cosine_reg0 <= 36'sb101110010100000100111000010010000001;
            sine_reg0   <= 36'sb11010101010110001000100011100011101;
        end
        5624: begin
            cosine_reg0 <= 36'sb101110010011011010111111101000111100;
            sine_reg0   <= 36'sb11010101010010101010001111010001010;
        end
        5625: begin
            cosine_reg0 <= 36'sb101110010010110001000111101011100001;
            sine_reg0   <= 36'sb11010101001111001011110010110000110;
        end
        5626: begin
            cosine_reg0 <= 36'sb101110010010000111010000011001110011;
            sine_reg0   <= 36'sb11010101001011101101001110000010000;
        end
        5627: begin
            cosine_reg0 <= 36'sb101110010001011101011001110011110010;
            sine_reg0   <= 36'sb11010101001000001110100001000101011;
        end
        5628: begin
            cosine_reg0 <= 36'sb101110010000110011100011111001100000;
            sine_reg0   <= 36'sb11010101000100101111101011111010110;
        end
        5629: begin
            cosine_reg0 <= 36'sb101110010000001001101110101011000000;
            sine_reg0   <= 36'sb11010101000001010000101110100010011;
        end
        5630: begin
            cosine_reg0 <= 36'sb101110001111011111111010001000010010;
            sine_reg0   <= 36'sb11010100111101110001101000111100100;
        end
        5631: begin
            cosine_reg0 <= 36'sb101110001110110110000110010001011001;
            sine_reg0   <= 36'sb11010100111010010010011011001001001;
        end
        5632: begin
            cosine_reg0 <= 36'sb101110001110001100010011000110010101;
            sine_reg0   <= 36'sb11010100110110110011000101001000011;
        end
        5633: begin
            cosine_reg0 <= 36'sb101110001101100010100000100111001001;
            sine_reg0   <= 36'sb11010100110011010011100110111010011;
        end
        5634: begin
            cosine_reg0 <= 36'sb101110001100111000101110110011110101;
            sine_reg0   <= 36'sb11010100101111110100000000011111011;
        end
        5635: begin
            cosine_reg0 <= 36'sb101110001100001110111101101100011101;
            sine_reg0   <= 36'sb11010100101100010100010001110111100;
        end
        5636: begin
            cosine_reg0 <= 36'sb101110001011100101001101010001000000;
            sine_reg0   <= 36'sb11010100101000110100011011000010110;
        end
        5637: begin
            cosine_reg0 <= 36'sb101110001010111011011101100001100010;
            sine_reg0   <= 36'sb11010100100101010100011100000001011;
        end
        5638: begin
            cosine_reg0 <= 36'sb101110001010010001101110011110000011;
            sine_reg0   <= 36'sb11010100100001110100010100110011011;
        end
        5639: begin
            cosine_reg0 <= 36'sb101110001001101000000000000110100101;
            sine_reg0   <= 36'sb11010100011110010100000101011001001;
        end
        5640: begin
            cosine_reg0 <= 36'sb101110001000111110010010011011001001;
            sine_reg0   <= 36'sb11010100011010110011101101110010100;
        end
        5641: begin
            cosine_reg0 <= 36'sb101110001000010100100101011011110011;
            sine_reg0   <= 36'sb11010100010111010011001101111111111;
        end
        5642: begin
            cosine_reg0 <= 36'sb101110000111101010111001001000100001;
            sine_reg0   <= 36'sb11010100010011110010100110000001001;
        end
        5643: begin
            cosine_reg0 <= 36'sb101110000111000001001101100001011000;
            sine_reg0   <= 36'sb11010100010000010001110101110110101;
        end
        5644: begin
            cosine_reg0 <= 36'sb101110000110010111100010100110011000;
            sine_reg0   <= 36'sb11010100001100110000111101100000011;
        end
        5645: begin
            cosine_reg0 <= 36'sb101110000101101101111000010111100010;
            sine_reg0   <= 36'sb11010100001001001111111100111110100;
        end
        5646: begin
            cosine_reg0 <= 36'sb101110000101000100001110110100111001;
            sine_reg0   <= 36'sb11010100000101101110110100010001010;
        end
        5647: begin
            cosine_reg0 <= 36'sb101110000100011010100101111110011101;
            sine_reg0   <= 36'sb11010100000010001101100011011000101;
        end
        5648: begin
            cosine_reg0 <= 36'sb101110000011110000111101110100010001;
            sine_reg0   <= 36'sb11010011111110101100001010010100111;
        end
        5649: begin
            cosine_reg0 <= 36'sb101110000011000111010110010110010111;
            sine_reg0   <= 36'sb11010011111011001010101001000110001;
        end
        5650: begin
            cosine_reg0 <= 36'sb101110000010011101101111100100101111;
            sine_reg0   <= 36'sb11010011110111101000111111101100011;
        end
        5651: begin
            cosine_reg0 <= 36'sb101110000001110100001001011111011011;
            sine_reg0   <= 36'sb11010011110100000111001110000111111;
        end
        5652: begin
            cosine_reg0 <= 36'sb101110000001001010100100000110011110;
            sine_reg0   <= 36'sb11010011110000100101010100011000110;
        end
        5653: begin
            cosine_reg0 <= 36'sb101110000000100000111111011001111000;
            sine_reg0   <= 36'sb11010011101101000011010010011111010;
        end
        5654: begin
            cosine_reg0 <= 36'sb101101111111110111011011011001101011;
            sine_reg0   <= 36'sb11010011101001100001001000011011010;
        end
        5655: begin
            cosine_reg0 <= 36'sb101101111111001101111000000101111001;
            sine_reg0   <= 36'sb11010011100101111110110110001101001;
        end
        5656: begin
            cosine_reg0 <= 36'sb101101111110100100010101011110100011;
            sine_reg0   <= 36'sb11010011100010011100011011110100111;
        end
        5657: begin
            cosine_reg0 <= 36'sb101101111101111010110011100011101100;
            sine_reg0   <= 36'sb11010011011110111001111001010010101;
        end
        5658: begin
            cosine_reg0 <= 36'sb101101111101010001010010010101010011;
            sine_reg0   <= 36'sb11010011011011010111001110100110101;
        end
        5659: begin
            cosine_reg0 <= 36'sb101101111100100111110001110011011100;
            sine_reg0   <= 36'sb11010011010111110100011011110000111;
        end
        5660: begin
            cosine_reg0 <= 36'sb101101111011111110010001111110001000;
            sine_reg0   <= 36'sb11010011010100010001100000110001101;
        end
        5661: begin
            cosine_reg0 <= 36'sb101101111011010100110010110101011001;
            sine_reg0   <= 36'sb11010011010000101110011101101001000;
        end
        5662: begin
            cosine_reg0 <= 36'sb101101111010101011010100011001001111;
            sine_reg0   <= 36'sb11010011001101001011010010010111001;
        end
        5663: begin
            cosine_reg0 <= 36'sb101101111010000001110110101001101101;
            sine_reg0   <= 36'sb11010011001001100111111110111100000;
        end
        5664: begin
            cosine_reg0 <= 36'sb101101111001011000011001100110110100;
            sine_reg0   <= 36'sb11010011000110000100100011011000000;
        end
        5665: begin
            cosine_reg0 <= 36'sb101101111000101110111101010000100101;
            sine_reg0   <= 36'sb11010011000010100000111111101011001;
        end
        5666: begin
            cosine_reg0 <= 36'sb101101111000000101100001100111000011;
            sine_reg0   <= 36'sb11010010111110111101010011110101100;
        end
        5667: begin
            cosine_reg0 <= 36'sb101101110111011100000110101010010000;
            sine_reg0   <= 36'sb11010010111011011001011111110111010;
        end
        5668: begin
            cosine_reg0 <= 36'sb101101110110110010101100011010001011;
            sine_reg0   <= 36'sb11010010110111110101100011110000101;
        end
        5669: begin
            cosine_reg0 <= 36'sb101101110110001001010010110110111000;
            sine_reg0   <= 36'sb11010010110100010001011111100001110;
        end
        5670: begin
            cosine_reg0 <= 36'sb101101110101011111111010000000011000;
            sine_reg0   <= 36'sb11010010110000101101010011001010101;
        end
        5671: begin
            cosine_reg0 <= 36'sb101101110100110110100001110110101100;
            sine_reg0   <= 36'sb11010010101101001000111110101011100;
        end
        5672: begin
            cosine_reg0 <= 36'sb101101110100001101001010011001110110;
            sine_reg0   <= 36'sb11010010101001100100100010000100011;
        end
        5673: begin
            cosine_reg0 <= 36'sb101101110011100011110011101001110111;
            sine_reg0   <= 36'sb11010010100101111111111101010101101;
        end
        5674: begin
            cosine_reg0 <= 36'sb101101110010111010011101100110110010;
            sine_reg0   <= 36'sb11010010100010011011010000011111010;
        end
        5675: begin
            cosine_reg0 <= 36'sb101101110010010001001000010000100111;
            sine_reg0   <= 36'sb11010010011110110110011011100001011;
        end
        5676: begin
            cosine_reg0 <= 36'sb101101110001100111110011100111011001;
            sine_reg0   <= 36'sb11010010011011010001011110011100001;
        end
        5677: begin
            cosine_reg0 <= 36'sb101101110000111110011111101011001000;
            sine_reg0   <= 36'sb11010010010111101100011001001111101;
        end
        5678: begin
            cosine_reg0 <= 36'sb101101110000010101001100011011110111;
            sine_reg0   <= 36'sb11010010010100000111001011111100001;
        end
        5679: begin
            cosine_reg0 <= 36'sb101101101111101011111001111001100111;
            sine_reg0   <= 36'sb11010010010000100001110110100001101;
        end
        5680: begin
            cosine_reg0 <= 36'sb101101101111000010101000000100011010;
            sine_reg0   <= 36'sb11010010001100111100011001000000100;
        end
        5681: begin
            cosine_reg0 <= 36'sb101101101110011001010110111100010010;
            sine_reg0   <= 36'sb11010010001001010110110011011000100;
        end
        5682: begin
            cosine_reg0 <= 36'sb101101101101110000000110100001001111;
            sine_reg0   <= 36'sb11010010000101110001000101101010001;
        end
        5683: begin
            cosine_reg0 <= 36'sb101101101101000110110110110011010011;
            sine_reg0   <= 36'sb11010010000010001011001111110101011;
        end
        5684: begin
            cosine_reg0 <= 36'sb101101101100011101100111110010100001;
            sine_reg0   <= 36'sb11010001111110100101010001111010011;
        end
        5685: begin
            cosine_reg0 <= 36'sb101101101011110100011001011110111001;
            sine_reg0   <= 36'sb11010001111010111111001011111001010;
        end
        5686: begin
            cosine_reg0 <= 36'sb101101101011001011001011111000011110;
            sine_reg0   <= 36'sb11010001110111011000111101110010001;
        end
        5687: begin
            cosine_reg0 <= 36'sb101101101010100001111110111111010000;
            sine_reg0   <= 36'sb11010001110011110010100111100101010;
        end
        5688: begin
            cosine_reg0 <= 36'sb101101101001111000110010110011010010;
            sine_reg0   <= 36'sb11010001110000001100001001010010101;
        end
        5689: begin
            cosine_reg0 <= 36'sb101101101001001111100111010100100100;
            sine_reg0   <= 36'sb11010001101100100101100010111010100;
        end
        5690: begin
            cosine_reg0 <= 36'sb101101101000100110011100100011001010;
            sine_reg0   <= 36'sb11010001101000111110110100011101000;
        end
        5691: begin
            cosine_reg0 <= 36'sb101101100111111101010010011111000011;
            sine_reg0   <= 36'sb11010001100101010111111101111010010;
        end
        5692: begin
            cosine_reg0 <= 36'sb101101100111010100001001001000010011;
            sine_reg0   <= 36'sb11010001100001110000111111010010010;
        end
        5693: begin
            cosine_reg0 <= 36'sb101101100110101011000000011110111001;
            sine_reg0   <= 36'sb11010001011110001001111000100101011;
        end
        5694: begin
            cosine_reg0 <= 36'sb101101100110000001111000100010111001;
            sine_reg0   <= 36'sb11010001011010100010101001110011101;
        end
        5695: begin
            cosine_reg0 <= 36'sb101101100101011000110001010100010011;
            sine_reg0   <= 36'sb11010001010110111011010010111101001;
        end
        5696: begin
            cosine_reg0 <= 36'sb101101100100101111101010110011001001;
            sine_reg0   <= 36'sb11010001010011010011110100000010001;
        end
        5697: begin
            cosine_reg0 <= 36'sb101101100100000110100100111111011101;
            sine_reg0   <= 36'sb11010001001111101100001101000010101;
        end
        5698: begin
            cosine_reg0 <= 36'sb101101100011011101011111111001010000;
            sine_reg0   <= 36'sb11010001001100000100011101111110111;
        end
        5699: begin
            cosine_reg0 <= 36'sb101101100010110100011011100000100101;
            sine_reg0   <= 36'sb11010001001000011100100110110110111;
        end
        5700: begin
            cosine_reg0 <= 36'sb101101100010001011010111110101011011;
            sine_reg0   <= 36'sb11010001000100110100100111101011000;
        end
        5701: begin
            cosine_reg0 <= 36'sb101101100001100010010100110111110110;
            sine_reg0   <= 36'sb11010001000001001100100000011011001;
        end
        5702: begin
            cosine_reg0 <= 36'sb101101100000111001010010100111110110;
            sine_reg0   <= 36'sb11010000111101100100010001000111101;
        end
        5703: begin
            cosine_reg0 <= 36'sb101101100000010000010001000101011101;
            sine_reg0   <= 36'sb11010000111001111011111001110000100;
        end
        5704: begin
            cosine_reg0 <= 36'sb101101011111100111010000010000101101;
            sine_reg0   <= 36'sb11010000110110010011011010010101111;
        end
        5705: begin
            cosine_reg0 <= 36'sb101101011110111110010000001001101000;
            sine_reg0   <= 36'sb11010000110010101010110010111000000;
        end
        5706: begin
            cosine_reg0 <= 36'sb101101011110010101010000110000001110;
            sine_reg0   <= 36'sb11010000101111000010000011010111000;
        end
        5707: begin
            cosine_reg0 <= 36'sb101101011101101100010010000100100010;
            sine_reg0   <= 36'sb11010000101011011001001011110010111;
        end
        5708: begin
            cosine_reg0 <= 36'sb101101011101000011010100000110100101;
            sine_reg0   <= 36'sb11010000100111110000001100001011111;
        end
        5709: begin
            cosine_reg0 <= 36'sb101101011100011010010110110110011001;
            sine_reg0   <= 36'sb11010000100100000111000100100010001;
        end
        5710: begin
            cosine_reg0 <= 36'sb101101011011110001011010010011111111;
            sine_reg0   <= 36'sb11010000100000011101110100110101110;
        end
        5711: begin
            cosine_reg0 <= 36'sb101101011011001000011110011111011001;
            sine_reg0   <= 36'sb11010000011100110100011101000110111;
        end
        5712: begin
            cosine_reg0 <= 36'sb101101011010011111100011011000101000;
            sine_reg0   <= 36'sb11010000011001001010111101010101110;
        end
        5713: begin
            cosine_reg0 <= 36'sb101101011001110110101000111111101110;
            sine_reg0   <= 36'sb11010000010101100001010101100010011;
        end
        5714: begin
            cosine_reg0 <= 36'sb101101011001001101101111010100101101;
            sine_reg0   <= 36'sb11010000010001110111100101101101000;
        end
        5715: begin
            cosine_reg0 <= 36'sb101101011000100100110110010111100110;
            sine_reg0   <= 36'sb11010000001110001101101101110101101;
        end
        5716: begin
            cosine_reg0 <= 36'sb101101010111111011111110001000011011;
            sine_reg0   <= 36'sb11010000001010100011101101111100101;
        end
        5717: begin
            cosine_reg0 <= 36'sb101101010111010011000110100111001100;
            sine_reg0   <= 36'sb11010000000110111001100110000001111;
        end
        5718: begin
            cosine_reg0 <= 36'sb101101010110101010001111110011111101;
            sine_reg0   <= 36'sb11010000000011001111010110000101110;
        end
        5719: begin
            cosine_reg0 <= 36'sb101101010110000001011001101110101111;
            sine_reg0   <= 36'sb11001111111111100100111110001000001;
        end
        5720: begin
            cosine_reg0 <= 36'sb101101010101011000100100010111100010;
            sine_reg0   <= 36'sb11001111111011111010011110001001100;
        end
        5721: begin
            cosine_reg0 <= 36'sb101101010100101111101111101110011001;
            sine_reg0   <= 36'sb11001111111000001111110110001001101;
        end
        5722: begin
            cosine_reg0 <= 36'sb101101010100000110111011110011010101;
            sine_reg0   <= 36'sb11001111110100100101000110001000111;
        end
        5723: begin
            cosine_reg0 <= 36'sb101101010011011110001000100110011000;
            sine_reg0   <= 36'sb11001111110000111010001110000111011;
        end
        5724: begin
            cosine_reg0 <= 36'sb101101010010110101010110000111100011;
            sine_reg0   <= 36'sb11001111101101001111001110000101010;
        end
        5725: begin
            cosine_reg0 <= 36'sb101101010010001100100100010110111000;
            sine_reg0   <= 36'sb11001111101001100100000110000010101;
        end
        5726: begin
            cosine_reg0 <= 36'sb101101010001100011110011010100011000;
            sine_reg0   <= 36'sb11001111100101111000110101111111101;
        end
        5727: begin
            cosine_reg0 <= 36'sb101101010000111011000011000000000110;
            sine_reg0   <= 36'sb11001111100010001101011101111100100;
        end
        5728: begin
            cosine_reg0 <= 36'sb101101010000010010010011011010000010;
            sine_reg0   <= 36'sb11001111011110100001111101111001010;
        end
        5729: begin
            cosine_reg0 <= 36'sb101101001111101001100100100010001110;
            sine_reg0   <= 36'sb11001111011010110110010101110110000;
        end
        5730: begin
            cosine_reg0 <= 36'sb101101001111000000110110011000101100;
            sine_reg0   <= 36'sb11001111010111001010100101110011000;
        end
        5731: begin
            cosine_reg0 <= 36'sb101101001110011000001000111101011110;
            sine_reg0   <= 36'sb11001111010011011110101101110000011;
        end
        5732: begin
            cosine_reg0 <= 36'sb101101001101101111011100010000100100;
            sine_reg0   <= 36'sb11001111001111110010101101101110010;
        end
        5733: begin
            cosine_reg0 <= 36'sb101101001101000110110000010010000000;
            sine_reg0   <= 36'sb11001111001100000110100101101100110;
        end
        5734: begin
            cosine_reg0 <= 36'sb101101001100011110000101000001110101;
            sine_reg0   <= 36'sb11001111001000011010010101101100000;
        end
        5735: begin
            cosine_reg0 <= 36'sb101101001011110101011010100000000011;
            sine_reg0   <= 36'sb11001111000100101101111101101100010;
        end
        5736: begin
            cosine_reg0 <= 36'sb101101001011001100110000101100101101;
            sine_reg0   <= 36'sb11001111000001000001011101101101100;
        end
        5737: begin
            cosine_reg0 <= 36'sb101101001010100100000111100111110011;
            sine_reg0   <= 36'sb11001110111101010100110101110000000;
        end
        5738: begin
            cosine_reg0 <= 36'sb101101001001111011011111010001011000;
            sine_reg0   <= 36'sb11001110111001101000000101110011111;
        end
        5739: begin
            cosine_reg0 <= 36'sb101101001001010010110111101001011100;
            sine_reg0   <= 36'sb11001110110101111011001101111001001;
        end
        5740: begin
            cosine_reg0 <= 36'sb101101001000101010010000110000000010;
            sine_reg0   <= 36'sb11001110110010001110001110000000001;
        end
        5741: begin
            cosine_reg0 <= 36'sb101101001000000001101010100101001010;
            sine_reg0   <= 36'sb11001110101110100001000110001000111;
        end
        5742: begin
            cosine_reg0 <= 36'sb101101000111011001000101001000111000;
            sine_reg0   <= 36'sb11001110101010110011110110010011100;
        end
        5743: begin
            cosine_reg0 <= 36'sb101101000110110000100000011011001011;
            sine_reg0   <= 36'sb11001110100111000110011110100000010;
        end
        5744: begin
            cosine_reg0 <= 36'sb101101000110000111111100011100000110;
            sine_reg0   <= 36'sb11001110100011011000111110101111010;
        end
        5745: begin
            cosine_reg0 <= 36'sb101101000101011111011001001011101011;
            sine_reg0   <= 36'sb11001110011111101011010111000000100;
        end
        5746: begin
            cosine_reg0 <= 36'sb101101000100110110110110101001111010;
            sine_reg0   <= 36'sb11001110011011111101100111010100010;
        end
        5747: begin
            cosine_reg0 <= 36'sb101101000100001110010100110110110101;
            sine_reg0   <= 36'sb11001110011000001111101111101010110;
        end
        5748: begin
            cosine_reg0 <= 36'sb101101000011100101110011110010011111;
            sine_reg0   <= 36'sb11001110010100100001110000000011111;
        end
        5749: begin
            cosine_reg0 <= 36'sb101101000010111101010011011100111000;
            sine_reg0   <= 36'sb11001110010000110011101000100000000;
        end
        5750: begin
            cosine_reg0 <= 36'sb101101000010010100110011110110000010;
            sine_reg0   <= 36'sb11001110001101000101011000111111010;
        end
        5751: begin
            cosine_reg0 <= 36'sb101101000001101100010100111101111111;
            sine_reg0   <= 36'sb11001110001001010111000001100001101;
        end
        5752: begin
            cosine_reg0 <= 36'sb101101000001000011110110110100110000;
            sine_reg0   <= 36'sb11001110000101101000100010000111011;
        end
        5753: begin
            cosine_reg0 <= 36'sb101101000000011011011001011010010110;
            sine_reg0   <= 36'sb11001110000001111001111010110000101;
        end
        5754: begin
            cosine_reg0 <= 36'sb101100111111110010111100101110110100;
            sine_reg0   <= 36'sb11001101111110001011001011011101101;
        end
        5755: begin
            cosine_reg0 <= 36'sb101100111111001010100000110010001011;
            sine_reg0   <= 36'sb11001101111010011100010100001110010;
        end
        5756: begin
            cosine_reg0 <= 36'sb101100111110100010000101100100011100;
            sine_reg0   <= 36'sb11001101110110101101010101000010111;
        end
        5757: begin
            cosine_reg0 <= 36'sb101100111101111001101011000101101001;
            sine_reg0   <= 36'sb11001101110010111110001101111011100;
        end
        5758: begin
            cosine_reg0 <= 36'sb101100111101010001010001010101110100;
            sine_reg0   <= 36'sb11001101101111001110111110111000100;
        end
        5759: begin
            cosine_reg0 <= 36'sb101100111100101000111000010100111110;
            sine_reg0   <= 36'sb11001101101011011111100111111001110;
        end
        5760: begin
            cosine_reg0 <= 36'sb101100111100000000100000000011001000;
            sine_reg0   <= 36'sb11001101100111110000001000111111100;
        end
        5761: begin
            cosine_reg0 <= 36'sb101100111011011000001000100000010101;
            sine_reg0   <= 36'sb11001101100100000000100010001001111;
        end
        5762: begin
            cosine_reg0 <= 36'sb101100111010101111110001101100100101;
            sine_reg0   <= 36'sb11001101100000010000110011011001001;
        end
        5763: begin
            cosine_reg0 <= 36'sb101100111010000111011011100111111011;
            sine_reg0   <= 36'sb11001101011100100000111100101101010;
        end
        5764: begin
            cosine_reg0 <= 36'sb101100111001011111000110010010011000;
            sine_reg0   <= 36'sb11001101011000110000111110000110100;
        end
        5765: begin
            cosine_reg0 <= 36'sb101100111000110110110001101011111101;
            sine_reg0   <= 36'sb11001101010101000000110111100101000;
        end
        5766: begin
            cosine_reg0 <= 36'sb101100111000001110011101110100101100;
            sine_reg0   <= 36'sb11001101010001010000101001001000111;
        end
        5767: begin
            cosine_reg0 <= 36'sb101100110111100110001010101100100110;
            sine_reg0   <= 36'sb11001101001101100000010010110010010;
        end
        5768: begin
            cosine_reg0 <= 36'sb101100110110111101111000010011101110;
            sine_reg0   <= 36'sb11001101001001101111110100100001010;
        end
        5769: begin
            cosine_reg0 <= 36'sb101100110110010101100110101010000101;
            sine_reg0   <= 36'sb11001101000101111111001110010110001;
        end
        5770: begin
            cosine_reg0 <= 36'sb101100110101101101010101101111101011;
            sine_reg0   <= 36'sb11001101000010001110100000010000111;
        end
        5771: begin
            cosine_reg0 <= 36'sb101100110101000101000101100100100011;
            sine_reg0   <= 36'sb11001100111110011101101010010001110;
        end
        5772: begin
            cosine_reg0 <= 36'sb101100110100011100110110001000101111;
            sine_reg0   <= 36'sb11001100111010101100101100011000111;
        end
        5773: begin
            cosine_reg0 <= 36'sb101100110011110100100111011100001111;
            sine_reg0   <= 36'sb11001100110110111011100110100110011;
        end
        5774: begin
            cosine_reg0 <= 36'sb101100110011001100011001011111000110;
            sine_reg0   <= 36'sb11001100110011001010011000111010011;
        end
        5775: begin
            cosine_reg0 <= 36'sb101100110010100100001100010001010101;
            sine_reg0   <= 36'sb11001100101111011001000011010101001;
        end
        5776: begin
            cosine_reg0 <= 36'sb101100110001111011111111110010111101;
            sine_reg0   <= 36'sb11001100101011100111100101110110101;
        end
        5777: begin
            cosine_reg0 <= 36'sb101100110001010011110100000100000001;
            sine_reg0   <= 36'sb11001100100111110110000000011111001;
        end
        5778: begin
            cosine_reg0 <= 36'sb101100110000101011101001000100100001;
            sine_reg0   <= 36'sb11001100100100000100010011001110110;
        end
        5779: begin
            cosine_reg0 <= 36'sb101100110000000011011110110100011111;
            sine_reg0   <= 36'sb11001100100000010010011110000101101;
        end
        5780: begin
            cosine_reg0 <= 36'sb101100101111011011010101010011111101;
            sine_reg0   <= 36'sb11001100011100100000100001000100000;
        end
        5781: begin
            cosine_reg0 <= 36'sb101100101110110011001100100010111100;
            sine_reg0   <= 36'sb11001100011000101110011100001001110;
        end
        5782: begin
            cosine_reg0 <= 36'sb101100101110001011000100100001011110;
            sine_reg0   <= 36'sb11001100010100111100001111010111011;
        end
        5783: begin
            cosine_reg0 <= 36'sb101100101101100010111101001111100100;
            sine_reg0   <= 36'sb11001100010001001001111010101100110;
        end
        5784: begin
            cosine_reg0 <= 36'sb101100101100111010110110101101010000;
            sine_reg0   <= 36'sb11001100001101010111011110001010001;
        end
        5785: begin
            cosine_reg0 <= 36'sb101100101100010010110000111010100100;
            sine_reg0   <= 36'sb11001100001001100100111001101111101;
        end
        5786: begin
            cosine_reg0 <= 36'sb101100101011101010101011110111100000;
            sine_reg0   <= 36'sb11001100000101110010001101011101011;
        end
        5787: begin
            cosine_reg0 <= 36'sb101100101011000010100111100100001000;
            sine_reg0   <= 36'sb11001100000001111111011001010011101;
        end
        5788: begin
            cosine_reg0 <= 36'sb101100101010011010100100000000011011;
            sine_reg0   <= 36'sb11001011111110001100011101010010011;
        end
        5789: begin
            cosine_reg0 <= 36'sb101100101001110010100001001100011011;
            sine_reg0   <= 36'sb11001011111010011001011001011001111;
        end
        5790: begin
            cosine_reg0 <= 36'sb101100101001001010011111001000001011;
            sine_reg0   <= 36'sb11001011110110100110001101101010010;
        end
        5791: begin
            cosine_reg0 <= 36'sb101100101000100010011101110011101100;
            sine_reg0   <= 36'sb11001011110010110010111010000011101;
        end
        5792: begin
            cosine_reg0 <= 36'sb101100100111111010011101001110111111;
            sine_reg0   <= 36'sb11001011101110111111011110100110001;
        end
        5793: begin
            cosine_reg0 <= 36'sb101100100111010010011101011010000110;
            sine_reg0   <= 36'sb11001011101011001011111011010010000;
        end
        5794: begin
            cosine_reg0 <= 36'sb101100100110101010011110010101000010;
            sine_reg0   <= 36'sb11001011100111011000010000000111010;
        end
        5795: begin
            cosine_reg0 <= 36'sb101100100110000010011111111111110101;
            sine_reg0   <= 36'sb11001011100011100100011101000110010;
        end
        5796: begin
            cosine_reg0 <= 36'sb101100100101011010100010011010100000;
            sine_reg0   <= 36'sb11001011011111110000100010001110111;
        end
        5797: begin
            cosine_reg0 <= 36'sb101100100100110010100101100101000101;
            sine_reg0   <= 36'sb11001011011011111100011111100001011;
        end
        5798: begin
            cosine_reg0 <= 36'sb101100100100001010101001011111100110;
            sine_reg0   <= 36'sb11001011011000001000010100111110000;
        end
        5799: begin
            cosine_reg0 <= 36'sb101100100011100010101110001010000100;
            sine_reg0   <= 36'sb11001011010100010100000010100100110;
        end
        5800: begin
            cosine_reg0 <= 36'sb101100100010111010110011100100100000;
            sine_reg0   <= 36'sb11001011010000011111101000010101111;
        end
        5801: begin
            cosine_reg0 <= 36'sb101100100010010010111001101110111101;
            sine_reg0   <= 36'sb11001011001100101011000110010001011;
        end
        5802: begin
            cosine_reg0 <= 36'sb101100100001101011000000101001011011;
            sine_reg0   <= 36'sb11001011001000110110011100010111101;
        end
        5803: begin
            cosine_reg0 <= 36'sb101100100001000011001000010011111100;
            sine_reg0   <= 36'sb11001011000101000001101010101000101;
        end
        5804: begin
            cosine_reg0 <= 36'sb101100100000011011010000101110100010;
            sine_reg0   <= 36'sb11001011000001001100110001000100100;
        end
        5805: begin
            cosine_reg0 <= 36'sb101100011111110011011001111001001111;
            sine_reg0   <= 36'sb11001010111101010111101111101011100;
        end
        5806: begin
            cosine_reg0 <= 36'sb101100011111001011100011110100000011;
            sine_reg0   <= 36'sb11001010111001100010100110011101110;
        end
        5807: begin
            cosine_reg0 <= 36'sb101100011110100011101110011111000000;
            sine_reg0   <= 36'sb11001010110101101101010101011011010;
        end
        5808: begin
            cosine_reg0 <= 36'sb101100011101111011111001111010001001;
            sine_reg0   <= 36'sb11001010110001110111111100100100011;
        end
        5809: begin
            cosine_reg0 <= 36'sb101100011101010100000110000101011101;
            sine_reg0   <= 36'sb11001010101110000010011011111001001;
        end
        5810: begin
            cosine_reg0 <= 36'sb101100011100101100010011000001000000;
            sine_reg0   <= 36'sb11001010101010001100110011011001101;
        end
        5811: begin
            cosine_reg0 <= 36'sb101100011100000100100000101100110010;
            sine_reg0   <= 36'sb11001010100110010111000011000110001;
        end
        5812: begin
            cosine_reg0 <= 36'sb101100011011011100101111001000110101;
            sine_reg0   <= 36'sb11001010100010100001001010111110110;
        end
        5813: begin
            cosine_reg0 <= 36'sb101100011010110100111110010101001011;
            sine_reg0   <= 36'sb11001010011110101011001011000011101;
        end
        5814: begin
            cosine_reg0 <= 36'sb101100011010001101001110010001110101;
            sine_reg0   <= 36'sb11001010011010110101000011010100111;
        end
        5815: begin
            cosine_reg0 <= 36'sb101100011001100101011110111110110100;
            sine_reg0   <= 36'sb11001010010110111110110011110010110;
        end
        5816: begin
            cosine_reg0 <= 36'sb101100011000111101110000011100001011;
            sine_reg0   <= 36'sb11001010010011001000011100011101010;
        end
        5817: begin
            cosine_reg0 <= 36'sb101100011000010110000010101001111010;
            sine_reg0   <= 36'sb11001010001111010001111101010100101;
        end
        5818: begin
            cosine_reg0 <= 36'sb101100010111101110010101101000000100;
            sine_reg0   <= 36'sb11001010001011011011010110011001000;
        end
        5819: begin
            cosine_reg0 <= 36'sb101100010111000110101001010110101001;
            sine_reg0   <= 36'sb11001010000111100100100111101010100;
        end
        5820: begin
            cosine_reg0 <= 36'sb101100010110011110111101110101101011;
            sine_reg0   <= 36'sb11001010000011101101110001001001011;
        end
        5821: begin
            cosine_reg0 <= 36'sb101100010101110111010011000101001101;
            sine_reg0   <= 36'sb11001001111111110110110010110101101;
        end
        5822: begin
            cosine_reg0 <= 36'sb101100010101001111101001000101001110;
            sine_reg0   <= 36'sb11001001111011111111101100101111011;
        end
        5823: begin
            cosine_reg0 <= 36'sb101100010100100111111111110101110010;
            sine_reg0   <= 36'sb11001001111000001000011110110111000;
        end
        5824: begin
            cosine_reg0 <= 36'sb101100010100000000010111010110111001;
            sine_reg0   <= 36'sb11001001110100010001001001001100100;
        end
        5825: begin
            cosine_reg0 <= 36'sb101100010011011000101111101000100100;
            sine_reg0   <= 36'sb11001001110000011001101011110000000;
        end
        5826: begin
            cosine_reg0 <= 36'sb101100010010110001001000101010110110;
            sine_reg0   <= 36'sb11001001101100100010000110100001101;
        end
        5827: begin
            cosine_reg0 <= 36'sb101100010010001001100010011101110001;
            sine_reg0   <= 36'sb11001001101000101010011001100001110;
        end
        5828: begin
            cosine_reg0 <= 36'sb101100010001100001111101000001010100;
            sine_reg0   <= 36'sb11001001100100110010100100110000010;
        end
        5829: begin
            cosine_reg0 <= 36'sb101100010000111010011000010101100011;
            sine_reg0   <= 36'sb11001001100000111010101000001101011;
        end
        5830: begin
            cosine_reg0 <= 36'sb101100010000010010110100011010011110;
            sine_reg0   <= 36'sb11001001011101000010100011111001010;
        end
        5831: begin
            cosine_reg0 <= 36'sb101100001111101011010001010000000111;
            sine_reg0   <= 36'sb11001001011001001010010111110100001;
        end
        5832: begin
            cosine_reg0 <= 36'sb101100001111000011101110110110100000;
            sine_reg0   <= 36'sb11001001010101010010000011111110001;
        end
        5833: begin
            cosine_reg0 <= 36'sb101100001110011100001101001101101010;
            sine_reg0   <= 36'sb11001001010001011001101000010111010;
        end
        5834: begin
            cosine_reg0 <= 36'sb101100001101110100101100010101100111;
            sine_reg0   <= 36'sb11001001001101100001000100111111110;
        end
        5835: begin
            cosine_reg0 <= 36'sb101100001101001101001100001110011000;
            sine_reg0   <= 36'sb11001001001001101000011001110111111;
        end
        5836: begin
            cosine_reg0 <= 36'sb101100001100100101101100110111111110;
            sine_reg0   <= 36'sb11001001000101101111100110111111101;
        end
        5837: begin
            cosine_reg0 <= 36'sb101100001011111110001110010010011100;
            sine_reg0   <= 36'sb11001001000001110110101100010111010;
        end
        5838: begin
            cosine_reg0 <= 36'sb101100001011010110110000011101110010;
            sine_reg0   <= 36'sb11001000111101111101101001111110111;
        end
        5839: begin
            cosine_reg0 <= 36'sb101100001010101111010011011010000011;
            sine_reg0   <= 36'sb11001000111010000100011111110110100;
        end
        5840: begin
            cosine_reg0 <= 36'sb101100001010000111110111000111001111;
            sine_reg0   <= 36'sb11001000110110001011001101111110100;
        end
        5841: begin
            cosine_reg0 <= 36'sb101100001001100000011011100101011001;
            sine_reg0   <= 36'sb11001000110010010001110100010111000;
        end
        5842: begin
            cosine_reg0 <= 36'sb101100001000111001000000110100100010;
            sine_reg0   <= 36'sb11001000101110011000010011000000000;
        end
        5843: begin
            cosine_reg0 <= 36'sb101100001000010001100110110100101010;
            sine_reg0   <= 36'sb11001000101010011110101001111001110;
        end
        5844: begin
            cosine_reg0 <= 36'sb101100000111101010001101100101110101;
            sine_reg0   <= 36'sb11001000100110100100111001000100011;
        end
        5845: begin
            cosine_reg0 <= 36'sb101100000111000010110101001000000011;
            sine_reg0   <= 36'sb11001000100010101011000000100000000;
        end
        5846: begin
            cosine_reg0 <= 36'sb101100000110011011011101011011010110;
            sine_reg0   <= 36'sb11001000011110110001000000001100111;
        end
        5847: begin
            cosine_reg0 <= 36'sb101100000101110100000110011111110000;
            sine_reg0   <= 36'sb11001000011010110110111000001011000;
        end
        5848: begin
            cosine_reg0 <= 36'sb101100000101001100110000010101010001;
            sine_reg0   <= 36'sb11001000010110111100101000011010101;
        end
        5849: begin
            cosine_reg0 <= 36'sb101100000100100101011010111011111100;
            sine_reg0   <= 36'sb11001000010011000010010000111011111;
        end
        5850: begin
            cosine_reg0 <= 36'sb101100000011111110000110010011110010;
            sine_reg0   <= 36'sb11001000001111000111110001101111000;
        end
        5851: begin
            cosine_reg0 <= 36'sb101100000011010110110010011100110100;
            sine_reg0   <= 36'sb11001000001011001101001010110100000;
        end
        5852: begin
            cosine_reg0 <= 36'sb101100000010101111011111010111000100;
            sine_reg0   <= 36'sb11001000000111010010011100001011001;
        end
        5853: begin
            cosine_reg0 <= 36'sb101100000010001000001101000010100100;
            sine_reg0   <= 36'sb11001000000011010111100101110100011;
        end
        5854: begin
            cosine_reg0 <= 36'sb101100000001100000111011011111010101;
            sine_reg0   <= 36'sb11000111111111011100100111110000001;
        end
        5855: begin
            cosine_reg0 <= 36'sb101100000000111001101010101101011000;
            sine_reg0   <= 36'sb11000111111011100001100001111110011;
        end
        5856: begin
            cosine_reg0 <= 36'sb101100000000010010011010101100101111;
            sine_reg0   <= 36'sb11000111110111100110010100011111011;
        end
        5857: begin
            cosine_reg0 <= 36'sb101011111111101011001011011101011100;
            sine_reg0   <= 36'sb11000111110011101010111111010011010;
        end
        5858: begin
            cosine_reg0 <= 36'sb101011111111000011111100111111100000;
            sine_reg0   <= 36'sb11000111101111101111100010011010000;
        end
        5859: begin
            cosine_reg0 <= 36'sb101011111110011100101111010010111101;
            sine_reg0   <= 36'sb11000111101011110011111101110011111;
        end
        5860: begin
            cosine_reg0 <= 36'sb101011111101110101100010010111110011;
            sine_reg0   <= 36'sb11000111100111111000010001100001001;
        end
        5861: begin
            cosine_reg0 <= 36'sb101011111101001110010110001110000110;
            sine_reg0   <= 36'sb11000111100011111100011101100001111;
        end
        5862: begin
            cosine_reg0 <= 36'sb101011111100100111001010110101110101;
            sine_reg0   <= 36'sb11000111100000000000100001110110001;
        end
        5863: begin
            cosine_reg0 <= 36'sb101011111100000000000000001111000011;
            sine_reg0   <= 36'sb11000111011100000100011110011110010;
        end
        5864: begin
            cosine_reg0 <= 36'sb101011111011011000110110011001110001;
            sine_reg0   <= 36'sb11000111011000001000010011011010001;
        end
        5865: begin
            cosine_reg0 <= 36'sb101011111010110001101101010110000001;
            sine_reg0   <= 36'sb11000111010100001100000000101010001;
        end
        5866: begin
            cosine_reg0 <= 36'sb101011111010001010100101000011110100;
            sine_reg0   <= 36'sb11000111010000001111100110001110011;
        end
        5867: begin
            cosine_reg0 <= 36'sb101011111001100011011101100011001100;
            sine_reg0   <= 36'sb11000111001100010011000100000111000;
        end
        5868: begin
            cosine_reg0 <= 36'sb101011111000111100010110110100001010;
            sine_reg0   <= 36'sb11000111001000010110011010010100001;
        end
        5869: begin
            cosine_reg0 <= 36'sb101011111000010101010000110110101111;
            sine_reg0   <= 36'sb11000111000100011001101000110101111;
        end
        5870: begin
            cosine_reg0 <= 36'sb101011110111101110001011101010111110;
            sine_reg0   <= 36'sb11000111000000011100101111101100011;
        end
        5871: begin
            cosine_reg0 <= 36'sb101011110111000111000111010000110111;
            sine_reg0   <= 36'sb11000110111100011111101110111000000;
        end
        5872: begin
            cosine_reg0 <= 36'sb101011110110100000000011101000011101;
            sine_reg0   <= 36'sb11000110111000100010100110011000101;
        end
        5873: begin
            cosine_reg0 <= 36'sb101011110101111001000000110001110000;
            sine_reg0   <= 36'sb11000110110100100101010110001110100;
        end
        5874: begin
            cosine_reg0 <= 36'sb101011110101010001111110101100110011;
            sine_reg0   <= 36'sb11000110110000100111111110011001111;
        end
        5875: begin
            cosine_reg0 <= 36'sb101011110100101010111101011001100110;
            sine_reg0   <= 36'sb11000110101100101010011110111010111;
        end
        5876: begin
            cosine_reg0 <= 36'sb101011110100000011111100111000001100;
            sine_reg0   <= 36'sb11000110101000101100110111110001100;
        end
        5877: begin
            cosine_reg0 <= 36'sb101011110011011100111101001000100101;
            sine_reg0   <= 36'sb11000110100100101111001000111110001;
        end
        5878: begin
            cosine_reg0 <= 36'sb101011110010110101111110001010110011;
            sine_reg0   <= 36'sb11000110100000110001010010100000110;
        end
        5879: begin
            cosine_reg0 <= 36'sb101011110010001110111111111110111001;
            sine_reg0   <= 36'sb11000110011100110011010100011001100;
        end
        5880: begin
            cosine_reg0 <= 36'sb101011110001101000000010100100110110;
            sine_reg0   <= 36'sb11000110011000110101001110101000101;
        end
        5881: begin
            cosine_reg0 <= 36'sb101011110001000001000101111100101101;
            sine_reg0   <= 36'sb11000110010100110111000001001110010;
        end
        5882: begin
            cosine_reg0 <= 36'sb101011110000011010001010000110100000;
            sine_reg0   <= 36'sb11000110010000111000101100001010101;
        end
        5883: begin
            cosine_reg0 <= 36'sb101011101111110011001111000010001111;
            sine_reg0   <= 36'sb11000110001100111010001111011101101;
        end
        5884: begin
            cosine_reg0 <= 36'sb101011101111001100010100101111111100;
            sine_reg0   <= 36'sb11000110001000111011101011000111110;
        end
        5885: begin
            cosine_reg0 <= 36'sb101011101110100101011011001111101001;
            sine_reg0   <= 36'sb11000110000100111100111111001000111;
        end
        5886: begin
            cosine_reg0 <= 36'sb101011101101111110100010100001011000;
            sine_reg0   <= 36'sb11000110000000111110001011100001010;
        end
        5887: begin
            cosine_reg0 <= 36'sb101011101101010111101010100101001001;
            sine_reg0   <= 36'sb11000101111100111111010000010001001;
        end
        5888: begin
            cosine_reg0 <= 36'sb101011101100110000110011011010111110;
            sine_reg0   <= 36'sb11000101111001000000001101011000100;
        end
        5889: begin
            cosine_reg0 <= 36'sb101011101100001001111101000010111001;
            sine_reg0   <= 36'sb11000101110101000001000010110111110;
        end
        5890: begin
            cosine_reg0 <= 36'sb101011101011100011000111011100111100;
            sine_reg0   <= 36'sb11000101110001000001110000101110110;
        end
        5891: begin
            cosine_reg0 <= 36'sb101011101010111100010010101001000111;
            sine_reg0   <= 36'sb11000101101101000010010110111101110;
        end
        5892: begin
            cosine_reg0 <= 36'sb101011101010010101011110100111011100;
            sine_reg0   <= 36'sb11000101101001000010110101100101000;
        end
        5893: begin
            cosine_reg0 <= 36'sb101011101001101110101011010111111101;
            sine_reg0   <= 36'sb11000101100101000011001100100100100;
        end
        5894: begin
            cosine_reg0 <= 36'sb101011101001000111111000111010101100;
            sine_reg0   <= 36'sb11000101100001000011011011111100101;
        end
        5895: begin
            cosine_reg0 <= 36'sb101011101000100001000111001111101001;
            sine_reg0   <= 36'sb11000101011101000011100011101101011;
        end
        5896: begin
            cosine_reg0 <= 36'sb101011100111111010010110010110110110;
            sine_reg0   <= 36'sb11000101011001000011100011110110111;
        end
        5897: begin
            cosine_reg0 <= 36'sb101011100111010011100110010000010101;
            sine_reg0   <= 36'sb11000101010101000011011100011001011;
        end
        5898: begin
            cosine_reg0 <= 36'sb101011100110101100110110111100000111;
            sine_reg0   <= 36'sb11000101010001000011001101010100111;
        end
        5899: begin
            cosine_reg0 <= 36'sb101011100110000110001000011010001110;
            sine_reg0   <= 36'sb11000101001101000010110110101001110;
        end
        5900: begin
            cosine_reg0 <= 36'sb101011100101011111011010101010101011;
            sine_reg0   <= 36'sb11000101001001000010011000011000000;
        end
        5901: begin
            cosine_reg0 <= 36'sb101011100100111000101101101101011111;
            sine_reg0   <= 36'sb11000101000101000001110010011111111;
        end
        5902: begin
            cosine_reg0 <= 36'sb101011100100010010000001100010101101;
            sine_reg0   <= 36'sb11000101000001000001000101000001011;
        end
        5903: begin
            cosine_reg0 <= 36'sb101011100011101011010110001010010110;
            sine_reg0   <= 36'sb11000100111101000000001111111100111;
        end
        5904: begin
            cosine_reg0 <= 36'sb101011100011000100101011100100011011;
            sine_reg0   <= 36'sb11000100111000111111010011010010011;
        end
        5905: begin
            cosine_reg0 <= 36'sb101011100010011110000001110000111101;
            sine_reg0   <= 36'sb11000100110100111110001111000010000;
        end
        5906: begin
            cosine_reg0 <= 36'sb101011100001110111011000101111111110;
            sine_reg0   <= 36'sb11000100110000111101000011001100000;
        end
        5907: begin
            cosine_reg0 <= 36'sb101011100001010000110000100001100000;
            sine_reg0   <= 36'sb11000100101100111011101111110000101;
        end
        5908: begin
            cosine_reg0 <= 36'sb101011100000101010001001000101100101;
            sine_reg0   <= 36'sb11000100101000111010010100101111110;
        end
        5909: begin
            cosine_reg0 <= 36'sb101011100000000011100010011100001101;
            sine_reg0   <= 36'sb11000100100100111000110010001001110;
        end
        5910: begin
            cosine_reg0 <= 36'sb101011011111011100111100100101011001;
            sine_reg0   <= 36'sb11000100100000110111000111111110110;
        end
        5911: begin
            cosine_reg0 <= 36'sb101011011110110110010111100001001101;
            sine_reg0   <= 36'sb11000100011100110101010110001110110;
        end
        5912: begin
            cosine_reg0 <= 36'sb101011011110001111110011001111101000;
            sine_reg0   <= 36'sb11000100011000110011011100111010001;
        end
        5913: begin
            cosine_reg0 <= 36'sb101011011101101001001111110000101110;
            sine_reg0   <= 36'sb11000100010100110001011100000001000;
        end
        5914: begin
            cosine_reg0 <= 36'sb101011011101000010101101000100011110;
            sine_reg0   <= 36'sb11000100010000101111010011100011011;
        end
        5915: begin
            cosine_reg0 <= 36'sb101011011100011100001011001010111010;
            sine_reg0   <= 36'sb11000100001100101101000011100001100;
        end
        5916: begin
            cosine_reg0 <= 36'sb101011011011110101101010000100000101;
            sine_reg0   <= 36'sb11000100001000101010101011111011100;
        end
        5917: begin
            cosine_reg0 <= 36'sb101011011011001111001001101111111111;
            sine_reg0   <= 36'sb11000100000100101000001100110001101;
        end
        5918: begin
            cosine_reg0 <= 36'sb101011011010101000101010001110101011;
            sine_reg0   <= 36'sb11000100000000100101100110000011111;
        end
        5919: begin
            cosine_reg0 <= 36'sb101011011010000010001011100000001000;
            sine_reg0   <= 36'sb11000011111100100010110111110010100;
        end
        5920: begin
            cosine_reg0 <= 36'sb101011011001011011101101100100011010;
            sine_reg0   <= 36'sb11000011111000100000000001111101110;
        end
        5921: begin
            cosine_reg0 <= 36'sb101011011000110101010000011011100001;
            sine_reg0   <= 36'sb11000011110100011101000100100101101;
        end
        5922: begin
            cosine_reg0 <= 36'sb101011011000001110110100000101011111;
            sine_reg0   <= 36'sb11000011110000011001111111101010010;
        end
        5923: begin
            cosine_reg0 <= 36'sb101011010111101000011000100010010101;
            sine_reg0   <= 36'sb11000011101100010110110011001100000;
        end
        5924: begin
            cosine_reg0 <= 36'sb101011010111000001111101110010000101;
            sine_reg0   <= 36'sb11000011101000010011011111001010110;
        end
        5925: begin
            cosine_reg0 <= 36'sb101011010110011011100011110100110001;
            sine_reg0   <= 36'sb11000011100100010000000011100111000;
        end
        5926: begin
            cosine_reg0 <= 36'sb101011010101110101001010101010011010;
            sine_reg0   <= 36'sb11000011100000001100100000100000100;
        end
        5927: begin
            cosine_reg0 <= 36'sb101011010101001110110010010011000000;
            sine_reg0   <= 36'sb11000011011100001000110101110111110;
        end
        5928: begin
            cosine_reg0 <= 36'sb101011010100101000011010101110100111;
            sine_reg0   <= 36'sb11000011011000000101000011101100110;
        end
        5929: begin
            cosine_reg0 <= 36'sb101011010100000010000011111101001111;
            sine_reg0   <= 36'sb11000011010100000001001001111111101;
        end
        5930: begin
            cosine_reg0 <= 36'sb101011010011011011101101111110111001;
            sine_reg0   <= 36'sb11000011001111111101001000110000101;
        end
        5931: begin
            cosine_reg0 <= 36'sb101011010010110101011000110011101000;
            sine_reg0   <= 36'sb11000011001011111000111111111111111;
        end
        5932: begin
            cosine_reg0 <= 36'sb101011010010001111000100011011011101;
            sine_reg0   <= 36'sb11000011000111110100101111101101100;
        end
        5933: begin
            cosine_reg0 <= 36'sb101011010001101000110000110110011000;
            sine_reg0   <= 36'sb11000011000011110000010111111001110;
        end
        5934: begin
            cosine_reg0 <= 36'sb101011010001000010011110000100011101;
            sine_reg0   <= 36'sb11000010111111101011111000100100101;
        end
        5935: begin
            cosine_reg0 <= 36'sb101011010000011100001100000101101011;
            sine_reg0   <= 36'sb11000010111011100111010001101110011;
        end
        5936: begin
            cosine_reg0 <= 36'sb101011001111110101111010111010000110;
            sine_reg0   <= 36'sb11000010110111100010100011010111010;
        end
        5937: begin
            cosine_reg0 <= 36'sb101011001111001111101010100001101101;
            sine_reg0   <= 36'sb11000010110011011101101101011111001;
        end
        5938: begin
            cosine_reg0 <= 36'sb101011001110101001011010111100100011;
            sine_reg0   <= 36'sb11000010101111011000110000000110100;
        end
        5939: begin
            cosine_reg0 <= 36'sb101011001110000011001100001010101001;
            sine_reg0   <= 36'sb11000010101011010011101011001101011;
        end
        5940: begin
            cosine_reg0 <= 36'sb101011001101011100111110001100000000;
            sine_reg0   <= 36'sb11000010100111001110011110110011110;
        end
        5941: begin
            cosine_reg0 <= 36'sb101011001100110110110001000000101011;
            sine_reg0   <= 36'sb11000010100011001001001010111010001;
        end
        5942: begin
            cosine_reg0 <= 36'sb101011001100010000100100101000101001;
            sine_reg0   <= 36'sb11000010011111000011101111100000011;
        end
        5943: begin
            cosine_reg0 <= 36'sb101011001011101010011001000011111110;
            sine_reg0   <= 36'sb11000010011010111110001100100110110;
        end
        5944: begin
            cosine_reg0 <= 36'sb101011001011000100001110010010101010;
            sine_reg0   <= 36'sb11000010010110111000100010001101011;
        end
        5945: begin
            cosine_reg0 <= 36'sb101011001010011110000100010100110000;
            sine_reg0   <= 36'sb11000010010010110010110000010100100;
        end
        5946: begin
            cosine_reg0 <= 36'sb101011001001110111111011001010001111;
            sine_reg0   <= 36'sb11000010001110101100110110111100010;
        end
        5947: begin
            cosine_reg0 <= 36'sb101011001001010001110010110011001010;
            sine_reg0   <= 36'sb11000010001010100110110110000100101;
        end
        5948: begin
            cosine_reg0 <= 36'sb101011001000101011101011001111100011;
            sine_reg0   <= 36'sb11000010000110100000101101101110000;
        end
        5949: begin
            cosine_reg0 <= 36'sb101011001000000101100100011111011010;
            sine_reg0   <= 36'sb11000010000010011010011101111000100;
        end
        5950: begin
            cosine_reg0 <= 36'sb101011000111011111011110100010110010;
            sine_reg0   <= 36'sb11000001111110010100000110100100010;
        end
        5951: begin
            cosine_reg0 <= 36'sb101011000110111001011001011001101011;
            sine_reg0   <= 36'sb11000001111010001101100111110001010;
        end
        5952: begin
            cosine_reg0 <= 36'sb101011000110010011010101000100001000;
            sine_reg0   <= 36'sb11000001110110000111000001011111111;
        end
        5953: begin
            cosine_reg0 <= 36'sb101011000101101101010001100010001001;
            sine_reg0   <= 36'sb11000001110010000000010011110000010;
        end
        5954: begin
            cosine_reg0 <= 36'sb101011000101000111001110110011110000;
            sine_reg0   <= 36'sb11000001101101111001011110100010011;
        end
        5955: begin
            cosine_reg0 <= 36'sb101011000100100001001100111000111111;
            sine_reg0   <= 36'sb11000001101001110010100001110110101;
        end
        5956: begin
            cosine_reg0 <= 36'sb101011000011111011001011110001110111;
            sine_reg0   <= 36'sb11000001100101101011011101101101000;
        end
        5957: begin
            cosine_reg0 <= 36'sb101011000011010101001011011110011001;
            sine_reg0   <= 36'sb11000001100001100100010010000101110;
        end
        5958: begin
            cosine_reg0 <= 36'sb101011000010101111001011111110100111;
            sine_reg0   <= 36'sb11000001011101011100111111000001000;
        end
        5959: begin
            cosine_reg0 <= 36'sb101011000010001001001101010010100011;
            sine_reg0   <= 36'sb11000001011001010101100100011110111;
        end
        5960: begin
            cosine_reg0 <= 36'sb101011000001100011001111011010001101;
            sine_reg0   <= 36'sb11000001010101001110000010011111101;
        end
        5961: begin
            cosine_reg0 <= 36'sb101011000000111101010010010101101000;
            sine_reg0   <= 36'sb11000001010001000110011001000011010;
        end
        5962: begin
            cosine_reg0 <= 36'sb101011000000010111010110000100110101;
            sine_reg0   <= 36'sb11000001001100111110101000001010000;
        end
        5963: begin
            cosine_reg0 <= 36'sb101010111111110001011010100111110101;
            sine_reg0   <= 36'sb11000001001000110110101111110100001;
        end
        5964: begin
            cosine_reg0 <= 36'sb101010111111001011011111111110101010;
            sine_reg0   <= 36'sb11000001000100101110110000000001110;
        end
        5965: begin
            cosine_reg0 <= 36'sb101010111110100101100110001001010101;
            sine_reg0   <= 36'sb11000001000000100110101000110010111;
        end
        5966: begin
            cosine_reg0 <= 36'sb101010111101111111101101000111111000;
            sine_reg0   <= 36'sb11000000111100011110011010000111110;
        end
        5967: begin
            cosine_reg0 <= 36'sb101010111101011001110100111010010100;
            sine_reg0   <= 36'sb11000000111000010110000100000000101;
        end
        5968: begin
            cosine_reg0 <= 36'sb101010111100110011111101100000101010;
            sine_reg0   <= 36'sb11000000110100001101100110011101101;
        end
        5969: begin
            cosine_reg0 <= 36'sb101010111100001110000110111010111101;
            sine_reg0   <= 36'sb11000000110000000101000001011110110;
        end
        5970: begin
            cosine_reg0 <= 36'sb101010111011101000010001001001001101;
            sine_reg0   <= 36'sb11000000101011111100010101000100011;
        end
        5971: begin
            cosine_reg0 <= 36'sb101010111011000010011100001011011100;
            sine_reg0   <= 36'sb11000000100111110011100001001110100;
        end
        5972: begin
            cosine_reg0 <= 36'sb101010111010011100101000000001101011;
            sine_reg0   <= 36'sb11000000100011101010100101111101011;
        end
        5973: begin
            cosine_reg0 <= 36'sb101010111001110110110100101011111100;
            sine_reg0   <= 36'sb11000000011111100001100011010001001;
        end
        5974: begin
            cosine_reg0 <= 36'sb101010111001010001000010001010010001;
            sine_reg0   <= 36'sb11000000011011011000011001001010000;
        end
        5975: begin
            cosine_reg0 <= 36'sb101010111000101011010000011100101011;
            sine_reg0   <= 36'sb11000000010111001111000111101000000;
        end
        5976: begin
            cosine_reg0 <= 36'sb101010111000000101011111100011001010;
            sine_reg0   <= 36'sb11000000010011000101101110101011011;
        end
        5977: begin
            cosine_reg0 <= 36'sb101010110111011111101111011101110010;
            sine_reg0   <= 36'sb11000000001110111100001110010100010;
        end
        5978: begin
            cosine_reg0 <= 36'sb101010110110111010000000001100100010;
            sine_reg0   <= 36'sb11000000001010110010100110100010111;
        end
        5979: begin
            cosine_reg0 <= 36'sb101010110110010100010001101111011101;
            sine_reg0   <= 36'sb11000000000110101000110111010111010;
        end
        5980: begin
            cosine_reg0 <= 36'sb101010110101101110100100000110100101;
            sine_reg0   <= 36'sb11000000000010011111000000110001101;
        end
        5981: begin
            cosine_reg0 <= 36'sb101010110101001000110111010001111010;
            sine_reg0   <= 36'sb10111111111110010101000010110010010;
        end
        5982: begin
            cosine_reg0 <= 36'sb101010110100100011001011010001011101;
            sine_reg0   <= 36'sb10111111111010001010111101011001010;
        end
        5983: begin
            cosine_reg0 <= 36'sb101010110011111101100000000101010010;
            sine_reg0   <= 36'sb10111111110110000000110000100110101;
        end
        5984: begin
            cosine_reg0 <= 36'sb101010110011010111110101101101011000;
            sine_reg0   <= 36'sb10111111110001110110011100011010101;
        end
        5985: begin
            cosine_reg0 <= 36'sb101010110010110010001100001001110001;
            sine_reg0   <= 36'sb10111111101101101100000000110101100;
        end
        5986: begin
            cosine_reg0 <= 36'sb101010110010001100100011011010100000;
            sine_reg0   <= 36'sb10111111101001100001011101110111010;
        end
        5987: begin
            cosine_reg0 <= 36'sb101010110001100110111011011111100100;
            sine_reg0   <= 36'sb10111111100101010110110011100000010;
        end
        5988: begin
            cosine_reg0 <= 36'sb101010110001000001010100011001000000;
            sine_reg0   <= 36'sb10111111100001001100000001110000100;
        end
        5989: begin
            cosine_reg0 <= 36'sb101010110000011011101110000110110110;
            sine_reg0   <= 36'sb10111111011101000001001000101000001;
        end
        5990: begin
            cosine_reg0 <= 36'sb101010101111110110001000101001000110;
            sine_reg0   <= 36'sb10111111011000110110001000000111011;
        end
        5991: begin
            cosine_reg0 <= 36'sb101010101111010000100011111111110010;
            sine_reg0   <= 36'sb10111111010100101011000000001110100;
        end
        5992: begin
            cosine_reg0 <= 36'sb101010101110101011000000001010111011;
            sine_reg0   <= 36'sb10111111010000011111110000111101011;
        end
        5993: begin
            cosine_reg0 <= 36'sb101010101110000101011101001010100100;
            sine_reg0   <= 36'sb10111111001100010100011010010100100;
        end
        5994: begin
            cosine_reg0 <= 36'sb101010101101011111111010111110101101;
            sine_reg0   <= 36'sb10111111001000001000111100010011110;
        end
        5995: begin
            cosine_reg0 <= 36'sb101010101100111010011001100111010111;
            sine_reg0   <= 36'sb10111111000011111101010110111011100;
        end
        5996: begin
            cosine_reg0 <= 36'sb101010101100010100111001000100100101;
            sine_reg0   <= 36'sb10111110111111110001101010001011111;
        end
        5997: begin
            cosine_reg0 <= 36'sb101010101011101111011001010110011000;
            sine_reg0   <= 36'sb10111110111011100101110110000100111;
        end
        5998: begin
            cosine_reg0 <= 36'sb101010101011001001111010011100110001;
            sine_reg0   <= 36'sb10111110110111011001111010100110110;
        end
        5999: begin
            cosine_reg0 <= 36'sb101010101010100100011100010111110001;
            sine_reg0   <= 36'sb10111110110011001101110111110001110;
        end
        6000: begin
            cosine_reg0 <= 36'sb101010101001111110111111000111011011;
            sine_reg0   <= 36'sb10111110101111000001101101100110000;
        end
        6001: begin
            cosine_reg0 <= 36'sb101010101001011001100010101011101111;
            sine_reg0   <= 36'sb10111110101010110101011100000011101;
        end
        6002: begin
            cosine_reg0 <= 36'sb101010101000110100000111000100101111;
            sine_reg0   <= 36'sb10111110100110101001000011001010110;
        end
        6003: begin
            cosine_reg0 <= 36'sb101010101000001110101100010010011100;
            sine_reg0   <= 36'sb10111110100010011100100010111011101;
        end
        6004: begin
            cosine_reg0 <= 36'sb101010100111101001010010010100111001;
            sine_reg0   <= 36'sb10111110011110001111111011010110010;
        end
        6005: begin
            cosine_reg0 <= 36'sb101010100111000011111001001100000101;
            sine_reg0   <= 36'sb10111110011010000011001100011011000;
        end
        6006: begin
            cosine_reg0 <= 36'sb101010100110011110100000111000000011;
            sine_reg0   <= 36'sb10111110010101110110010110001001111;
        end
        6007: begin
            cosine_reg0 <= 36'sb101010100101111001001001011000110101;
            sine_reg0   <= 36'sb10111110010001101001011000100011010;
        end
        6008: begin
            cosine_reg0 <= 36'sb101010100101010011110010101110011011;
            sine_reg0   <= 36'sb10111110001101011100010011100111000;
        end
        6009: begin
            cosine_reg0 <= 36'sb101010100100101110011100111000110111;
            sine_reg0   <= 36'sb10111110001001001111000111010101100;
        end
        6010: begin
            cosine_reg0 <= 36'sb101010100100001001000111111000001010;
            sine_reg0   <= 36'sb10111110000101000001110011101110110;
        end
        6011: begin
            cosine_reg0 <= 36'sb101010100011100011110011101100010111;
            sine_reg0   <= 36'sb10111110000000110100011000110011000;
        end
        6012: begin
            cosine_reg0 <= 36'sb101010100010111110100000010101011110;
            sine_reg0   <= 36'sb10111101111100100110110110100010100;
        end
        6013: begin
            cosine_reg0 <= 36'sb101010100010011001001101110011100000;
            sine_reg0   <= 36'sb10111101111000011001001100111101010;
        end
        6014: begin
            cosine_reg0 <= 36'sb101010100001110011111100000110100000;
            sine_reg0   <= 36'sb10111101110100001011011100000011101;
        end
        6015: begin
            cosine_reg0 <= 36'sb101010100001001110101011001110011111;
            sine_reg0   <= 36'sb10111101101111111101100011110101100;
        end
        6016: begin
            cosine_reg0 <= 36'sb101010100000101001011011001011011101;
            sine_reg0   <= 36'sb10111101101011101111100100010011010;
        end
        6017: begin
            cosine_reg0 <= 36'sb101010100000000100001011111101011110;
            sine_reg0   <= 36'sb10111101100111100001011101011101000;
        end
        6018: begin
            cosine_reg0 <= 36'sb101010011111011110111101100100100001;
            sine_reg0   <= 36'sb10111101100011010011001111010010110;
        end
        6019: begin
            cosine_reg0 <= 36'sb101010011110111001110000000000101000;
            sine_reg0   <= 36'sb10111101011111000100111001110101000;
        end
        6020: begin
            cosine_reg0 <= 36'sb101010011110010100100011010001110110;
            sine_reg0   <= 36'sb10111101011010110110011101000011100;
        end
        6021: begin
            cosine_reg0 <= 36'sb101010011101101111010111011000001011;
            sine_reg0   <= 36'sb10111101010110100111111000111110110;
        end
        6022: begin
            cosine_reg0 <= 36'sb101010011101001010001100010011101000;
            sine_reg0   <= 36'sb10111101010010011001001101100110111;
        end
        6023: begin
            cosine_reg0 <= 36'sb101010011100100101000010000100010000;
            sine_reg0   <= 36'sb10111101001110001010011010111011110;
        end
        6024: begin
            cosine_reg0 <= 36'sb101010011011111111111000101010000011;
            sine_reg0   <= 36'sb10111101001001111011100000111101111;
        end
        6025: begin
            cosine_reg0 <= 36'sb101010011011011010110000000101000011;
            sine_reg0   <= 36'sb10111101000101101100011111101101010;
        end
        6026: begin
            cosine_reg0 <= 36'sb101010011010110101101000010101010010;
            sine_reg0   <= 36'sb10111101000001011101010111001010001;
        end
        6027: begin
            cosine_reg0 <= 36'sb101010011010010000100001011010110000;
            sine_reg0   <= 36'sb10111100111101001110000111010100100;
        end
        6028: begin
            cosine_reg0 <= 36'sb101010011001101011011011010101100000;
            sine_reg0   <= 36'sb10111100111000111110110000001100101;
        end
        6029: begin
            cosine_reg0 <= 36'sb101010011001000110010110000101100011;
            sine_reg0   <= 36'sb10111100110100101111010001110010110;
        end
        6030: begin
            cosine_reg0 <= 36'sb101010011000100001010001101010111010;
            sine_reg0   <= 36'sb10111100110000011111101100000111000;
        end
        6031: begin
            cosine_reg0 <= 36'sb101010010111111100001110000101100110;
            sine_reg0   <= 36'sb10111100101100001111111111001001100;
        end
        6032: begin
            cosine_reg0 <= 36'sb101010010111010111001011010101101001;
            sine_reg0   <= 36'sb10111100101000000000001010111010011;
        end
        6033: begin
            cosine_reg0 <= 36'sb101010010110110010001001011011000101;
            sine_reg0   <= 36'sb10111100100011110000001111011001111;
        end
        6034: begin
            cosine_reg0 <= 36'sb101010010110001101001000010101111011;
            sine_reg0   <= 36'sb10111100011111100000001100101000001;
        end
        6035: begin
            cosine_reg0 <= 36'sb101010010101101000001000000110001100;
            sine_reg0   <= 36'sb10111100011011010000000010100101010;
        end
        6036: begin
            cosine_reg0 <= 36'sb101010010101000011001000101011111010;
            sine_reg0   <= 36'sb10111100010110111111110001010001100;
        end
        6037: begin
            cosine_reg0 <= 36'sb101010010100011110001010000111000110;
            sine_reg0   <= 36'sb10111100010010101111011000101101000;
        end
        6038: begin
            cosine_reg0 <= 36'sb101010010011111001001100010111110001;
            sine_reg0   <= 36'sb10111100001110011110111000110111110;
        end
        6039: begin
            cosine_reg0 <= 36'sb101010010011010100001111011101111110;
            sine_reg0   <= 36'sb10111100001010001110010001110010010;
        end
        6040: begin
            cosine_reg0 <= 36'sb101010010010101111010011011001101101;
            sine_reg0   <= 36'sb10111100000101111101100011011100011;
        end
        6041: begin
            cosine_reg0 <= 36'sb101010010010001010011000001011000000;
            sine_reg0   <= 36'sb10111100000001101100101101110110100;
        end
        6042: begin
            cosine_reg0 <= 36'sb101010010001100101011101110001111000;
            sine_reg0   <= 36'sb10111011111101011011110001000000101;
        end
        6043: begin
            cosine_reg0 <= 36'sb101010010001000000100100001110010111;
            sine_reg0   <= 36'sb10111011111001001010101100111011000;
        end
        6044: begin
            cosine_reg0 <= 36'sb101010010000011011101011100000011110;
            sine_reg0   <= 36'sb10111011110100111001100001100101110;
        end
        6045: begin
            cosine_reg0 <= 36'sb101010001111110110110011101000001110;
            sine_reg0   <= 36'sb10111011110000101000001111000001001;
        end
        6046: begin
            cosine_reg0 <= 36'sb101010001111010001111100100101101010;
            sine_reg0   <= 36'sb10111011101100010110110101001101001;
        end
        6047: begin
            cosine_reg0 <= 36'sb101010001110101101000110011000110010;
            sine_reg0   <= 36'sb10111011101000000101010100001010000;
        end
        6048: begin
            cosine_reg0 <= 36'sb101010001110001000010001000001100111;
            sine_reg0   <= 36'sb10111011100011110011101011111000000;
        end
        6049: begin
            cosine_reg0 <= 36'sb101010001101100011011100100000001100;
            sine_reg0   <= 36'sb10111011011111100001111100010111010;
        end
        6050: begin
            cosine_reg0 <= 36'sb101010001100111110101000110100100010;
            sine_reg0   <= 36'sb10111011011011010000000101100111110;
        end
        6051: begin
            cosine_reg0 <= 36'sb101010001100011001110101111110101010;
            sine_reg0   <= 36'sb10111011010110111110000111101001111;
        end
        6052: begin
            cosine_reg0 <= 36'sb101010001011110101000011111110100101;
            sine_reg0   <= 36'sb10111011010010101100000010011101110;
        end
        6053: begin
            cosine_reg0 <= 36'sb101010001011010000010010110100010101;
            sine_reg0   <= 36'sb10111011001110011001110110000011011;
        end
        6054: begin
            cosine_reg0 <= 36'sb101010001010101011100010011111111100;
            sine_reg0   <= 36'sb10111011001010000111100010011011001;
        end
        6055: begin
            cosine_reg0 <= 36'sb101010001010000110110011000001011010;
            sine_reg0   <= 36'sb10111011000101110101000111100101001;
        end
        6056: begin
            cosine_reg0 <= 36'sb101010001001100010000100011000110001;
            sine_reg0   <= 36'sb10111011000001100010100101100001011;
        end
        6057: begin
            cosine_reg0 <= 36'sb101010001000111101010110100110000011;
            sine_reg0   <= 36'sb10111010111101001111111100010000010;
        end
        6058: begin
            cosine_reg0 <= 36'sb101010001000011000101001101001010001;
            sine_reg0   <= 36'sb10111010111000111101001011110001111;
        end
        6059: begin
            cosine_reg0 <= 36'sb101010000111110011111101100010011100;
            sine_reg0   <= 36'sb10111010110100101010010100000110010;
        end
        6060: begin
            cosine_reg0 <= 36'sb101010000111001111010010010001100111;
            sine_reg0   <= 36'sb10111010110000010111010101001101110;
        end
        6061: begin
            cosine_reg0 <= 36'sb101010000110101010100111110110110001;
            sine_reg0   <= 36'sb10111010101100000100001111001000011;
        end
        6062: begin
            cosine_reg0 <= 36'sb101010000110000101111110010001111101;
            sine_reg0   <= 36'sb10111010100111110001000001110110011;
        end
        6063: begin
            cosine_reg0 <= 36'sb101010000101100001010101100011001100;
            sine_reg0   <= 36'sb10111010100011011101101101011000000;
        end
        6064: begin
            cosine_reg0 <= 36'sb101010000100111100101101101010100000;
            sine_reg0   <= 36'sb10111010011111001010010001101101001;
        end
        6065: begin
            cosine_reg0 <= 36'sb101010000100011000000110100111111001;
            sine_reg0   <= 36'sb10111010011010110110101110110110010;
        end
        6066: begin
            cosine_reg0 <= 36'sb101010000011110011100000011011011010;
            sine_reg0   <= 36'sb10111010010110100011000100110011011;
        end
        6067: begin
            cosine_reg0 <= 36'sb101010000011001110111011000101000100;
            sine_reg0   <= 36'sb10111010010010001111010011100100110;
        end
        6068: begin
            cosine_reg0 <= 36'sb101010000010101010010110100100110111;
            sine_reg0   <= 36'sb10111010001101111011011011001010100;
        end
        6069: begin
            cosine_reg0 <= 36'sb101010000010000101110010111010110111;
            sine_reg0   <= 36'sb10111010001001100111011011100100101;
        end
        6070: begin
            cosine_reg0 <= 36'sb101010000001100001010000000111000011;
            sine_reg0   <= 36'sb10111010000101010011010100110011101;
        end
        6071: begin
            cosine_reg0 <= 36'sb101010000000111100101110001001011101;
            sine_reg0   <= 36'sb10111010000000111111000110110111011;
        end
        6072: begin
            cosine_reg0 <= 36'sb101010000000011000001101000010000111;
            sine_reg0   <= 36'sb10111001111100101010110001110000001;
        end
        6073: begin
            cosine_reg0 <= 36'sb101001111111110011101100110001000011;
            sine_reg0   <= 36'sb10111001111000010110010101011110001;
        end
        6074: begin
            cosine_reg0 <= 36'sb101001111111001111001101010110010001;
            sine_reg0   <= 36'sb10111001110100000001110010000001100;
        end
        6075: begin
            cosine_reg0 <= 36'sb101001111110101010101110110001110011;
            sine_reg0   <= 36'sb10111001101111101101000111011010011;
        end
        6076: begin
            cosine_reg0 <= 36'sb101001111110000110010001000011101010;
            sine_reg0   <= 36'sb10111001101011011000010101101000111;
        end
        6077: begin
            cosine_reg0 <= 36'sb101001111101100001110100001011111000;
            sine_reg0   <= 36'sb10111001100111000011011100101101011;
        end
        6078: begin
            cosine_reg0 <= 36'sb101001111100111101011000001010011110;
            sine_reg0   <= 36'sb10111001100010101110011100100111110;
        end
        6079: begin
            cosine_reg0 <= 36'sb101001111100011000111100111111011110;
            sine_reg0   <= 36'sb10111001011110011001010101011000011;
        end
        6080: begin
            cosine_reg0 <= 36'sb101001111011110100100010101010111001;
            sine_reg0   <= 36'sb10111001011010000100000110111111011;
        end
        6081: begin
            cosine_reg0 <= 36'sb101001111011010000001001001100110001;
            sine_reg0   <= 36'sb10111001010101101110110001011100111;
        end
        6082: begin
            cosine_reg0 <= 36'sb101001111010101011110000100101000110;
            sine_reg0   <= 36'sb10111001010001011001010100110001001;
        end
        6083: begin
            cosine_reg0 <= 36'sb101001111010000111011000110011111010;
            sine_reg0   <= 36'sb10111001001101000011110000111100010;
        end
        6084: begin
            cosine_reg0 <= 36'sb101001111001100011000001111001001111;
            sine_reg0   <= 36'sb10111001001000101110000101111110011;
        end
        6085: begin
            cosine_reg0 <= 36'sb101001111000111110101011110101000110;
            sine_reg0   <= 36'sb10111001000100011000010011110111101;
        end
        6086: begin
            cosine_reg0 <= 36'sb101001111000011010010110100111100001;
            sine_reg0   <= 36'sb10111001000000000010011010101000010;
        end
        6087: begin
            cosine_reg0 <= 36'sb101001110111110110000010010000100000;
            sine_reg0   <= 36'sb10111000111011101100011010010000100;
        end
        6088: begin
            cosine_reg0 <= 36'sb101001110111010001101110110000000110;
            sine_reg0   <= 36'sb10111000110111010110010010110000011;
        end
        6089: begin
            cosine_reg0 <= 36'sb101001110110101101011100000110010011;
            sine_reg0   <= 36'sb10111000110011000000000100001000001;
        end
        6090: begin
            cosine_reg0 <= 36'sb101001110110001001001010010011001001;
            sine_reg0   <= 36'sb10111000101110101001101110010111111;
        end
        6091: begin
            cosine_reg0 <= 36'sb101001110101100100111001010110101010;
            sine_reg0   <= 36'sb10111000101010010011010001011111111;
        end
        6092: begin
            cosine_reg0 <= 36'sb101001110101000000101001010000110110;
            sine_reg0   <= 36'sb10111000100101111100101101100000010;
        end
        6093: begin
            cosine_reg0 <= 36'sb101001110100011100011010000001110000;
            sine_reg0   <= 36'sb10111000100001100110000010011001001;
        end
        6094: begin
            cosine_reg0 <= 36'sb101001110011111000001011101001011000;
            sine_reg0   <= 36'sb10111000011101001111010000001010101;
        end
        6095: begin
            cosine_reg0 <= 36'sb101001110011010011111110000111110000;
            sine_reg0   <= 36'sb10111000011000111000010110110101001;
        end
        6096: begin
            cosine_reg0 <= 36'sb101001110010101111110001011100111010;
            sine_reg0   <= 36'sb10111000010100100001010110011000101;
        end
        6097: begin
            cosine_reg0 <= 36'sb101001110010001011100101101000110110;
            sine_reg0   <= 36'sb10111000010000001010001110110101011;
        end
        6098: begin
            cosine_reg0 <= 36'sb101001110001100111011010101011100111;
            sine_reg0   <= 36'sb10111000001011110011000000001011011;
        end
        6099: begin
            cosine_reg0 <= 36'sb101001110001000011010000100101001101;
            sine_reg0   <= 36'sb10111000000111011011101010011011000;
        end
        6100: begin
            cosine_reg0 <= 36'sb101001110000011111000111010101101010;
            sine_reg0   <= 36'sb10111000000011000100001101100100011;
        end
        6101: begin
            cosine_reg0 <= 36'sb101001101111111010111110111101000000;
            sine_reg0   <= 36'sb10110111111110101100101001100111101;
        end
        6102: begin
            cosine_reg0 <= 36'sb101001101111010110110111011011001111;
            sine_reg0   <= 36'sb10110111111010010100111110100100111;
        end
        6103: begin
            cosine_reg0 <= 36'sb101001101110110010110000110000011010;
            sine_reg0   <= 36'sb10110111110101111101001100011100011;
        end
        6104: begin
            cosine_reg0 <= 36'sb101001101110001110101010111100100001;
            sine_reg0   <= 36'sb10110111110001100101010011001110010;
        end
        6105: begin
            cosine_reg0 <= 36'sb101001101101101010100101111111100110;
            sine_reg0   <= 36'sb10110111101101001101010010111010101;
        end
        6106: begin
            cosine_reg0 <= 36'sb101001101101000110100001111001101010;
            sine_reg0   <= 36'sb10110111101000110101001011100001110;
        end
        6107: begin
            cosine_reg0 <= 36'sb101001101100100010011110101010101111;
            sine_reg0   <= 36'sb10110111100100011100111101000011110;
        end
        6108: begin
            cosine_reg0 <= 36'sb101001101011111110011100010010110111;
            sine_reg0   <= 36'sb10110111100000000100100111100000111;
        end
        6109: begin
            cosine_reg0 <= 36'sb101001101011011010011010110010000001;
            sine_reg0   <= 36'sb10110111011011101100001010111001010;
        end
        6110: begin
            cosine_reg0 <= 36'sb101001101010110110011010001000010001;
            sine_reg0   <= 36'sb10110111010111010011100111001100111;
        end
        6111: begin
            cosine_reg0 <= 36'sb101001101010010010011010010101100111;
            sine_reg0   <= 36'sb10110111010010111010111100011100010;
        end
        6112: begin
            cosine_reg0 <= 36'sb101001101001101110011011011010000101;
            sine_reg0   <= 36'sb10110111001110100010001010100111010;
        end
        6113: begin
            cosine_reg0 <= 36'sb101001101001001010011101010101101011;
            sine_reg0   <= 36'sb10110111001010001001010001101110001;
        end
        6114: begin
            cosine_reg0 <= 36'sb101001101000100110100000001000011100;
            sine_reg0   <= 36'sb10110111000101110000010001110001001;
        end
        6115: begin
            cosine_reg0 <= 36'sb101001101000000010100011110010011001;
            sine_reg0   <= 36'sb10110111000001010111001010110000011;
        end
        6116: begin
            cosine_reg0 <= 36'sb101001100111011110101000010011100011;
            sine_reg0   <= 36'sb10110110111100111101111100101100001;
        end
        6117: begin
            cosine_reg0 <= 36'sb101001100110111010101101101011111100;
            sine_reg0   <= 36'sb10110110111000100100100111100100011;
        end
        6118: begin
            cosine_reg0 <= 36'sb101001100110010110110011111011100101;
            sine_reg0   <= 36'sb10110110110100001011001011011001011;
        end
        6119: begin
            cosine_reg0 <= 36'sb101001100101110010111011000010011111;
            sine_reg0   <= 36'sb10110110101111110001101000001011010;
        end
        6120: begin
            cosine_reg0 <= 36'sb101001100101001111000011000000101100;
            sine_reg0   <= 36'sb10110110101011010111111101111010010;
        end
        6121: begin
            cosine_reg0 <= 36'sb101001100100101011001011110110001101;
            sine_reg0   <= 36'sb10110110100110111110001100100110100;
        end
        6122: begin
            cosine_reg0 <= 36'sb101001100100000111010101100011000100;
            sine_reg0   <= 36'sb10110110100010100100010100010000010;
        end
        6123: begin
            cosine_reg0 <= 36'sb101001100011100011100000000111010001;
            sine_reg0   <= 36'sb10110110011110001010010100110111100;
        end
        6124: begin
            cosine_reg0 <= 36'sb101001100010111111101011100010110111;
            sine_reg0   <= 36'sb10110110011001110000001110011100101;
        end
        6125: begin
            cosine_reg0 <= 36'sb101001100010011011110111110101110110;
            sine_reg0   <= 36'sb10110110010101010110000000111111101;
        end
        6126: begin
            cosine_reg0 <= 36'sb101001100001111000000101000000010001;
            sine_reg0   <= 36'sb10110110010000111011101100100000110;
        end
        6127: begin
            cosine_reg0 <= 36'sb101001100001010100010011000010001000;
            sine_reg0   <= 36'sb10110110001100100001010001000000001;
        end
        6128: begin
            cosine_reg0 <= 36'sb101001100000110000100001111011011100;
            sine_reg0   <= 36'sb10110110001000000110101110011110000;
        end
        6129: begin
            cosine_reg0 <= 36'sb101001100000001100110001101100010000;
            sine_reg0   <= 36'sb10110110000011101100000100111010011;
        end
        6130: begin
            cosine_reg0 <= 36'sb101001011111101001000010010100100101;
            sine_reg0   <= 36'sb10110101111111010001010100010101110;
        end
        6131: begin
            cosine_reg0 <= 36'sb101001011111000101010011110100011011;
            sine_reg0   <= 36'sb10110101111010110110011100101111111;
        end
        6132: begin
            cosine_reg0 <= 36'sb101001011110100001100110001011110101;
            sine_reg0   <= 36'sb10110101110110011011011110001001010;
        end
        6133: begin
            cosine_reg0 <= 36'sb101001011101111101111001011010110011;
            sine_reg0   <= 36'sb10110101110010000000011000100001111;
        end
        6134: begin
            cosine_reg0 <= 36'sb101001011101011010001101100001011000;
            sine_reg0   <= 36'sb10110101101101100101001011111010000;
        end
        6135: begin
            cosine_reg0 <= 36'sb101001011100110110100010011111100100;
            sine_reg0   <= 36'sb10110101101001001001111000010001111;
        end
        6136: begin
            cosine_reg0 <= 36'sb101001011100010010111000010101011000;
            sine_reg0   <= 36'sb10110101100100101110011101101001011;
        end
        6137: begin
            cosine_reg0 <= 36'sb101001011011101111001111000010110111;
            sine_reg0   <= 36'sb10110101100000010010111100000001000;
        end
        6138: begin
            cosine_reg0 <= 36'sb101001011011001011100110101000000010;
            sine_reg0   <= 36'sb10110101011011110111010011011000110;
        end
        6139: begin
            cosine_reg0 <= 36'sb101001011010100111111111000100111001;
            sine_reg0   <= 36'sb10110101010111011011100011110000110;
        end
        6140: begin
            cosine_reg0 <= 36'sb101001011010000100011000011001011111;
            sine_reg0   <= 36'sb10110101010010111111101101001001010;
        end
        6141: begin
            cosine_reg0 <= 36'sb101001011001100000110010100101110101;
            sine_reg0   <= 36'sb10110101001110100011101111100010100;
        end
        6142: begin
            cosine_reg0 <= 36'sb101001011000111101001101101001111011;
            sine_reg0   <= 36'sb10110101001010000111101010111100101;
        end
        6143: begin
            cosine_reg0 <= 36'sb101001011000011001101001100101110100;
            sine_reg0   <= 36'sb10110101000101101011011111010111101;
        end
        6144: begin
            cosine_reg0 <= 36'sb101001010111110110000110011001100001;
            sine_reg0   <= 36'sb10110101000001001111001100110011111;
        end
        6145: begin
            cosine_reg0 <= 36'sb101001010111010010100100000101000011;
            sine_reg0   <= 36'sb10110100111100110010110011010001100;
        end
        6146: begin
            cosine_reg0 <= 36'sb101001010110101111000010101000011011;
            sine_reg0   <= 36'sb10110100111000010110010010110000101;
        end
        6147: begin
            cosine_reg0 <= 36'sb101001010110001011100010000011101100;
            sine_reg0   <= 36'sb10110100110011111001101011010001011;
        end
        6148: begin
            cosine_reg0 <= 36'sb101001010101101000000010010110110110;
            sine_reg0   <= 36'sb10110100101111011100111100110100001;
        end
        6149: begin
            cosine_reg0 <= 36'sb101001010101000100100011100001111010;
            sine_reg0   <= 36'sb10110100101011000000000111011000111;
        end
        6150: begin
            cosine_reg0 <= 36'sb101001010100100001000101100100111010;
            sine_reg0   <= 36'sb10110100100110100011001010111111110;
        end
        6151: begin
            cosine_reg0 <= 36'sb101001010011111101101000011111111000;
            sine_reg0   <= 36'sb10110100100010000110000111101001001;
        end
        6152: begin
            cosine_reg0 <= 36'sb101001010011011010001100010010110101;
            sine_reg0   <= 36'sb10110100011101101000111101010101000;
        end
        6153: begin
            cosine_reg0 <= 36'sb101001010010110110110000111101110001;
            sine_reg0   <= 36'sb10110100011001001011101100000011100;
        end
        6154: begin
            cosine_reg0 <= 36'sb101001010010010011010110100000110000;
            sine_reg0   <= 36'sb10110100010100101110010011110101000;
        end
        6155: begin
            cosine_reg0 <= 36'sb101001010001101111111100111011110001;
            sine_reg0   <= 36'sb10110100010000010000110100101001101;
        end
        6156: begin
            cosine_reg0 <= 36'sb101001010001001100100100001110110110;
            sine_reg0   <= 36'sb10110100001011110011001110100001011;
        end
        6157: begin
            cosine_reg0 <= 36'sb101001010000101001001100011010000001;
            sine_reg0   <= 36'sb10110100000111010101100001011100101;
        end
        6158: begin
            cosine_reg0 <= 36'sb101001010000000101110101011101010010;
            sine_reg0   <= 36'sb10110100000010110111101101011011011;
        end
        6159: begin
            cosine_reg0 <= 36'sb101001001111100010011111011000101101;
            sine_reg0   <= 36'sb10110011111110011001110010011110000;
        end
        6160: begin
            cosine_reg0 <= 36'sb101001001110111111001010001100010000;
            sine_reg0   <= 36'sb10110011111001111011110000100100100;
        end
        6161: begin
            cosine_reg0 <= 36'sb101001001110011011110101110111111111;
            sine_reg0   <= 36'sb10110011110101011101100111101111000;
        end
        6162: begin
            cosine_reg0 <= 36'sb101001001101111000100010011011111010;
            sine_reg0   <= 36'sb10110011110000111111010111111101111;
        end
        6163: begin
            cosine_reg0 <= 36'sb101001001101010101001111111000000011;
            sine_reg0   <= 36'sb10110011101100100001000001010001010;
        end
        6164: begin
            cosine_reg0 <= 36'sb101001001100110001111110001100011011;
            sine_reg0   <= 36'sb10110011101000000010100011101001001;
        end
        6165: begin
            cosine_reg0 <= 36'sb101001001100001110101101011001000100;
            sine_reg0   <= 36'sb10110011100011100011111111000101111;
        end
        6166: begin
            cosine_reg0 <= 36'sb101001001011101011011101011101111110;
            sine_reg0   <= 36'sb10110011011111000101010011100111100;
        end
        6167: begin
            cosine_reg0 <= 36'sb101001001011001000001110011011001100;
            sine_reg0   <= 36'sb10110011011010100110100001001110011;
        end
        6168: begin
            cosine_reg0 <= 36'sb101001001010100101000000010000101110;
            sine_reg0   <= 36'sb10110011010110000111100111111010100;
        end
        6169: begin
            cosine_reg0 <= 36'sb101001001010000001110010111110100110;
            sine_reg0   <= 36'sb10110011010001101000100111101100001;
        end
        6170: begin
            cosine_reg0 <= 36'sb101001001001011110100110100100110101;
            sine_reg0   <= 36'sb10110011001101001001100000100011011;
        end
        6171: begin
            cosine_reg0 <= 36'sb101001001000111011011011000011011101;
            sine_reg0   <= 36'sb10110011001000101010010010100000100;
        end
        6172: begin
            cosine_reg0 <= 36'sb101001001000011000010000011010011111;
            sine_reg0   <= 36'sb10110011000100001010111101100011101;
        end
        6173: begin
            cosine_reg0 <= 36'sb101001000111110101000110101001111101;
            sine_reg0   <= 36'sb10110010111111101011100001101100111;
        end
        6174: begin
            cosine_reg0 <= 36'sb101001000111010001111101110001110111;
            sine_reg0   <= 36'sb10110010111011001011111110111100100;
        end
        6175: begin
            cosine_reg0 <= 36'sb101001000110101110110101110010001111;
            sine_reg0   <= 36'sb10110010110110101100010101010010101;
        end
        6176: begin
            cosine_reg0 <= 36'sb101001000110001011101110101011000110;
            sine_reg0   <= 36'sb10110010110010001100100100101111011;
        end
        6177: begin
            cosine_reg0 <= 36'sb101001000101101000101000011100011110;
            sine_reg0   <= 36'sb10110010101101101100101101010011001;
        end
        6178: begin
            cosine_reg0 <= 36'sb101001000101000101100011000110011001;
            sine_reg0   <= 36'sb10110010101001001100101110111101111;
        end
        6179: begin
            cosine_reg0 <= 36'sb101001000100100010011110101000110110;
            sine_reg0   <= 36'sb10110010100100101100101001101111111;
        end
        6180: begin
            cosine_reg0 <= 36'sb101001000011111111011011000011111001;
            sine_reg0   <= 36'sb10110010100000001100011101101001001;
        end
        6181: begin
            cosine_reg0 <= 36'sb101001000011011100011000010111100010;
            sine_reg0   <= 36'sb10110010011011101100001010101010001;
        end
        6182: begin
            cosine_reg0 <= 36'sb101001000010111001010110100011110010;
            sine_reg0   <= 36'sb10110010010111001011110000110010110;
        end
        6183: begin
            cosine_reg0 <= 36'sb101001000010010110010101101000101011;
            sine_reg0   <= 36'sb10110010010010101011010000000011010;
        end
        6184: begin
            cosine_reg0 <= 36'sb101001000001110011010101100110001110;
            sine_reg0   <= 36'sb10110010001110001010101000011011111;
        end
        6185: begin
            cosine_reg0 <= 36'sb101001000001010000010110011100011101;
            sine_reg0   <= 36'sb10110010001001101001111001111100110;
        end
        6186: begin
            cosine_reg0 <= 36'sb101001000000101101011000001011011001;
            sine_reg0   <= 36'sb10110010000101001001000100100110001;
        end
        6187: begin
            cosine_reg0 <= 36'sb101001000000001010011010110011000011;
            sine_reg0   <= 36'sb10110010000000101000001000011000000;
        end
        6188: begin
            cosine_reg0 <= 36'sb101000111111100111011110010011011101;
            sine_reg0   <= 36'sb10110001111100000111000101010010110;
        end
        6189: begin
            cosine_reg0 <= 36'sb101000111111000100100010101100101000;
            sine_reg0   <= 36'sb10110001110111100101111011010110011;
        end
        6190: begin
            cosine_reg0 <= 36'sb101000111110100001100111111110100101;
            sine_reg0   <= 36'sb10110001110011000100101010100011001;
        end
        6191: begin
            cosine_reg0 <= 36'sb101000111101111110101110001001010101;
            sine_reg0   <= 36'sb10110001101110100011010010111001010;
        end
        6192: begin
            cosine_reg0 <= 36'sb101000111101011011110101001100111011;
            sine_reg0   <= 36'sb10110001101010000001110100011000110;
        end
        6193: begin
            cosine_reg0 <= 36'sb101000111100111000111101001001010111;
            sine_reg0   <= 36'sb10110001100101100000001111000010000;
        end
        6194: begin
            cosine_reg0 <= 36'sb101000111100010110000101111110101011;
            sine_reg0   <= 36'sb10110001100000111110100010110101000;
        end
        6195: begin
            cosine_reg0 <= 36'sb101000111011110011001111101100110111;
            sine_reg0   <= 36'sb10110001011100011100101111110010000;
        end
        6196: begin
            cosine_reg0 <= 36'sb101000111011010000011010010011111110;
            sine_reg0   <= 36'sb10110001010111111010110101111001010;
        end
        6197: begin
            cosine_reg0 <= 36'sb101000111010101101100101110100000001;
            sine_reg0   <= 36'sb10110001010011011000110101001010110;
        end
        6198: begin
            cosine_reg0 <= 36'sb101000111010001010110010001101000001;
            sine_reg0   <= 36'sb10110001001110110110101101100110111;
        end
        6199: begin
            cosine_reg0 <= 36'sb101000111001100111111111011110111111;
            sine_reg0   <= 36'sb10110001001010010100011111001101101;
        end
        6200: begin
            cosine_reg0 <= 36'sb101000111001000101001101101001111101;
            sine_reg0   <= 36'sb10110001000101110010001001111111010;
        end
        6201: begin
            cosine_reg0 <= 36'sb101000111000100010011100101101111100;
            sine_reg0   <= 36'sb10110001000001001111101101111100000;
        end
        6202: begin
            cosine_reg0 <= 36'sb101000110111111111101100101010111110;
            sine_reg0   <= 36'sb10110000111100101101001011000011111;
        end
        6203: begin
            cosine_reg0 <= 36'sb101000110111011100111101100001000011;
            sine_reg0   <= 36'sb10110000111000001010100001010111010;
        end
        6204: begin
            cosine_reg0 <= 36'sb101000110110111010001111010000001101;
            sine_reg0   <= 36'sb10110000110011100111110000110110001;
        end
        6205: begin
            cosine_reg0 <= 36'sb101000110110010111100001111000011110;
            sine_reg0   <= 36'sb10110000101111000100111001100000110;
        end
        6206: begin
            cosine_reg0 <= 36'sb101000110101110100110101011001110111;
            sine_reg0   <= 36'sb10110000101010100001111011010111010;
        end
        6207: begin
            cosine_reg0 <= 36'sb101000110101010010001001110100011001;
            sine_reg0   <= 36'sb10110000100101111110110110011001111;
        end
        6208: begin
            cosine_reg0 <= 36'sb101000110100101111011111001000000101;
            sine_reg0   <= 36'sb10110000100001011011101010101000111;
        end
        6209: begin
            cosine_reg0 <= 36'sb101000110100001100110101010100111101;
            sine_reg0   <= 36'sb10110000011100111000011000000100010;
        end
        6210: begin
            cosine_reg0 <= 36'sb101000110011101010001100011011000010;
            sine_reg0   <= 36'sb10110000011000010100111110101100010;
        end
        6211: begin
            cosine_reg0 <= 36'sb101000110011000111100100011010010101;
            sine_reg0   <= 36'sb10110000010011110001011110100001000;
        end
        6212: begin
            cosine_reg0 <= 36'sb101000110010100100111101010010111001;
            sine_reg0   <= 36'sb10110000001111001101110111100010110;
        end
        6213: begin
            cosine_reg0 <= 36'sb101000110010000010010111000100101101;
            sine_reg0   <= 36'sb10110000001010101010001001110001101;
        end
        6214: begin
            cosine_reg0 <= 36'sb101000110001011111110001101111110100;
            sine_reg0   <= 36'sb10110000000110000110010101001101111;
        end
        6215: begin
            cosine_reg0 <= 36'sb101000110000111101001101010100001111;
            sine_reg0   <= 36'sb10110000000001100010011001110111101;
        end
        6216: begin
            cosine_reg0 <= 36'sb101000110000011010101001110001111111;
            sine_reg0   <= 36'sb10101111111100111110010111101111001;
        end
        6217: begin
            cosine_reg0 <= 36'sb101000101111111000000111001001000101;
            sine_reg0   <= 36'sb10101111111000011010001110110100011;
        end
        6218: begin
            cosine_reg0 <= 36'sb101000101111010101100101011001100011;
            sine_reg0   <= 36'sb10101111110011110101111111000111101;
        end
        6219: begin
            cosine_reg0 <= 36'sb101000101110110011000100100011011011;
            sine_reg0   <= 36'sb10101111101111010001101000101001001;
        end
        6220: begin
            cosine_reg0 <= 36'sb101000101110010000100100100110101100;
            sine_reg0   <= 36'sb10101111101010101101001011011001001;
        end
        6221: begin
            cosine_reg0 <= 36'sb101000101101101110000101100011011010;
            sine_reg0   <= 36'sb10101111100110001000100111010111100;
        end
        6222: begin
            cosine_reg0 <= 36'sb101000101101001011100111011001100101;
            sine_reg0   <= 36'sb10101111100001100011111100100100110;
        end
        6223: begin
            cosine_reg0 <= 36'sb101000101100101001001010001001001110;
            sine_reg0   <= 36'sb10101111011100111111001011000000111;
        end
        6224: begin
            cosine_reg0 <= 36'sb101000101100000110101101110010010111;
            sine_reg0   <= 36'sb10101111011000011010010010101100000;
        end
        6225: begin
            cosine_reg0 <= 36'sb101000101011100100010010010101000000;
            sine_reg0   <= 36'sb10101111010011110101010011100110100;
        end
        6226: begin
            cosine_reg0 <= 36'sb101000101011000001110111110001001101;
            sine_reg0   <= 36'sb10101111001111010000001101110000011;
        end
        6227: begin
            cosine_reg0 <= 36'sb101000101010011111011110000110111101;
            sine_reg0   <= 36'sb10101111001010101011000001001001111;
        end
        6228: begin
            cosine_reg0 <= 36'sb101000101001111101000101010110010010;
            sine_reg0   <= 36'sb10101111000110000101101101110011001;
        end
        6229: begin
            cosine_reg0 <= 36'sb101000101001011010101101011111001110;
            sine_reg0   <= 36'sb10101111000001100000010011101100100;
        end
        6230: begin
            cosine_reg0 <= 36'sb101000101000111000010110100001110001;
            sine_reg0   <= 36'sb10101110111100111010110010110101111;
        end
        6231: begin
            cosine_reg0 <= 36'sb101000101000010110000000011101111110;
            sine_reg0   <= 36'sb10101110111000010101001011001111101;
        end
        6232: begin
            cosine_reg0 <= 36'sb101000100111110011101011010011110101;
            sine_reg0   <= 36'sb10101110110011101111011100111001111;
        end
        6233: begin
            cosine_reg0 <= 36'sb101000100111010001010111000011010111;
            sine_reg0   <= 36'sb10101110101111001001100111110100110;
        end
        6234: begin
            cosine_reg0 <= 36'sb101000100110101111000011101100100111;
            sine_reg0   <= 36'sb10101110101010100011101100000000100;
        end
        6235: begin
            cosine_reg0 <= 36'sb101000100110001100110001001111100101;
            sine_reg0   <= 36'sb10101110100101111101101001011101011;
        end
        6236: begin
            cosine_reg0 <= 36'sb101000100101101010011111101100010010;
            sine_reg0   <= 36'sb10101110100001010111100000001011011;
        end
        6237: begin
            cosine_reg0 <= 36'sb101000100101001000001111000010110001;
            sine_reg0   <= 36'sb10101110011100110001010000001010110;
        end
        6238: begin
            cosine_reg0 <= 36'sb101000100100100101111111010011000010;
            sine_reg0   <= 36'sb10101110011000001010111001011011110;
        end
        6239: begin
            cosine_reg0 <= 36'sb101000100100000011110000011101000110;
            sine_reg0   <= 36'sb10101110010011100100011011111110100;
        end
        6240: begin
            cosine_reg0 <= 36'sb101000100011100001100010100001000000;
            sine_reg0   <= 36'sb10101110001110111101110111110011001;
        end
        6241: begin
            cosine_reg0 <= 36'sb101000100010111111010101011110110000;
            sine_reg0   <= 36'sb10101110001010010111001100111001110;
        end
        6242: begin
            cosine_reg0 <= 36'sb101000100010011101001001010110010111;
            sine_reg0   <= 36'sb10101110000101110000011011010010110;
        end
        6243: begin
            cosine_reg0 <= 36'sb101000100001111010111110000111110111;
            sine_reg0   <= 36'sb10101110000001001001100010111110010;
        end
        6244: begin
            cosine_reg0 <= 36'sb101000100001011000110011110011010010;
            sine_reg0   <= 36'sb10101101111100100010100011111100010;
        end
        6245: begin
            cosine_reg0 <= 36'sb101000100000110110101010011000101000;
            sine_reg0   <= 36'sb10101101110111111011011110001101001;
        end
        6246: begin
            cosine_reg0 <= 36'sb101000100000010100100001110111111011;
            sine_reg0   <= 36'sb10101101110011010100010001110001000;
        end
        6247: begin
            cosine_reg0 <= 36'sb101000011111110010011010010001001100;
            sine_reg0   <= 36'sb10101101101110101100111110101000000;
        end
        6248: begin
            cosine_reg0 <= 36'sb101000011111010000010011100100011101;
            sine_reg0   <= 36'sb10101101101010000101100100110010011;
        end
        6249: begin
            cosine_reg0 <= 36'sb101000011110101110001101110001101110;
            sine_reg0   <= 36'sb10101101100101011110000100010000010;
        end
        6250: begin
            cosine_reg0 <= 36'sb101000011110001100001000111001000010;
            sine_reg0   <= 36'sb10101101100000110110011101000001111;
        end
        6251: begin
            cosine_reg0 <= 36'sb101000011101101010000100111010011000;
            sine_reg0   <= 36'sb10101101011100001110101111000111010;
        end
        6252: begin
            cosine_reg0 <= 36'sb101000011101001000000001110101110100;
            sine_reg0   <= 36'sb10101101010111100110111010100000110;
        end
        6253: begin
            cosine_reg0 <= 36'sb101000011100100101111111101011010110;
            sine_reg0   <= 36'sb10101101010010111110111111001110100;
        end
        6254: begin
            cosine_reg0 <= 36'sb101000011100000011111110011010111111;
            sine_reg0   <= 36'sb10101101001110010110111101010000101;
        end
        6255: begin
            cosine_reg0 <= 36'sb101000011011100001111110000100110001;
            sine_reg0   <= 36'sb10101101001001101110110100100111011;
        end
        6256: begin
            cosine_reg0 <= 36'sb101000011010111111111110101000101101;
            sine_reg0   <= 36'sb10101101000101000110100101010010111;
        end
        6257: begin
            cosine_reg0 <= 36'sb101000011010011110000000000110110100;
            sine_reg0   <= 36'sb10101101000000011110001111010011010;
        end
        6258: begin
            cosine_reg0 <= 36'sb101000011001111100000010011111001000;
            sine_reg0   <= 36'sb10101100111011110101110010101000110;
        end
        6259: begin
            cosine_reg0 <= 36'sb101000011001011010000101110001101010;
            sine_reg0   <= 36'sb10101100110111001101001111010011101;
        end
        6260: begin
            cosine_reg0 <= 36'sb101000011000111000001001111110011011;
            sine_reg0   <= 36'sb10101100110010100100100101010100000;
        end
        6261: begin
            cosine_reg0 <= 36'sb101000011000010110001111000101011100;
            sine_reg0   <= 36'sb10101100101101111011110100101010000;
        end
        6262: begin
            cosine_reg0 <= 36'sb101000010111110100010101000110101111;
            sine_reg0   <= 36'sb10101100101001010010111101010101110;
        end
        6263: begin
            cosine_reg0 <= 36'sb101000010111010010011100000010010110;
            sine_reg0   <= 36'sb10101100100100101001111111010111101;
        end
        6264: begin
            cosine_reg0 <= 36'sb101000010110110000100011111000010001;
            sine_reg0   <= 36'sb10101100100000000000111010101111101;
        end
        6265: begin
            cosine_reg0 <= 36'sb101000010110001110101100101000100010;
            sine_reg0   <= 36'sb10101100011011010111101111011110000;
        end
        6266: begin
            cosine_reg0 <= 36'sb101000010101101100110110010011001001;
            sine_reg0   <= 36'sb10101100010110101110011101100011000;
        end
        6267: begin
            cosine_reg0 <= 36'sb101000010101001011000000111000001010;
            sine_reg0   <= 36'sb10101100010010000101000100111110101;
        end
        6268: begin
            cosine_reg0 <= 36'sb101000010100101001001100010111100100;
            sine_reg0   <= 36'sb10101100001101011011100101110001010;
        end
        6269: begin
            cosine_reg0 <= 36'sb101000010100000111011000110001011000;
            sine_reg0   <= 36'sb10101100001000110001111111111011000;
        end
        6270: begin
            cosine_reg0 <= 36'sb101000010011100101100110000101101010;
            sine_reg0   <= 36'sb10101100000100001000010011011011111;
        end
        6271: begin
            cosine_reg0 <= 36'sb101000010011000011110100010100011000;
            sine_reg0   <= 36'sb10101011111111011110100000010100010;
        end
        6272: begin
            cosine_reg0 <= 36'sb101000010010100010000011011101100110;
            sine_reg0   <= 36'sb10101011111010110100100110100100011;
        end
        6273: begin
            cosine_reg0 <= 36'sb101000010010000000010011100001010100;
            sine_reg0   <= 36'sb10101011110110001010100110001100001;
        end
        6274: begin
            cosine_reg0 <= 36'sb101000010001011110100100011111100011;
            sine_reg0   <= 36'sb10101011110001100000011111001100000;
        end
        6275: begin
            cosine_reg0 <= 36'sb101000010000111100110110011000010110;
            sine_reg0   <= 36'sb10101011101100110110010001100100000;
        end
        6276: begin
            cosine_reg0 <= 36'sb101000010000011011001001001011101100;
            sine_reg0   <= 36'sb10101011101000001011111101010100010;
        end
        6277: begin
            cosine_reg0 <= 36'sb101000001111111001011100111001101000;
            sine_reg0   <= 36'sb10101011100011100001100010011101001;
        end
        6278: begin
            cosine_reg0 <= 36'sb101000001111010111110001100010001010;
            sine_reg0   <= 36'sb10101011011110110111000000111110110;
        end
        6279: begin
            cosine_reg0 <= 36'sb101000001110110110000111000101010100;
            sine_reg0   <= 36'sb10101011011010001100011000111001001;
        end
        6280: begin
            cosine_reg0 <= 36'sb101000001110010100011101100011001000;
            sine_reg0   <= 36'sb10101011010101100001101010001100101;
        end
        6281: begin
            cosine_reg0 <= 36'sb101000001101110010110100111011100110;
            sine_reg0   <= 36'sb10101011010000110110110100111001011;
        end
        6282: begin
            cosine_reg0 <= 36'sb101000001101010001001101001110110001;
            sine_reg0   <= 36'sb10101011001100001011111000111111101;
        end
        6283: begin
            cosine_reg0 <= 36'sb101000001100101111100110011100101000;
            sine_reg0   <= 36'sb10101011000111100000110110011111011;
        end
        6284: begin
            cosine_reg0 <= 36'sb101000001100001110000000100101001110;
            sine_reg0   <= 36'sb10101011000010110101101101011000111;
        end
        6285: begin
            cosine_reg0 <= 36'sb101000001011101100011011101000100011;
            sine_reg0   <= 36'sb10101010111110001010011101101100100;
        end
        6286: begin
            cosine_reg0 <= 36'sb101000001011001010110111100110101010;
            sine_reg0   <= 36'sb10101010111001011111000111011010001;
        end
        6287: begin
            cosine_reg0 <= 36'sb101000001010101001010100011111100011;
            sine_reg0   <= 36'sb10101010110100110011101010100010001;
        end
        6288: begin
            cosine_reg0 <= 36'sb101000001010000111110010010011010000;
            sine_reg0   <= 36'sb10101010110000001000000111000100101;
        end
        6289: begin
            cosine_reg0 <= 36'sb101000001001100110010001000001110010;
            sine_reg0   <= 36'sb10101010101011011100011101000001111;
        end
        6290: begin
            cosine_reg0 <= 36'sb101000001001000100110000101011001010;
            sine_reg0   <= 36'sb10101010100110110000101100011001111;
        end
        6291: begin
            cosine_reg0 <= 36'sb101000001000100011010001001111011001;
            sine_reg0   <= 36'sb10101010100010000100110101001101000;
        end
        6292: begin
            cosine_reg0 <= 36'sb101000001000000001110010101110100001;
            sine_reg0   <= 36'sb10101010011101011000110111011011011;
        end
        6293: begin
            cosine_reg0 <= 36'sb101000000111100000010101001000100100;
            sine_reg0   <= 36'sb10101010011000101100110011000101001;
        end
        6294: begin
            cosine_reg0 <= 36'sb101000000110111110111000011101100010;
            sine_reg0   <= 36'sb10101010010100000000101000001010011;
        end
        6295: begin
            cosine_reg0 <= 36'sb101000000110011101011100101101011100;
            sine_reg0   <= 36'sb10101010001111010100010110101011100;
        end
        6296: begin
            cosine_reg0 <= 36'sb101000000101111100000001111000010101;
            sine_reg0   <= 36'sb10101010001010100111111110101000101;
        end
        6297: begin
            cosine_reg0 <= 36'sb101000000101011010100111111110001100;
            sine_reg0   <= 36'sb10101010000101111011100000000001110;
        end
        6298: begin
            cosine_reg0 <= 36'sb101000000100111001001110111111000101;
            sine_reg0   <= 36'sb10101010000001001110111010110111010;
        end
        6299: begin
            cosine_reg0 <= 36'sb101000000100010111110110111010111111;
            sine_reg0   <= 36'sb10101001111100100010001111001001010;
        end
        6300: begin
            cosine_reg0 <= 36'sb101000000011110110011111110001111100;
            sine_reg0   <= 36'sb10101001110111110101011100111000000;
        end
        6301: begin
            cosine_reg0 <= 36'sb101000000011010101001001100011111110;
            sine_reg0   <= 36'sb10101001110011001000100100000011100;
        end
        6302: begin
            cosine_reg0 <= 36'sb101000000010110011110100010001000110;
            sine_reg0   <= 36'sb10101001101110011011100100101100000;
        end
        6303: begin
            cosine_reg0 <= 36'sb101000000010010010011111111001010100;
            sine_reg0   <= 36'sb10101001101001101110011110110001111;
        end
        6304: begin
            cosine_reg0 <= 36'sb101000000001110001001100011100101011;
            sine_reg0   <= 36'sb10101001100101000001010010010101000;
        end
        6305: begin
            cosine_reg0 <= 36'sb101000000001001111111001111011001011;
            sine_reg0   <= 36'sb10101001100000010011111111010101110;
        end
        6306: begin
            cosine_reg0 <= 36'sb101000000000101110101000010100110110;
            sine_reg0   <= 36'sb10101001011011100110100101110100011;
        end
        6307: begin
            cosine_reg0 <= 36'sb101000000000001101010111101001101110;
            sine_reg0   <= 36'sb10101001010110111001000101110000110;
        end
        6308: begin
            cosine_reg0 <= 36'sb100111111111101100000111111001110011;
            sine_reg0   <= 36'sb10101001010010001011011111001011011;
        end
        6309: begin
            cosine_reg0 <= 36'sb100111111111001010111001000101000110;
            sine_reg0   <= 36'sb10101001001101011101110010000100011;
        end
        6310: begin
            cosine_reg0 <= 36'sb100111111110101001101011001011101001;
            sine_reg0   <= 36'sb10101001001000101111111110011011110;
        end
        6311: begin
            cosine_reg0 <= 36'sb100111111110001000011110001101011110;
            sine_reg0   <= 36'sb10101001000100000010000100010001110;
        end
        6312: begin
            cosine_reg0 <= 36'sb100111111101100111010010001010100101;
            sine_reg0   <= 36'sb10101000111111010100000011100110110;
        end
        6313: begin
            cosine_reg0 <= 36'sb100111111101000110000111000011000000;
            sine_reg0   <= 36'sb10101000111010100101111100011010101;
        end
        6314: begin
            cosine_reg0 <= 36'sb100111111100100100111100110110110000;
            sine_reg0   <= 36'sb10101000110101110111101110101101111;
        end
        6315: begin
            cosine_reg0 <= 36'sb100111111100000011110011100101110111;
            sine_reg0   <= 36'sb10101000110001001001011010100000100;
        end
        6316: begin
            cosine_reg0 <= 36'sb100111111011100010101011010000010101;
            sine_reg0   <= 36'sb10101000101100011010111111110010101;
        end
        6317: begin
            cosine_reg0 <= 36'sb100111111011000001100011110110001100;
            sine_reg0   <= 36'sb10101000100111101100011110100100100;
        end
        6318: begin
            cosine_reg0 <= 36'sb100111111010100000011101010111011101;
            sine_reg0   <= 36'sb10101000100010111101110110110110011;
        end
        6319: begin
            cosine_reg0 <= 36'sb100111111001111111010111110100001010;
            sine_reg0   <= 36'sb10101000011110001111001000101000011;
        end
        6320: begin
            cosine_reg0 <= 36'sb100111111001011110010011001100010011;
            sine_reg0   <= 36'sb10101000011001100000010011111010110;
        end
        6321: begin
            cosine_reg0 <= 36'sb100111111000111101001111011111111011;
            sine_reg0   <= 36'sb10101000010100110001011000101101100;
        end
        6322: begin
            cosine_reg0 <= 36'sb100111111000011100001100101111000010;
            sine_reg0   <= 36'sb10101000010000000010010111000001000;
        end
        6323: begin
            cosine_reg0 <= 36'sb100111110111111011001010111001101001;
            sine_reg0   <= 36'sb10101000001011010011001110110101011;
        end
        6324: begin
            cosine_reg0 <= 36'sb100111110111011010001001111111110010;
            sine_reg0   <= 36'sb10101000000110100100000000001010110;
        end
        6325: begin
            cosine_reg0 <= 36'sb100111110110111001001010000001011111;
            sine_reg0   <= 36'sb10101000000001110100101011000001011;
        end
        6326: begin
            cosine_reg0 <= 36'sb100111110110011000001010111110110000;
            sine_reg0   <= 36'sb10100111111101000101001111011001011;
        end
        6327: begin
            cosine_reg0 <= 36'sb100111110101110111001100110111100110;
            sine_reg0   <= 36'sb10100111111000010101101101010011000;
        end
        6328: begin
            cosine_reg0 <= 36'sb100111110101010110001111101100000011;
            sine_reg0   <= 36'sb10100111110011100110000100101110011;
        end
        6329: begin
            cosine_reg0 <= 36'sb100111110100110101010011011100001001;
            sine_reg0   <= 36'sb10100111101110110110010101101011101;
        end
        6330: begin
            cosine_reg0 <= 36'sb100111110100010100011000000111111000;
            sine_reg0   <= 36'sb10100111101010000110100000001011001;
        end
        6331: begin
            cosine_reg0 <= 36'sb100111110011110011011101101111010010;
            sine_reg0   <= 36'sb10100111100101010110100100001100111;
        end
        6332: begin
            cosine_reg0 <= 36'sb100111110011010010100100010010011000;
            sine_reg0   <= 36'sb10100111100000100110100001110001001;
        end
        6333: begin
            cosine_reg0 <= 36'sb100111110010110001101011110001001011;
            sine_reg0   <= 36'sb10100111011011110110011000111000001;
        end
        6334: begin
            cosine_reg0 <= 36'sb100111110010010000110100001011101101;
            sine_reg0   <= 36'sb10100111010111000110001001100010000;
        end
        6335: begin
            cosine_reg0 <= 36'sb100111110001101111111101100001111110;
            sine_reg0   <= 36'sb10100111010010010101110011101110111;
        end
        6336: begin
            cosine_reg0 <= 36'sb100111110001001111000111110100000001;
            sine_reg0   <= 36'sb10100111001101100101010111011111000;
        end
        6337: begin
            cosine_reg0 <= 36'sb100111110000101110010011000001110110;
            sine_reg0   <= 36'sb10100111001000110100110100110010101;
        end
        6338: begin
            cosine_reg0 <= 36'sb100111110000001101011111001011011110;
            sine_reg0   <= 36'sb10100111000100000100001011101001110;
        end
        6339: begin
            cosine_reg0 <= 36'sb100111101111101100101100010000111100;
            sine_reg0   <= 36'sb10100110111111010011011100000100110;
        end
        6340: begin
            cosine_reg0 <= 36'sb100111101111001011111010010010010000;
            sine_reg0   <= 36'sb10100110111010100010100110000011101;
        end
        6341: begin
            cosine_reg0 <= 36'sb100111101110101011001001001111011011;
            sine_reg0   <= 36'sb10100110110101110001101001100110110;
        end
        6342: begin
            cosine_reg0 <= 36'sb100111101110001010011001001000011110;
            sine_reg0   <= 36'sb10100110110001000000100110101110001;
        end
        6343: begin
            cosine_reg0 <= 36'sb100111101101101001101001111101011100;
            sine_reg0   <= 36'sb10100110101100001111011101011010000;
        end
        6344: begin
            cosine_reg0 <= 36'sb100111101101001000111011101110010101;
            sine_reg0   <= 36'sb10100110100111011110001101101010110;
        end
        6345: begin
            cosine_reg0 <= 36'sb100111101100101000001110011011001010;
            sine_reg0   <= 36'sb10100110100010101100110111100000010;
        end
        6346: begin
            cosine_reg0 <= 36'sb100111101100000111100010000011111101;
            sine_reg0   <= 36'sb10100110011101111011011010111010111;
        end
        6347: begin
            cosine_reg0 <= 36'sb100111101011100110110110101000101111;
            sine_reg0   <= 36'sb10100110011001001001110111111010101;
        end
        6348: begin
            cosine_reg0 <= 36'sb100111101011000110001100001001100010;
            sine_reg0   <= 36'sb10100110010100011000001110100000000;
        end
        6349: begin
            cosine_reg0 <= 36'sb100111101010100101100010100110010101;
            sine_reg0   <= 36'sb10100110001111100110011110101010111;
        end
        6350: begin
            cosine_reg0 <= 36'sb100111101010000100111001111111001100;
            sine_reg0   <= 36'sb10100110001010110100101000011011101;
        end
        6351: begin
            cosine_reg0 <= 36'sb100111101001100100010010010100000111;
            sine_reg0   <= 36'sb10100110000110000010101011110010011;
        end
        6352: begin
            cosine_reg0 <= 36'sb100111101001000011101011100101000110;
            sine_reg0   <= 36'sb10100110000001010000101000101111010;
        end
        6353: begin
            cosine_reg0 <= 36'sb100111101000100011000101110010001101;
            sine_reg0   <= 36'sb10100101111100011110011111010010101;
        end
        6354: begin
            cosine_reg0 <= 36'sb100111101000000010100000111011011011;
            sine_reg0   <= 36'sb10100101110111101100001111011100011;
        end
        6355: begin
            cosine_reg0 <= 36'sb100111100111100001111101000000110010;
            sine_reg0   <= 36'sb10100101110010111001111001001101000;
        end
        6356: begin
            cosine_reg0 <= 36'sb100111100111000001011010000010010100;
            sine_reg0   <= 36'sb10100101101110000111011100100100011;
        end
        6357: begin
            cosine_reg0 <= 36'sb100111100110100000111000000000000001;
            sine_reg0   <= 36'sb10100101101001010100111001100011000;
        end
        6358: begin
            cosine_reg0 <= 36'sb100111100110000000010110111001111011;
            sine_reg0   <= 36'sb10100101100100100010010000001000111;
        end
        6359: begin
            cosine_reg0 <= 36'sb100111100101011111110110110000000011;
            sine_reg0   <= 36'sb10100101011111101111100000010110001;
        end
        6360: begin
            cosine_reg0 <= 36'sb100111100100111111010111100010011010;
            sine_reg0   <= 36'sb10100101011010111100101010001011001;
        end
        6361: begin
            cosine_reg0 <= 36'sb100111100100011110111001010001000010;
            sine_reg0   <= 36'sb10100101010110001001101101101000000;
        end
        6362: begin
            cosine_reg0 <= 36'sb100111100011111110011011111011111100;
            sine_reg0   <= 36'sb10100101010001010110101010101100110;
        end
        6363: begin
            cosine_reg0 <= 36'sb100111100011011101111111100011001000;
            sine_reg0   <= 36'sb10100101001100100011100001011001111;
        end
        6364: begin
            cosine_reg0 <= 36'sb100111100010111101100100000110101010;
            sine_reg0   <= 36'sb10100101000111110000010001101111011;
        end
        6365: begin
            cosine_reg0 <= 36'sb100111100010011101001001100110100000;
            sine_reg0   <= 36'sb10100101000010111100111011101101011;
        end
        6366: begin
            cosine_reg0 <= 36'sb100111100001111100110000000010101110;
            sine_reg0   <= 36'sb10100100111110001001011111010100001;
        end
        6367: begin
            cosine_reg0 <= 36'sb100111100001011100010111011011010011;
            sine_reg0   <= 36'sb10100100111001010101111100100011111;
        end
        6368: begin
            cosine_reg0 <= 36'sb100111100000111011111111110000010010;
            sine_reg0   <= 36'sb10100100110100100010010011011100110;
        end
        6369: begin
            cosine_reg0 <= 36'sb100111100000011011101001000001101100;
            sine_reg0   <= 36'sb10100100101111101110100011111111000;
        end
        6370: begin
            cosine_reg0 <= 36'sb100111011111111011010011001111100001;
            sine_reg0   <= 36'sb10100100101010111010101110001010101;
        end
        6371: begin
            cosine_reg0 <= 36'sb100111011111011010111110011001110011;
            sine_reg0   <= 36'sb10100100100110000110110010000000001;
        end
        6372: begin
            cosine_reg0 <= 36'sb100111011110111010101010100000100100;
            sine_reg0   <= 36'sb10100100100001010010101111011111011;
        end
        6373: begin
            cosine_reg0 <= 36'sb100111011110011010010111100011110100;
            sine_reg0   <= 36'sb10100100011100011110100110101000110;
        end
        6374: begin
            cosine_reg0 <= 36'sb100111011101111010000101100011100101;
            sine_reg0   <= 36'sb10100100010111101010010111011100010;
        end
        6375: begin
            cosine_reg0 <= 36'sb100111011101011001110100011111111000;
            sine_reg0   <= 36'sb10100100010010110110000001111010010;
        end
        6376: begin
            cosine_reg0 <= 36'sb100111011100111001100100011000101111;
            sine_reg0   <= 36'sb10100100001110000001100110000011000;
        end
        6377: begin
            cosine_reg0 <= 36'sb100111011100011001010101001110001010;
            sine_reg0   <= 36'sb10100100001001001101000011110110011;
        end
        6378: begin
            cosine_reg0 <= 36'sb100111011011111001000111000000001010;
            sine_reg0   <= 36'sb10100100000100011000011011010100111;
        end
        6379: begin
            cosine_reg0 <= 36'sb100111011011011000111001101110110010;
            sine_reg0   <= 36'sb10100011111111100011101100011110011;
        end
        6380: begin
            cosine_reg0 <= 36'sb100111011010111000101101011010000010;
            sine_reg0   <= 36'sb10100011111010101110110111010011011;
        end
        6381: begin
            cosine_reg0 <= 36'sb100111011010011000100010000001111011;
            sine_reg0   <= 36'sb10100011110101111001111011110100000;
        end
        6382: begin
            cosine_reg0 <= 36'sb100111011001111000010111100110100000;
            sine_reg0   <= 36'sb10100011110001000100111010000000010;
        end
        6383: begin
            cosine_reg0 <= 36'sb100111011001011000001110000111110000;
            sine_reg0   <= 36'sb10100011101100001111110001111000011;
        end
        6384: begin
            cosine_reg0 <= 36'sb100111011000111000000101100101101101;
            sine_reg0   <= 36'sb10100011100111011010100011011100101;
        end
        6385: begin
            cosine_reg0 <= 36'sb100111011000010111111110000000011001;
            sine_reg0   <= 36'sb10100011100010100101001110101101010;
        end
        6386: begin
            cosine_reg0 <= 36'sb100111010111110111110111010111110101;
            sine_reg0   <= 36'sb10100011011101101111110011101010011;
        end
        6387: begin
            cosine_reg0 <= 36'sb100111010111010111110001101100000001;
            sine_reg0   <= 36'sb10100011011000111010010010010100001;
        end
        6388: begin
            cosine_reg0 <= 36'sb100111010110110111101100111101000000;
            sine_reg0   <= 36'sb10100011010100000100101010101010101;
        end
        6389: begin
            cosine_reg0 <= 36'sb100111010110010111101001001010110010;
            sine_reg0   <= 36'sb10100011001111001110111100101110010;
        end
        6390: begin
            cosine_reg0 <= 36'sb100111010101110111100110010101011001;
            sine_reg0   <= 36'sb10100011001010011001001000011111001;
        end
        6391: begin
            cosine_reg0 <= 36'sb100111010101010111100100011100110101;
            sine_reg0   <= 36'sb10100011000101100011001101111101011;
        end
        6392: begin
            cosine_reg0 <= 36'sb100111010100110111100011100001001001;
            sine_reg0   <= 36'sb10100011000000101101001101001001010;
        end
        6393: begin
            cosine_reg0 <= 36'sb100111010100010111100011100010010101;
            sine_reg0   <= 36'sb10100010111011110111000110000010111;
        end
        6394: begin
            cosine_reg0 <= 36'sb100111010011110111100100100000011011;
            sine_reg0   <= 36'sb10100010110111000000111000101010100;
        end
        6395: begin
            cosine_reg0 <= 36'sb100111010011010111100110011011011100;
            sine_reg0   <= 36'sb10100010110010001010100101000000011;
        end
        6396: begin
            cosine_reg0 <= 36'sb100111010010110111101001010011011000;
            sine_reg0   <= 36'sb10100010101101010100001011000100100;
        end
        6397: begin
            cosine_reg0 <= 36'sb100111010010010111101101001000010010;
            sine_reg0   <= 36'sb10100010101000011101101010110111001;
        end
        6398: begin
            cosine_reg0 <= 36'sb100111010001110111110001111010001010;
            sine_reg0   <= 36'sb10100010100011100111000100011000100;
        end
        6399: begin
            cosine_reg0 <= 36'sb100111010001010111110111101001000010;
            sine_reg0   <= 36'sb10100010011110110000010111101000111;
        end
        6400: begin
            cosine_reg0 <= 36'sb100111010000110111111110010100111100;
            sine_reg0   <= 36'sb10100010011001111001100100101000010;
        end
        6401: begin
            cosine_reg0 <= 36'sb100111010000011000000101111101110111;
            sine_reg0   <= 36'sb10100010010101000010101011010110111;
        end
        6402: begin
            cosine_reg0 <= 36'sb100111001111111000001110100011110110;
            sine_reg0   <= 36'sb10100010010000001011101011110101000;
        end
        6403: begin
            cosine_reg0 <= 36'sb100111001111011000011000000110111001;
            sine_reg0   <= 36'sb10100010001011010100100110000010111;
        end
        6404: begin
            cosine_reg0 <= 36'sb100111001110111000100010100111000010;
            sine_reg0   <= 36'sb10100010000110011101011010000000100;
        end
        6405: begin
            cosine_reg0 <= 36'sb100111001110011000101110000100010011;
            sine_reg0   <= 36'sb10100010000001100110000111101110001;
        end
        6406: begin
            cosine_reg0 <= 36'sb100111001101111000111010011110101011;
            sine_reg0   <= 36'sb10100001111100101110101111001100000;
        end
        6407: begin
            cosine_reg0 <= 36'sb100111001101011001000111110110001110;
            sine_reg0   <= 36'sb10100001110111110111010000011010011;
        end
        6408: begin
            cosine_reg0 <= 36'sb100111001100111001010110001010111011;
            sine_reg0   <= 36'sb10100001110010111111101011011001010;
        end
        6409: begin
            cosine_reg0 <= 36'sb100111001100011001100101011100110100;
            sine_reg0   <= 36'sb10100001101110001000000000001000111;
        end
        6410: begin
            cosine_reg0 <= 36'sb100111001011111001110101101011111010;
            sine_reg0   <= 36'sb10100001101001010000001110101001101;
        end
        6411: begin
            cosine_reg0 <= 36'sb100111001011011010000110111000001111;
            sine_reg0   <= 36'sb10100001100100011000010110111011011;
        end
        6412: begin
            cosine_reg0 <= 36'sb100111001010111010011001000001110100;
            sine_reg0   <= 36'sb10100001011111100000011000111110100;
        end
        6413: begin
            cosine_reg0 <= 36'sb100111001010011010101100001000101001;
            sine_reg0   <= 36'sb10100001011010101000010100110011010;
        end
        6414: begin
            cosine_reg0 <= 36'sb100111001001111011000000001100110001;
            sine_reg0   <= 36'sb10100001010101110000001010011001101;
        end
        6415: begin
            cosine_reg0 <= 36'sb100111001001011011010101001110001100;
            sine_reg0   <= 36'sb10100001010000110111111001110010000;
        end
        6416: begin
            cosine_reg0 <= 36'sb100111001000111011101011001100111011;
            sine_reg0   <= 36'sb10100001001011111111100010111100011;
        end
        6417: begin
            cosine_reg0 <= 36'sb100111001000011100000010001001000000;
            sine_reg0   <= 36'sb10100001000111000111000101111001001;
        end
        6418: begin
            cosine_reg0 <= 36'sb100111000111111100011010000010011101;
            sine_reg0   <= 36'sb10100001000010001110100010101000010;
        end
        6419: begin
            cosine_reg0 <= 36'sb100111000111011100110010111001010001;
            sine_reg0   <= 36'sb10100000111101010101111001001010001;
        end
        6420: begin
            cosine_reg0 <= 36'sb100111000110111101001100101101011111;
            sine_reg0   <= 36'sb10100000111000011101001001011110110;
        end
        6421: begin
            cosine_reg0 <= 36'sb100111000110011101100111011111001000;
            sine_reg0   <= 36'sb10100000110011100100010011100110100;
        end
        6422: begin
            cosine_reg0 <= 36'sb100111000101111110000011001110001101;
            sine_reg0   <= 36'sb10100000101110101011010111100001100;
        end
        6423: begin
            cosine_reg0 <= 36'sb100111000101011110011111111010101111;
            sine_reg0   <= 36'sb10100000101001110010010101001111111;
        end
        6424: begin
            cosine_reg0 <= 36'sb100111000100111110111101100100101111;
            sine_reg0   <= 36'sb10100000100100111001001100110001111;
        end
        6425: begin
            cosine_reg0 <= 36'sb100111000100011111011100001100001110;
            sine_reg0   <= 36'sb10100000011111111111111110000111101;
        end
        6426: begin
            cosine_reg0 <= 36'sb100111000011111111111011110001001111;
            sine_reg0   <= 36'sb10100000011011000110101001010001011;
        end
        6427: begin
            cosine_reg0 <= 36'sb100111000011100000011100010011110001;
            sine_reg0   <= 36'sb10100000010110001101001110001111010;
        end
        6428: begin
            cosine_reg0 <= 36'sb100111000011000000111101110011110111;
            sine_reg0   <= 36'sb10100000010001010011101101000001101;
        end
        6429: begin
            cosine_reg0 <= 36'sb100111000010100001100000010001100001;
            sine_reg0   <= 36'sb10100000001100011010000101101000011;
        end
        6430: begin
            cosine_reg0 <= 36'sb100111000010000010000011101100110000;
            sine_reg0   <= 36'sb10100000000111100000011000000100000;
        end
        6431: begin
            cosine_reg0 <= 36'sb100111000001100010101000000101100110;
            sine_reg0   <= 36'sb10100000000010100110100100010100100;
        end
        6432: begin
            cosine_reg0 <= 36'sb100111000001000011001101011100000101;
            sine_reg0   <= 36'sb10011111111101101100101010011010001;
        end
        6433: begin
            cosine_reg0 <= 36'sb100111000000100011110011110000001101;
            sine_reg0   <= 36'sb10011111111000110010101010010101000;
        end
        6434: begin
            cosine_reg0 <= 36'sb100111000000000100011011000001111111;
            sine_reg0   <= 36'sb10011111110011111000100100000101011;
        end
        6435: begin
            cosine_reg0 <= 36'sb100110111111100101000011010001011101;
            sine_reg0   <= 36'sb10011111101110111110010111101011100;
        end
        6436: begin
            cosine_reg0 <= 36'sb100110111111000101101100011110100111;
            sine_reg0   <= 36'sb10011111101010000100000101000111100;
        end
        6437: begin
            cosine_reg0 <= 36'sb100110111110100110010110101001100000;
            sine_reg0   <= 36'sb10011111100101001001101100011001100;
        end
        6438: begin
            cosine_reg0 <= 36'sb100110111110000111000001110010001000;
            sine_reg0   <= 36'sb10011111100000001111001101100001110;
        end
        6439: begin
            cosine_reg0 <= 36'sb100110111101100111101101111000100001;
            sine_reg0   <= 36'sb10011111011011010100101000100000100;
        end
        6440: begin
            cosine_reg0 <= 36'sb100110111101001000011010111100101011;
            sine_reg0   <= 36'sb10011111010110011001111101010101111;
        end
        6441: begin
            cosine_reg0 <= 36'sb100110111100101001001000111110101000;
            sine_reg0   <= 36'sb10011111010001011111001100000010000;
        end
        6442: begin
            cosine_reg0 <= 36'sb100110111100001001110111111110011001;
            sine_reg0   <= 36'sb10011111001100100100010100100101010;
        end
        6443: begin
            cosine_reg0 <= 36'sb100110111011101010100111111100000000;
            sine_reg0   <= 36'sb10011111000111101001010110111111101;
        end
        6444: begin
            cosine_reg0 <= 36'sb100110111011001011011000110111011101;
            sine_reg0   <= 36'sb10011111000010101110010011010001011;
        end
        6445: begin
            cosine_reg0 <= 36'sb100110111010101100001010110000110010;
            sine_reg0   <= 36'sb10011110111101110011001001011010110;
        end
        6446: begin
            cosine_reg0 <= 36'sb100110111010001100111101101000000000;
            sine_reg0   <= 36'sb10011110111000110111111001011011110;
        end
        6447: begin
            cosine_reg0 <= 36'sb100110111001101101110001011101001000;
            sine_reg0   <= 36'sb10011110110011111100100011010100111;
        end
        6448: begin
            cosine_reg0 <= 36'sb100110111001001110100110010000001100;
            sine_reg0   <= 36'sb10011110101111000001000111000110001;
        end
        6449: begin
            cosine_reg0 <= 36'sb100110111000101111011100000001001100;
            sine_reg0   <= 36'sb10011110101010000101100100101111101;
        end
        6450: begin
            cosine_reg0 <= 36'sb100110111000010000010010110000001001;
            sine_reg0   <= 36'sb10011110100101001001111100010001110;
        end
        6451: begin
            cosine_reg0 <= 36'sb100110110111110001001010011101000110;
            sine_reg0   <= 36'sb10011110100000001110001101101100100;
        end
        6452: begin
            cosine_reg0 <= 36'sb100110110111010010000011001000000011;
            sine_reg0   <= 36'sb10011110011011010010011001000000010;
        end
        6453: begin
            cosine_reg0 <= 36'sb100110110110110010111100110001000001;
            sine_reg0   <= 36'sb10011110010110010110011110001101000;
        end
        6454: begin
            cosine_reg0 <= 36'sb100110110110010011110111011000000010;
            sine_reg0   <= 36'sb10011110010001011010011101010011001;
        end
        6455: begin
            cosine_reg0 <= 36'sb100110110101110100110010111101000110;
            sine_reg0   <= 36'sb10011110001100011110010110010010110;
        end
        6456: begin
            cosine_reg0 <= 36'sb100110110101010101101111100000001111;
            sine_reg0   <= 36'sb10011110000111100010001001001100000;
        end
        6457: begin
            cosine_reg0 <= 36'sb100110110100110110101101000001011111;
            sine_reg0   <= 36'sb10011110000010100101110101111111001;
        end
        6458: begin
            cosine_reg0 <= 36'sb100110110100010111101011100000110110;
            sine_reg0   <= 36'sb10011101111101101001011100101100010;
        end
        6459: begin
            cosine_reg0 <= 36'sb100110110011111000101010111110010101;
            sine_reg0   <= 36'sb10011101111000101100111101010011101;
        end
        6460: begin
            cosine_reg0 <= 36'sb100110110011011001101011011001111110;
            sine_reg0   <= 36'sb10011101110011110000010111110101100;
        end
        6461: begin
            cosine_reg0 <= 36'sb100110110010111010101100110011110010;
            sine_reg0   <= 36'sb10011101101110110011101100010001111;
        end
        6462: begin
            cosine_reg0 <= 36'sb100110110010011011101111001011110011;
            sine_reg0   <= 36'sb10011101101001110110111010101001010;
        end
        6463: begin
            cosine_reg0 <= 36'sb100110110001111100110010100010000000;
            sine_reg0   <= 36'sb10011101100100111010000010111011100;
        end
        6464: begin
            cosine_reg0 <= 36'sb100110110001011101110110110110011100;
            sine_reg0   <= 36'sb10011101011111111101000101001000111;
        end
        6465: begin
            cosine_reg0 <= 36'sb100110110000111110111100001001001000;
            sine_reg0   <= 36'sb10011101011011000000000001010001110;
        end
        6466: begin
            cosine_reg0 <= 36'sb100110110000100000000010011010000101;
            sine_reg0   <= 36'sb10011101010110000010110111010110010;
        end
        6467: begin
            cosine_reg0 <= 36'sb100110110000000001001001101001010011;
            sine_reg0   <= 36'sb10011101010001000101100111010110011;
        end
        6468: begin
            cosine_reg0 <= 36'sb100110101111100010010001110110110101;
            sine_reg0   <= 36'sb10011101001100001000010001010010101;
        end
        6469: begin
            cosine_reg0 <= 36'sb100110101111000011011011000010101100;
            sine_reg0   <= 36'sb10011101000111001010110101001010111;
        end
        6470: begin
            cosine_reg0 <= 36'sb100110101110100100100101001100111000;
            sine_reg0   <= 36'sb10011101000010001101010010111111100;
        end
        6471: begin
            cosine_reg0 <= 36'sb100110101110000101110000010101011011;
            sine_reg0   <= 36'sb10011100111101001111101010110000110;
        end
        6472: begin
            cosine_reg0 <= 36'sb100110101101100110111100011100010110;
            sine_reg0   <= 36'sb10011100111000010001111100011110101;
        end
        6473: begin
            cosine_reg0 <= 36'sb100110101101001000001001100001101010;
            sine_reg0   <= 36'sb10011100110011010100001000001001100;
        end
        6474: begin
            cosine_reg0 <= 36'sb100110101100101001010111100101011001;
            sine_reg0   <= 36'sb10011100101110010110001101110001011;
        end
        6475: begin
            cosine_reg0 <= 36'sb100110101100001010100110100111100011;
            sine_reg0   <= 36'sb10011100101001011000001101010110101;
        end
        6476: begin
            cosine_reg0 <= 36'sb100110101011101011110110101000001010;
            sine_reg0   <= 36'sb10011100100100011010000110111001011;
        end
        6477: begin
            cosine_reg0 <= 36'sb100110101011001101000111100111001111;
            sine_reg0   <= 36'sb10011100011111011011111010011001110;
        end
        6478: begin
            cosine_reg0 <= 36'sb100110101010101110011001100100110011;
            sine_reg0   <= 36'sb10011100011010011101100111111000000;
        end
        6479: begin
            cosine_reg0 <= 36'sb100110101010001111101100100000110111;
            sine_reg0   <= 36'sb10011100010101011111001111010100011;
        end
        6480: begin
            cosine_reg0 <= 36'sb100110101001110001000000011011011101;
            sine_reg0   <= 36'sb10011100010000100000110000101110111;
        end
        6481: begin
            cosine_reg0 <= 36'sb100110101001010010010101010100100110;
            sine_reg0   <= 36'sb10011100001011100010001100001000000;
        end
        6482: begin
            cosine_reg0 <= 36'sb100110101000110011101011001100010010;
            sine_reg0   <= 36'sb10011100000110100011100001011111101;
        end
        6483: begin
            cosine_reg0 <= 36'sb100110101000010101000010000010100100;
            sine_reg0   <= 36'sb10011100000001100100110000110110001;
        end
        6484: begin
            cosine_reg0 <= 36'sb100110100111110110011001110111011100;
            sine_reg0   <= 36'sb10011011111100100101111010001011110;
        end
        6485: begin
            cosine_reg0 <= 36'sb100110100111010111110010101010111011;
            sine_reg0   <= 36'sb10011011110111100110111101100000100;
        end
        6486: begin
            cosine_reg0 <= 36'sb100110100110111001001100011101000011;
            sine_reg0   <= 36'sb10011011110010100111111010110100101;
        end
        6487: begin
            cosine_reg0 <= 36'sb100110100110011010100111001101110101;
            sine_reg0   <= 36'sb10011011101101101000110010001000011;
        end
        6488: begin
            cosine_reg0 <= 36'sb100110100101111100000010111101010001;
            sine_reg0   <= 36'sb10011011101000101001100011011100000;
        end
        6489: begin
            cosine_reg0 <= 36'sb100110100101011101011111101011011010;
            sine_reg0   <= 36'sb10011011100011101010001110101111100;
        end
        6490: begin
            cosine_reg0 <= 36'sb100110100100111110111101011000010000;
            sine_reg0   <= 36'sb10011011011110101010110100000011010;
        end
        6491: begin
            cosine_reg0 <= 36'sb100110100100100000011100000011110101;
            sine_reg0   <= 36'sb10011011011001101011010011010111011;
        end
        6492: begin
            cosine_reg0 <= 36'sb100110100100000001111011101110001001;
            sine_reg0   <= 36'sb10011011010100101011101100101100000;
        end
        6493: begin
            cosine_reg0 <= 36'sb100110100011100011011100010111001110;
            sine_reg0   <= 36'sb10011011001111101100000000000001011;
        end
        6494: begin
            cosine_reg0 <= 36'sb100110100011000100111101111111000110;
            sine_reg0   <= 36'sb10011011001010101100001101010111110;
        end
        6495: begin
            cosine_reg0 <= 36'sb100110100010100110100000100101110000;
            sine_reg0   <= 36'sb10011011000101101100010100101111010;
        end
        6496: begin
            cosine_reg0 <= 36'sb100110100010001000000100001011001111;
            sine_reg0   <= 36'sb10011011000000101100010110001000001;
        end
        6497: begin
            cosine_reg0 <= 36'sb100110100001101001101000101111100011;
            sine_reg0   <= 36'sb10011010111011101100010001100010100;
        end
        6498: begin
            cosine_reg0 <= 36'sb100110100001001011001110010010101110;
            sine_reg0   <= 36'sb10011010110110101100000110111110101;
        end
        6499: begin
            cosine_reg0 <= 36'sb100110100000101100110100110100110001;
            sine_reg0   <= 36'sb10011010110001101011110110011100101;
        end
        6500: begin
            cosine_reg0 <= 36'sb100110100000001110011100010101101101;
            sine_reg0   <= 36'sb10011010101100101011011111111100101;
        end
        6501: begin
            cosine_reg0 <= 36'sb100110011111110000000100110101100011;
            sine_reg0   <= 36'sb10011010100111101011000011011111000;
        end
        6502: begin
            cosine_reg0 <= 36'sb100110011111010001101110010100010101;
            sine_reg0   <= 36'sb10011010100010101010100001000100000;
        end
        6503: begin
            cosine_reg0 <= 36'sb100110011110110011011000110010000011;
            sine_reg0   <= 36'sb10011010011101101001111000101011100;
        end
        6504: begin
            cosine_reg0 <= 36'sb100110011110010101000100001110101111;
            sine_reg0   <= 36'sb10011010011000101001001010010110000;
        end
        6505: begin
            cosine_reg0 <= 36'sb100110011101110110110000101010011010;
            sine_reg0   <= 36'sb10011010010011101000010110000011100;
        end
        6506: begin
            cosine_reg0 <= 36'sb100110011101011000011110000101000101;
            sine_reg0   <= 36'sb10011010001110100111011011110100010;
        end
        6507: begin
            cosine_reg0 <= 36'sb100110011100111010001100011110110010;
            sine_reg0   <= 36'sb10011010001001100110011011101000100;
        end
        6508: begin
            cosine_reg0 <= 36'sb100110011100011011111011110111100000;
            sine_reg0   <= 36'sb10011010000100100101010101100000011;
        end
        6509: begin
            cosine_reg0 <= 36'sb100110011011111101101100001111010011;
            sine_reg0   <= 36'sb10011001111111100100001001011100001;
        end
        6510: begin
            cosine_reg0 <= 36'sb100110011011011111011101100110001010;
            sine_reg0   <= 36'sb10011001111010100010110111011011111;
        end
        6511: begin
            cosine_reg0 <= 36'sb100110011011000001001111111100000111;
            sine_reg0   <= 36'sb10011001110101100001011111011111111;
        end
        6512: begin
            cosine_reg0 <= 36'sb100110011010100011000011010001001011;
            sine_reg0   <= 36'sb10011001110000100000000001101000011;
        end
        6513: begin
            cosine_reg0 <= 36'sb100110011010000100110111100101010111;
            sine_reg0   <= 36'sb10011001101011011110011101110101011;
        end
        6514: begin
            cosine_reg0 <= 36'sb100110011001100110101100111000101101;
            sine_reg0   <= 36'sb10011001100110011100110100000111010;
        end
        6515: begin
            cosine_reg0 <= 36'sb100110011001001000100011001011001101;
            sine_reg0   <= 36'sb10011001100001011011000100011110001;
        end
        6516: begin
            cosine_reg0 <= 36'sb100110011000101010011010011100111001;
            sine_reg0   <= 36'sb10011001011100011001001110111010001;
        end
        6517: begin
            cosine_reg0 <= 36'sb100110011000001100010010101101110010;
            sine_reg0   <= 36'sb10011001010111010111010011011011101;
        end
        6518: begin
            cosine_reg0 <= 36'sb100110010111101110001011111101111001;
            sine_reg0   <= 36'sb10011001010010010101010010000010101;
        end
        6519: begin
            cosine_reg0 <= 36'sb100110010111010000000110001101001111;
            sine_reg0   <= 36'sb10011001001101010011001010101111011;
        end
        6520: begin
            cosine_reg0 <= 36'sb100110010110110010000001011011110110;
            sine_reg0   <= 36'sb10011001001000010000111101100010010;
        end
        6521: begin
            cosine_reg0 <= 36'sb100110010110010011111101101001101110;
            sine_reg0   <= 36'sb10011001000011001110101010011011010;
        end
        6522: begin
            cosine_reg0 <= 36'sb100110010101110101111010110110111001;
            sine_reg0   <= 36'sb10011000111110001100010001011010100;
        end
        6523: begin
            cosine_reg0 <= 36'sb100110010101010111111001000011011000;
            sine_reg0   <= 36'sb10011000111001001001110010100000011;
        end
        6524: begin
            cosine_reg0 <= 36'sb100110010100111001111000001111001100;
            sine_reg0   <= 36'sb10011000110100000111001101101101000;
        end
        6525: begin
            cosine_reg0 <= 36'sb100110010100011011111000011010010110;
            sine_reg0   <= 36'sb10011000101111000100100011000000101;
        end
        6526: begin
            cosine_reg0 <= 36'sb100110010011111101111001100100110111;
            sine_reg0   <= 36'sb10011000101010000001110010011011011;
        end
        6527: begin
            cosine_reg0 <= 36'sb100110010011011111111011101110110001;
            sine_reg0   <= 36'sb10011000100100111110111011111101011;
        end
        6528: begin
            cosine_reg0 <= 36'sb100110010011000001111110111000000100;
            sine_reg0   <= 36'sb10011000011111111011111111100111000;
        end
        6529: begin
            cosine_reg0 <= 36'sb100110010010100100000011000000110010;
            sine_reg0   <= 36'sb10011000011010111000111101011000010;
        end
        6530: begin
            cosine_reg0 <= 36'sb100110010010000110001000001000111100;
            sine_reg0   <= 36'sb10011000010101110101110101010001100;
        end
        6531: begin
            cosine_reg0 <= 36'sb100110010001101000001110010000100100;
            sine_reg0   <= 36'sb10011000010000110010100111010010111;
        end
        6532: begin
            cosine_reg0 <= 36'sb100110010001001010010101010111101001;
            sine_reg0   <= 36'sb10011000001011101111010011011100100;
        end
        6533: begin
            cosine_reg0 <= 36'sb100110010000101100011101011110001110;
            sine_reg0   <= 36'sb10011000000110101011111001101110101;
        end
        6534: begin
            cosine_reg0 <= 36'sb100110010000001110100110100100010011;
            sine_reg0   <= 36'sb10011000000001101000011010001001100;
        end
        6535: begin
            cosine_reg0 <= 36'sb100110001111110000110000101001111011;
            sine_reg0   <= 36'sb10010111111100100100110100101101010;
        end
        6536: begin
            cosine_reg0 <= 36'sb100110001111010010111011101111000101;
            sine_reg0   <= 36'sb10010111110111100001001001011010000;
        end
        6537: begin
            cosine_reg0 <= 36'sb100110001110110101000111110011110011;
            sine_reg0   <= 36'sb10010111110010011101011000010000001;
        end
        6538: begin
            cosine_reg0 <= 36'sb100110001110010111010100111000000110;
            sine_reg0   <= 36'sb10010111101101011001100001001111110;
        end
        6539: begin
            cosine_reg0 <= 36'sb100110001101111001100010111100000000;
            sine_reg0   <= 36'sb10010111101000010101100100011001000;
        end
        6540: begin
            cosine_reg0 <= 36'sb100110001101011011110001111111100001;
            sine_reg0   <= 36'sb10010111100011010001100001101100001;
        end
        6541: begin
            cosine_reg0 <= 36'sb100110001100111110000010000010101010;
            sine_reg0   <= 36'sb10010111011110001101011001001001011;
        end
        6542: begin
            cosine_reg0 <= 36'sb100110001100100000010011000101011110;
            sine_reg0   <= 36'sb10010111011001001001001010110000110;
        end
        6543: begin
            cosine_reg0 <= 36'sb100110001100000010100101000111111100;
            sine_reg0   <= 36'sb10010111010100000100110110100010101;
        end
        6544: begin
            cosine_reg0 <= 36'sb100110001011100100111000001010000110;
            sine_reg0   <= 36'sb10010111001111000000011100011111010;
        end
        6545: begin
            cosine_reg0 <= 36'sb100110001011000111001100001011111110;
            sine_reg0   <= 36'sb10010111001001111011111100100110101;
        end
        6546: begin
            cosine_reg0 <= 36'sb100110001010101001100001001101100100;
            sine_reg0   <= 36'sb10010111000100110111010110111001000;
        end
        6547: begin
            cosine_reg0 <= 36'sb100110001010001011110111001110111001;
            sine_reg0   <= 36'sb10010110111111110010101011010110110;
        end
        6548: begin
            cosine_reg0 <= 36'sb100110001001101110001110001111111111;
            sine_reg0   <= 36'sb10010110111010101101111001111111110;
        end
        6549: begin
            cosine_reg0 <= 36'sb100110001001010000100110010000110111;
            sine_reg0   <= 36'sb10010110110101101001000010110100100;
        end
        6550: begin
            cosine_reg0 <= 36'sb100110001000110010111111010001100001;
            sine_reg0   <= 36'sb10010110110000100100000101110101000;
        end
        6551: begin
            cosine_reg0 <= 36'sb100110001000010101011001010010000000;
            sine_reg0   <= 36'sb10010110101011011111000011000001101;
        end
        6552: begin
            cosine_reg0 <= 36'sb100110000111110111110100010010010100;
            sine_reg0   <= 36'sb10010110100110011001111010011010011;
        end
        6553: begin
            cosine_reg0 <= 36'sb100110000111011010010000010010011110;
            sine_reg0   <= 36'sb10010110100001010100101011111111101;
        end
        6554: begin
            cosine_reg0 <= 36'sb100110000110111100101101010010100000;
            sine_reg0   <= 36'sb10010110011100001111010111110001011;
        end
        6555: begin
            cosine_reg0 <= 36'sb100110000110011111001011010010011010;
            sine_reg0   <= 36'sb10010110010111001001111101110000000;
        end
        6556: begin
            cosine_reg0 <= 36'sb100110000110000001101010010010001110;
            sine_reg0   <= 36'sb10010110010010000100011101111011100;
        end
        6557: begin
            cosine_reg0 <= 36'sb100110000101100100001010010001111101;
            sine_reg0   <= 36'sb10010110001100111110111000010100010;
        end
        6558: begin
            cosine_reg0 <= 36'sb100110000101000110101011010001101000;
            sine_reg0   <= 36'sb10010110000111111001001100111010100;
        end
        6559: begin
            cosine_reg0 <= 36'sb100110000100101001001101010001010000;
            sine_reg0   <= 36'sb10010110000010110011011011101110010;
        end
        6560: begin
            cosine_reg0 <= 36'sb100110000100001011110000010000110110;
            sine_reg0   <= 36'sb10010101111101101101100100101111110;
        end
        6561: begin
            cosine_reg0 <= 36'sb100110000011101110010100010000011100;
            sine_reg0   <= 36'sb10010101111000100111100111111111010;
        end
        6562: begin
            cosine_reg0 <= 36'sb100110000011010000111001010000000011;
            sine_reg0   <= 36'sb10010101110011100001100101011101000;
        end
        6563: begin
            cosine_reg0 <= 36'sb100110000010110011011111001111101011;
            sine_reg0   <= 36'sb10010101101110011011011101001001000;
        end
        6564: begin
            cosine_reg0 <= 36'sb100110000010010110000110001111010110;
            sine_reg0   <= 36'sb10010101101001010101001111000011101;
        end
        6565: begin
            cosine_reg0 <= 36'sb100110000001111000101110001111000101;
            sine_reg0   <= 36'sb10010101100100001110111011001101000;
        end
        6566: begin
            cosine_reg0 <= 36'sb100110000001011011010111001110111001;
            sine_reg0   <= 36'sb10010101011111001000100001100101011;
        end
        6567: begin
            cosine_reg0 <= 36'sb100110000000111110000001001110110011;
            sine_reg0   <= 36'sb10010101011010000010000010001100111;
        end
        6568: begin
            cosine_reg0 <= 36'sb100110000000100000101100001110110100;
            sine_reg0   <= 36'sb10010101010100111011011101000011110;
        end
        6569: begin
            cosine_reg0 <= 36'sb100110000000000011011000001110111111;
            sine_reg0   <= 36'sb10010101001111110100110010001010001;
        end
        6570: begin
            cosine_reg0 <= 36'sb100101111111100110000101001111010010;
            sine_reg0   <= 36'sb10010101001010101110000001100000011;
        end
        6571: begin
            cosine_reg0 <= 36'sb100101111111001000110011001111110001;
            sine_reg0   <= 36'sb10010101000101100111001011000110100;
        end
        6572: begin
            cosine_reg0 <= 36'sb100101111110101011100010010000011011;
            sine_reg0   <= 36'sb10010101000000100000001110111100101;
        end
        6573: begin
            cosine_reg0 <= 36'sb100101111110001110010010010001010011;
            sine_reg0   <= 36'sb10010100111011011001001101000011010;
        end
        6574: begin
            cosine_reg0 <= 36'sb100101111101110001000011010010011000;
            sine_reg0   <= 36'sb10010100110110010010000101011010011;
        end
        6575: begin
            cosine_reg0 <= 36'sb100101111101010011110101010011101101;
            sine_reg0   <= 36'sb10010100110001001010111000000010010;
        end
        6576: begin
            cosine_reg0 <= 36'sb100101111100110110101000010101010010;
            sine_reg0   <= 36'sb10010100101100000011100100111011000;
        end
        6577: begin
            cosine_reg0 <= 36'sb100101111100011001011100010111001001;
            sine_reg0   <= 36'sb10010100100110111100001100000100111;
        end
        6578: begin
            cosine_reg0 <= 36'sb100101111011111100010001011001010010;
            sine_reg0   <= 36'sb10010100100001110100101101100000001;
        end
        6579: begin
            cosine_reg0 <= 36'sb100101111011011111000111011011101111;
            sine_reg0   <= 36'sb10010100011100101101001001001100111;
        end
        6580: begin
            cosine_reg0 <= 36'sb100101111011000001111110011110100001;
            sine_reg0   <= 36'sb10010100010111100101011111001011011;
        end
        6581: begin
            cosine_reg0 <= 36'sb100101111010100100110110100001101001;
            sine_reg0   <= 36'sb10010100010010011101101111011011110;
        end
        6582: begin
            cosine_reg0 <= 36'sb100101111010000111101111100101001000;
            sine_reg0   <= 36'sb10010100001101010101111001111110010;
        end
        6583: begin
            cosine_reg0 <= 36'sb100101111001101010101001101001000000;
            sine_reg0   <= 36'sb10010100001000001101111110110011000;
        end
        6584: begin
            cosine_reg0 <= 36'sb100101111001001101100100101101010001;
            sine_reg0   <= 36'sb10010100000011000101111101111010011;
        end
        6585: begin
            cosine_reg0 <= 36'sb100101111000110000100000110001111100;
            sine_reg0   <= 36'sb10010011111101111101110111010100011;
        end
        6586: begin
            cosine_reg0 <= 36'sb100101111000010011011101110111000011;
            sine_reg0   <= 36'sb10010011111000110101101011000001010;
        end
        6587: begin
            cosine_reg0 <= 36'sb100101110111110110011011111100100111;
            sine_reg0   <= 36'sb10010011110011101101011001000001010;
        end
        6588: begin
            cosine_reg0 <= 36'sb100101110111011001011011000010101000;
            sine_reg0   <= 36'sb10010011101110100101000001010100101;
        end
        6589: begin
            cosine_reg0 <= 36'sb100101110110111100011011001001001001;
            sine_reg0   <= 36'sb10010011101001011100100011111011011;
        end
        6590: begin
            cosine_reg0 <= 36'sb100101110110011111011100010000001001;
            sine_reg0   <= 36'sb10010011100100010100000000110110000;
        end
        6591: begin
            cosine_reg0 <= 36'sb100101110110000010011110010111101011;
            sine_reg0   <= 36'sb10010011011111001011011000000100011;
        end
        6592: begin
            cosine_reg0 <= 36'sb100101110101100101100001011111101111;
            sine_reg0   <= 36'sb10010011011010000010101001100110111;
        end
        6593: begin
            cosine_reg0 <= 36'sb100101110101001000100101101000010111;
            sine_reg0   <= 36'sb10010011010100111001110101011101101;
        end
        6594: begin
            cosine_reg0 <= 36'sb100101110100101011101010110001100011;
            sine_reg0   <= 36'sb10010011001111110000111011101000111;
        end
        6595: begin
            cosine_reg0 <= 36'sb100101110100001110110000111011010101;
            sine_reg0   <= 36'sb10010011001010100111111100001000111;
        end
        6596: begin
            cosine_reg0 <= 36'sb100101110011110001111000000101101110;
            sine_reg0   <= 36'sb10010011000101011110110110111101101;
        end
        6597: begin
            cosine_reg0 <= 36'sb100101110011010101000000010000101110;
            sine_reg0   <= 36'sb10010011000000010101101100000111101;
        end
        6598: begin
            cosine_reg0 <= 36'sb100101110010111000001001011100011000;
            sine_reg0   <= 36'sb10010010111011001100011011100110110;
        end
        6599: begin
            cosine_reg0 <= 36'sb100101110010011011010011101000101100;
            sine_reg0   <= 36'sb10010010110110000011000101011011100;
        end
        6600: begin
            cosine_reg0 <= 36'sb100101110001111110011110110101101011;
            sine_reg0   <= 36'sb10010010110000111001101001100101110;
        end
        6601: begin
            cosine_reg0 <= 36'sb100101110001100001101011000011010110;
            sine_reg0   <= 36'sb10010010101011110000001000000110000;
        end
        6602: begin
            cosine_reg0 <= 36'sb100101110001000100111000010001101111;
            sine_reg0   <= 36'sb10010010100110100110100000111100010;
        end
        6603: begin
            cosine_reg0 <= 36'sb100101110000101000000110100000110110;
            sine_reg0   <= 36'sb10010010100001011100110100001000111;
        end
        6604: begin
            cosine_reg0 <= 36'sb100101110000001011010101110000101101;
            sine_reg0   <= 36'sb10010010011100010011000001101011111;
        end
        6605: begin
            cosine_reg0 <= 36'sb100101101111101110100110000001010101;
            sine_reg0   <= 36'sb10010010010111001001001001100101101;
        end
        6606: begin
            cosine_reg0 <= 36'sb100101101111010001110111010010101111;
            sine_reg0   <= 36'sb10010010010001111111001011110110001;
        end
        6607: begin
            cosine_reg0 <= 36'sb100101101110110101001001100100111100;
            sine_reg0   <= 36'sb10010010001100110101001000011101110;
        end
        6608: begin
            cosine_reg0 <= 36'sb100101101110011000011100110111111100;
            sine_reg0   <= 36'sb10010010000111101010111111011100110;
        end
        6609: begin
            cosine_reg0 <= 36'sb100101101101111011110001001011110011;
            sine_reg0   <= 36'sb10010010000010100000110000110011001;
        end
        6610: begin
            cosine_reg0 <= 36'sb100101101101011111000110100000011111;
            sine_reg0   <= 36'sb10010001111101010110011100100001001;
        end
        6611: begin
            cosine_reg0 <= 36'sb100101101101000010011100110110000011;
            sine_reg0   <= 36'sb10010001111000001100000010100111000;
        end
        6612: begin
            cosine_reg0 <= 36'sb100101101100100101110100001100011111;
            sine_reg0   <= 36'sb10010001110011000001100011000100111;
        end
        6613: begin
            cosine_reg0 <= 36'sb100101101100001001001100100011110101;
            sine_reg0   <= 36'sb10010001101101110110111101111011001;
        end
        6614: begin
            cosine_reg0 <= 36'sb100101101011101100100101111100000110;
            sine_reg0   <= 36'sb10010001101000101100010011001001110;
        end
        6615: begin
            cosine_reg0 <= 36'sb100101101011010000000000010101010011;
            sine_reg0   <= 36'sb10010001100011100001100010110001001;
        end
        6616: begin
            cosine_reg0 <= 36'sb100101101010110011011011101111011101;
            sine_reg0   <= 36'sb10010001011110010110101100110001010;
        end
        6617: begin
            cosine_reg0 <= 36'sb100101101010010110111000001010100100;
            sine_reg0   <= 36'sb10010001011001001011110001001010100;
        end
        6618: begin
            cosine_reg0 <= 36'sb100101101001111010010101100110101011;
            sine_reg0   <= 36'sb10010001010100000000101111111101000;
        end
        6619: begin
            cosine_reg0 <= 36'sb100101101001011101110100000011110010;
            sine_reg0   <= 36'sb10010001001110110101101001001001000;
        end
        6620: begin
            cosine_reg0 <= 36'sb100101101001000001010011100001111011;
            sine_reg0   <= 36'sb10010001001001101010011100101110101;
        end
        6621: begin
            cosine_reg0 <= 36'sb100101101000100100110100000001000110;
            sine_reg0   <= 36'sb10010001000100011111001010101110000;
        end
        6622: begin
            cosine_reg0 <= 36'sb100101101000001000010101100001010100;
            sine_reg0   <= 36'sb10010000111111010011110011000111101;
        end
        6623: begin
            cosine_reg0 <= 36'sb100101100111101011111000000010100111;
            sine_reg0   <= 36'sb10010000111010001000010101111011011;
        end
        6624: begin
            cosine_reg0 <= 36'sb100101100111001111011011100101000000;
            sine_reg0   <= 36'sb10010000110100111100110011001001100;
        end
        6625: begin
            cosine_reg0 <= 36'sb100101100110110011000000001000100000;
            sine_reg0   <= 36'sb10010000101111110001001010110010011;
        end
        6626: begin
            cosine_reg0 <= 36'sb100101100110010110100101101101000111;
            sine_reg0   <= 36'sb10010000101010100101011100110110001;
        end
        6627: begin
            cosine_reg0 <= 36'sb100101100101111010001100010010111000;
            sine_reg0   <= 36'sb10010000100101011001101001010100111;
        end
        6628: begin
            cosine_reg0 <= 36'sb100101100101011101110011111001110011;
            sine_reg0   <= 36'sb10010000100000001101110000001111000;
        end
        6629: begin
            cosine_reg0 <= 36'sb100101100101000001011100100001111001;
            sine_reg0   <= 36'sb10010000011011000001110001100100100;
        end
        6630: begin
            cosine_reg0 <= 36'sb100101100100100101000110001011001011;
            sine_reg0   <= 36'sb10010000010101110101101101010101101;
        end
        6631: begin
            cosine_reg0 <= 36'sb100101100100001000110000110101101011;
            sine_reg0   <= 36'sb10010000010000101001100011100010100;
        end
        6632: begin
            cosine_reg0 <= 36'sb100101100011101100011100100001011001;
            sine_reg0   <= 36'sb10010000001011011101010100001011101;
        end
        6633: begin
            cosine_reg0 <= 36'sb100101100011010000001001001110010111;
            sine_reg0   <= 36'sb10010000000110010000111111010000111;
        end
        6634: begin
            cosine_reg0 <= 36'sb100101100010110011110110111100100110;
            sine_reg0   <= 36'sb10010000000001000100100100110010101;
        end
        6635: begin
            cosine_reg0 <= 36'sb100101100010010111100101101100000110;
            sine_reg0   <= 36'sb10001111111011111000000100110001000;
        end
        6636: begin
            cosine_reg0 <= 36'sb100101100001111011010101011100111010;
            sine_reg0   <= 36'sb10001111110110101011011111001100010;
        end
        6637: begin
            cosine_reg0 <= 36'sb100101100001011111000110001111000001;
            sine_reg0   <= 36'sb10001111110001011110110100000100101;
        end
        6638: begin
            cosine_reg0 <= 36'sb100101100001000010111000000010011101;
            sine_reg0   <= 36'sb10001111101100010010000011011010001;
        end
        6639: begin
            cosine_reg0 <= 36'sb100101100000100110101010110111001111;
            sine_reg0   <= 36'sb10001111100111000101001101001101001;
        end
        6640: begin
            cosine_reg0 <= 36'sb100101100000001010011110101101011001;
            sine_reg0   <= 36'sb10001111100001111000010001011101111;
        end
        6641: begin
            cosine_reg0 <= 36'sb100101011111101110010011100100111011;
            sine_reg0   <= 36'sb10001111011100101011010000001100011;
        end
        6642: begin
            cosine_reg0 <= 36'sb100101011111010010001001011101110110;
            sine_reg0   <= 36'sb10001111010111011110001001011000111;
        end
        6643: begin
            cosine_reg0 <= 36'sb100101011110110110000000011000001100;
            sine_reg0   <= 36'sb10001111010010010000111101000011110;
        end
        6644: begin
            cosine_reg0 <= 36'sb100101011110011001111000010011111101;
            sine_reg0   <= 36'sb10001111001101000011101011001101000;
        end
        6645: begin
            cosine_reg0 <= 36'sb100101011101111101110001010001001011;
            sine_reg0   <= 36'sb10001111000111110110010011110101000;
        end
        6646: begin
            cosine_reg0 <= 36'sb100101011101100001101011001111110111;
            sine_reg0   <= 36'sb10001111000010101000110110111011111;
        end
        6647: begin
            cosine_reg0 <= 36'sb100101011101000101100110010000000001;
            sine_reg0   <= 36'sb10001110111101011011010100100001101;
        end
        6648: begin
            cosine_reg0 <= 36'sb100101011100101001100010010001101100;
            sine_reg0   <= 36'sb10001110111000001101101100100110111;
        end
        6649: begin
            cosine_reg0 <= 36'sb100101011100001101011111010100110111;
            sine_reg0   <= 36'sb10001110110010111111111111001011011;
        end
        6650: begin
            cosine_reg0 <= 36'sb100101011011110001011101011001100101;
            sine_reg0   <= 36'sb10001110101101110010001100001111101;
        end
        6651: begin
            cosine_reg0 <= 36'sb100101011011010101011100011111110101;
            sine_reg0   <= 36'sb10001110101000100100010011110011110;
        end
        6652: begin
            cosine_reg0 <= 36'sb100101011010111001011100100111101010;
            sine_reg0   <= 36'sb10001110100011010110010101111000000;
        end
        6653: begin
            cosine_reg0 <= 36'sb100101011010011101011101110001000100;
            sine_reg0   <= 36'sb10001110011110001000010010011100011;
        end
        6654: begin
            cosine_reg0 <= 36'sb100101011010000001011111111100000101;
            sine_reg0   <= 36'sb10001110011000111010001001100001011;
        end
        6655: begin
            cosine_reg0 <= 36'sb100101011001100101100011001000101101;
            sine_reg0   <= 36'sb10001110010011101011111011000110111;
        end
        6656: begin
            cosine_reg0 <= 36'sb100101011001001001100111010110111101;
            sine_reg0   <= 36'sb10001110001110011101100111001101011;
        end
        6657: begin
            cosine_reg0 <= 36'sb100101011000101101101100100110110111;
            sine_reg0   <= 36'sb10001110001001001111001101110100111;
        end
        6658: begin
            cosine_reg0 <= 36'sb100101011000010001110010111000011100;
            sine_reg0   <= 36'sb10001110000100000000101110111101110;
        end
        6659: begin
            cosine_reg0 <= 36'sb100101010111110101111010001011101101;
            sine_reg0   <= 36'sb10001101111110110010001010101000000;
        end
        6660: begin
            cosine_reg0 <= 36'sb100101010111011010000010100000101010;
            sine_reg0   <= 36'sb10001101111001100011100000110100000;
        end
        6661: begin
            cosine_reg0 <= 36'sb100101010110111110001011110111010101;
            sine_reg0   <= 36'sb10001101110100010100110001100001110;
        end
        6662: begin
            cosine_reg0 <= 36'sb100101010110100010010110001111110000;
            sine_reg0   <= 36'sb10001101101111000101111100110001101;
        end
        6663: begin
            cosine_reg0 <= 36'sb100101010110000110100001101001111010;
            sine_reg0   <= 36'sb10001101101001110111000010100011111;
        end
        6664: begin
            cosine_reg0 <= 36'sb100101010101101010101110000101110110;
            sine_reg0   <= 36'sb10001101100100101000000010111000100;
        end
        6665: begin
            cosine_reg0 <= 36'sb100101010101001110111011100011100011;
            sine_reg0   <= 36'sb10001101011111011000111101101111111;
        end
        6666: begin
            cosine_reg0 <= 36'sb100101010100110011001010000011000100;
            sine_reg0   <= 36'sb10001101011010001001110011001010001;
        end
        6667: begin
            cosine_reg0 <= 36'sb100101010100010111011001100100011010;
            sine_reg0   <= 36'sb10001101010100111010100011000111100;
        end
        6668: begin
            cosine_reg0 <= 36'sb100101010011111011101010000111100100;
            sine_reg0   <= 36'sb10001101001111101011001101101000001;
        end
        6669: begin
            cosine_reg0 <= 36'sb100101010011011111111011101100100110;
            sine_reg0   <= 36'sb10001101001010011011110010101100010;
        end
        6670: begin
            cosine_reg0 <= 36'sb100101010011000100001110010011011111;
            sine_reg0   <= 36'sb10001101000101001100010010010100000;
        end
        6671: begin
            cosine_reg0 <= 36'sb100101010010101000100001111100010000;
            sine_reg0   <= 36'sb10001100111111111100101100011111110;
        end
        6672: begin
            cosine_reg0 <= 36'sb100101010010001100110110100110111011;
            sine_reg0   <= 36'sb10001100111010101101000001001111100;
        end
        6673: begin
            cosine_reg0 <= 36'sb100101010001110001001100010011100001;
            sine_reg0   <= 36'sb10001100110101011101010000100011101;
        end
        6674: begin
            cosine_reg0 <= 36'sb100101010001010101100011000010000011;
            sine_reg0   <= 36'sb10001100110000001101011010011100010;
        end
        6675: begin
            cosine_reg0 <= 36'sb100101010000111001111010110010100001;
            sine_reg0   <= 36'sb10001100101010111101011110111001100;
        end
        6676: begin
            cosine_reg0 <= 36'sb100101010000011110010011100100111110;
            sine_reg0   <= 36'sb10001100100101101101011101111011110;
        end
        6677: begin
            cosine_reg0 <= 36'sb100101010000000010101101011001011010;
            sine_reg0   <= 36'sb10001100100000011101010111100011001;
        end
        6678: begin
            cosine_reg0 <= 36'sb100101001111100111001000001111110101;
            sine_reg0   <= 36'sb10001100011011001101001011101111110;
        end
        6679: begin
            cosine_reg0 <= 36'sb100101001111001011100100001000010010;
            sine_reg0   <= 36'sb10001100010101111100111010100001111;
        end
        6680: begin
            cosine_reg0 <= 36'sb100101001110110000000001000010110001;
            sine_reg0   <= 36'sb10001100010000101100100011111001110;
        end
        6681: begin
            cosine_reg0 <= 36'sb100101001110010100011110111111010011;
            sine_reg0   <= 36'sb10001100001011011100000111110111100;
        end
        6682: begin
            cosine_reg0 <= 36'sb100101001101111000111101111101111010;
            sine_reg0   <= 36'sb10001100000110001011100110011011100;
        end
        6683: begin
            cosine_reg0 <= 36'sb100101001101011101011101111110100110;
            sine_reg0   <= 36'sb10001100000000111010111111100101110;
        end
        6684: begin
            cosine_reg0 <= 36'sb100101001101000001111111000001011001;
            sine_reg0   <= 36'sb10001011111011101010010011010110100;
        end
        6685: begin
            cosine_reg0 <= 36'sb100101001100100110100001000110010011;
            sine_reg0   <= 36'sb10001011110110011001100001101110000;
        end
        6686: begin
            cosine_reg0 <= 36'sb100101001100001011000100001101010101;
            sine_reg0   <= 36'sb10001011110001001000101010101100011;
        end
        6687: begin
            cosine_reg0 <= 36'sb100101001011101111101000010110100001;
            sine_reg0   <= 36'sb10001011101011110111101110010010000;
        end
        6688: begin
            cosine_reg0 <= 36'sb100101001011010100001101100001111000;
            sine_reg0   <= 36'sb10001011100110100110101100011110111;
        end
        6689: begin
            cosine_reg0 <= 36'sb100101001010111000110011101111011011;
            sine_reg0   <= 36'sb10001011100001010101100101010011011;
        end
        6690: begin
            cosine_reg0 <= 36'sb100101001010011101011010111111001011;
            sine_reg0   <= 36'sb10001011011100000100011000101111100;
        end
        6691: begin
            cosine_reg0 <= 36'sb100101001010000010000011010001001000;
            sine_reg0   <= 36'sb10001011010110110011000110110011110;
        end
        6692: begin
            cosine_reg0 <= 36'sb100101001001100110101100100101010100;
            sine_reg0   <= 36'sb10001011010001100001101111100000000;
        end
        6693: begin
            cosine_reg0 <= 36'sb100101001001001011010110111011110000;
            sine_reg0   <= 36'sb10001011001100010000010010110100101;
        end
        6694: begin
            cosine_reg0 <= 36'sb100101001000110000000010010100011110;
            sine_reg0   <= 36'sb10001011000110111110110000110001111;
        end
        6695: begin
            cosine_reg0 <= 36'sb100101001000010100101110101111011101;
            sine_reg0   <= 36'sb10001011000001101101001001010111111;
        end
        6696: begin
            cosine_reg0 <= 36'sb100101000111111001011100001100101111;
            sine_reg0   <= 36'sb10001010111100011011011100100110110;
        end
        6697: begin
            cosine_reg0 <= 36'sb100101000111011110001010101100010110;
            sine_reg0   <= 36'sb10001010110111001001101010011110111;
        end
        6698: begin
            cosine_reg0 <= 36'sb100101000111000010111010001110010010;
            sine_reg0   <= 36'sb10001010110001110111110011000000011;
        end
        6699: begin
            cosine_reg0 <= 36'sb100101000110100111101010110010100100;
            sine_reg0   <= 36'sb10001010101100100101110110001011100;
        end
        6700: begin
            cosine_reg0 <= 36'sb100101000110001100011100011001001110;
            sine_reg0   <= 36'sb10001010100111010011110100000000010;
        end
        6701: begin
            cosine_reg0 <= 36'sb100101000101110001001111000010001111;
            sine_reg0   <= 36'sb10001010100010000001101100011111001;
        end
        6702: begin
            cosine_reg0 <= 36'sb100101000101010110000010101101101011;
            sine_reg0   <= 36'sb10001010011100101111011111101000001;
        end
        6703: begin
            cosine_reg0 <= 36'sb100101000100111010110111011011100000;
            sine_reg0   <= 36'sb10001010010111011101001101011011100;
        end
        6704: begin
            cosine_reg0 <= 36'sb100101000100011111101101001011110010;
            sine_reg0   <= 36'sb10001010010010001010110101111001100;
        end
        6705: begin
            cosine_reg0 <= 36'sb100101000100000100100011111110100000;
            sine_reg0   <= 36'sb10001010001100111000011001000010011;
        end
        6706: begin
            cosine_reg0 <= 36'sb100101000011101001011011110011101011;
            sine_reg0   <= 36'sb10001010000111100101110110110110001;
        end
        6707: begin
            cosine_reg0 <= 36'sb100101000011001110010100101011010101;
            sine_reg0   <= 36'sb10001010000010010011001111010101001;
        end
        6708: begin
            cosine_reg0 <= 36'sb100101000010110011001110100101011111;
            sine_reg0   <= 36'sb10001001111101000000100010011111100;
        end
        6709: begin
            cosine_reg0 <= 36'sb100101000010011000001001100010001010;
            sine_reg0   <= 36'sb10001001110111101101110000010101101;
        end
        6710: begin
            cosine_reg0 <= 36'sb100101000001111101000101100001010110;
            sine_reg0   <= 36'sb10001001110010011010111000110111011;
        end
        6711: begin
            cosine_reg0 <= 36'sb100101000001100010000010100011000110;
            sine_reg0   <= 36'sb10001001101101000111111100000101010;
        end
        6712: begin
            cosine_reg0 <= 36'sb100101000001000111000000100111011001;
            sine_reg0   <= 36'sb10001001100111110100111001111111011;
        end
        6713: begin
            cosine_reg0 <= 36'sb100101000000101011111111101110010001;
            sine_reg0   <= 36'sb10001001100010100001110010100101111;
        end
        6714: begin
            cosine_reg0 <= 36'sb100101000000010000111111110111101111;
            sine_reg0   <= 36'sb10001001011101001110100101111001000;
        end
        6715: begin
            cosine_reg0 <= 36'sb100100111111110110000001000011110100;
            sine_reg0   <= 36'sb10001001010111111011010011111001000;
        end
        6716: begin
            cosine_reg0 <= 36'sb100100111111011011000011010010100010;
            sine_reg0   <= 36'sb10001001010010100111111100100110001;
        end
        6717: begin
            cosine_reg0 <= 36'sb100100111111000000000110100011111000;
            sine_reg0   <= 36'sb10001001001101010100100000000000011;
        end
        6718: begin
            cosine_reg0 <= 36'sb100100111110100101001010110111111000;
            sine_reg0   <= 36'sb10001001001000000000111110001000001;
        end
        6719: begin
            cosine_reg0 <= 36'sb100100111110001010010000001110100100;
            sine_reg0   <= 36'sb10001001000010101101010110111101100;
        end
        6720: begin
            cosine_reg0 <= 36'sb100100111101101111010110100111111100;
            sine_reg0   <= 36'sb10001000111101011001101010100000110;
        end
        6721: begin
            cosine_reg0 <= 36'sb100100111101010100011110000100000001;
            sine_reg0   <= 36'sb10001000111000000101111000110010001;
        end
        6722: begin
            cosine_reg0 <= 36'sb100100111100111001100110100010110100;
            sine_reg0   <= 36'sb10001000110010110010000001110001110;
        end
        6723: begin
            cosine_reg0 <= 36'sb100100111100011110110000000100010111;
            sine_reg0   <= 36'sb10001000101101011110000101011111110;
        end
        6724: begin
            cosine_reg0 <= 36'sb100100111100000011111010101000101010;
            sine_reg0   <= 36'sb10001000101000001010000011111100100;
        end
        6725: begin
            cosine_reg0 <= 36'sb100100111011101001000110001111101110;
            sine_reg0   <= 36'sb10001000100010110101111101001000001;
        end
        6726: begin
            cosine_reg0 <= 36'sb100100111011001110010010111001100101;
            sine_reg0   <= 36'sb10001000011101100001110001000010111;
        end
        6727: begin
            cosine_reg0 <= 36'sb100100111010110011100000100110001111;
            sine_reg0   <= 36'sb10001000011000001101011111101100111;
        end
        6728: begin
            cosine_reg0 <= 36'sb100100111010011000101111010101101110;
            sine_reg0   <= 36'sb10001000010010111001001001000110100;
        end
        6729: begin
            cosine_reg0 <= 36'sb100100111001111101111111001000000010;
            sine_reg0   <= 36'sb10001000001101100100101101001111101;
        end
        6730: begin
            cosine_reg0 <= 36'sb100100111001100011001111111101001101;
            sine_reg0   <= 36'sb10001000001000010000001100001000111;
        end
        6731: begin
            cosine_reg0 <= 36'sb100100111001001000100001110101001111;
            sine_reg0   <= 36'sb10001000000010111011100101110010001;
        end
        6732: begin
            cosine_reg0 <= 36'sb100100111000101101110100110000001010;
            sine_reg0   <= 36'sb10000111111101100110111010001011101;
        end
        6733: begin
            cosine_reg0 <= 36'sb100100111000010011001000101101111111;
            sine_reg0   <= 36'sb10000111111000010010001001010101110;
        end
        6734: begin
            cosine_reg0 <= 36'sb100100110111111000011101101110101110;
            sine_reg0   <= 36'sb10000111110010111101010011010000101;
        end
        6735: begin
            cosine_reg0 <= 36'sb100100110111011101110011110010011001;
            sine_reg0   <= 36'sb10000111101101101000010111111100011;
        end
        6736: begin
            cosine_reg0 <= 36'sb100100110111000011001010111001000001;
            sine_reg0   <= 36'sb10000111101000010011010111011001010;
        end
        6737: begin
            cosine_reg0 <= 36'sb100100110110101000100011000010100110;
            sine_reg0   <= 36'sb10000111100010111110010001100111100;
        end
        6738: begin
            cosine_reg0 <= 36'sb100100110110001101111100001111001011;
            sine_reg0   <= 36'sb10000111011101101001000110100111011;
        end
        6739: begin
            cosine_reg0 <= 36'sb100100110101110011010110011110101111;
            sine_reg0   <= 36'sb10000111011000010011110110011000111;
        end
        6740: begin
            cosine_reg0 <= 36'sb100100110101011000110001110001010100;
            sine_reg0   <= 36'sb10000111010010111110100000111100011;
        end
        6741: begin
            cosine_reg0 <= 36'sb100100110100111110001110000110111010;
            sine_reg0   <= 36'sb10000111001101101001000110010010001;
        end
        6742: begin
            cosine_reg0 <= 36'sb100100110100100011101011011111100100;
            sine_reg0   <= 36'sb10000111001000010011100110011010010;
        end
        6743: begin
            cosine_reg0 <= 36'sb100100110100001001001001111011010010;
            sine_reg0   <= 36'sb10000111000010111110000001010100111;
        end
        6744: begin
            cosine_reg0 <= 36'sb100100110011101110101001011010000100;
            sine_reg0   <= 36'sb10000110111101101000010111000010010;
        end
        6745: begin
            cosine_reg0 <= 36'sb100100110011010100001001111011111100;
            sine_reg0   <= 36'sb10000110111000010010100111100010110;
        end
        6746: begin
            cosine_reg0 <= 36'sb100100110010111001101011100000111100;
            sine_reg0   <= 36'sb10000110110010111100110010110110011;
        end
        6747: begin
            cosine_reg0 <= 36'sb100100110010011111001110001001000011;
            sine_reg0   <= 36'sb10000110101101100110111000111101011;
        end
        6748: begin
            cosine_reg0 <= 36'sb100100110010000100110001110100010100;
            sine_reg0   <= 36'sb10000110101000010000111001111000000;
        end
        6749: begin
            cosine_reg0 <= 36'sb100100110001101010010110100010101110;
            sine_reg0   <= 36'sb10000110100010111010110101100110100;
        end
        6750: begin
            cosine_reg0 <= 36'sb100100110001001111111100010100010011;
            sine_reg0   <= 36'sb10000110011101100100101100001001000;
        end
        6751: begin
            cosine_reg0 <= 36'sb100100110000110101100011001001000101;
            sine_reg0   <= 36'sb10000110011000001110011101011111110;
        end
        6752: begin
            cosine_reg0 <= 36'sb100100110000011011001011000001000100;
            sine_reg0   <= 36'sb10000110010010111000001001101010111;
        end
        6753: begin
            cosine_reg0 <= 36'sb100100110000000000110011111100010000;
            sine_reg0   <= 36'sb10000110001101100001110000101010101;
        end
        6754: begin
            cosine_reg0 <= 36'sb100100101111100110011101111010101100;
            sine_reg0   <= 36'sb10000110001000001011010010011111010;
        end
        6755: begin
            cosine_reg0 <= 36'sb100100101111001100001000111100011000;
            sine_reg0   <= 36'sb10000110000010110100101111001001000;
        end
        6756: begin
            cosine_reg0 <= 36'sb100100101110110001110101000001010101;
            sine_reg0   <= 36'sb10000101111101011110000110100111111;
        end
        6757: begin
            cosine_reg0 <= 36'sb100100101110010111100010001001100100;
            sine_reg0   <= 36'sb10000101111000000111011000111100011;
        end
        6758: begin
            cosine_reg0 <= 36'sb100100101101111101010000010101000111;
            sine_reg0   <= 36'sb10000101110010110000100110000110011;
        end
        6759: begin
            cosine_reg0 <= 36'sb100100101101100010111111100011111101;
            sine_reg0   <= 36'sb10000101101101011001101110000110011;
        end
        6760: begin
            cosine_reg0 <= 36'sb100100101101001000101111110110001001;
            sine_reg0   <= 36'sb10000101101000000010110000111100011;
        end
        6761: begin
            cosine_reg0 <= 36'sb100100101100101110100001001011101011;
            sine_reg0   <= 36'sb10000101100010101011101110101000110;
        end
        6762: begin
            cosine_reg0 <= 36'sb100100101100010100010011100100100101;
            sine_reg0   <= 36'sb10000101011101010100100111001011101;
        end
        6763: begin
            cosine_reg0 <= 36'sb100100101011111010000111000000110110;
            sine_reg0   <= 36'sb10000101010111111101011010100101001;
        end
        6764: begin
            cosine_reg0 <= 36'sb100100101011011111111011100000100001;
            sine_reg0   <= 36'sb10000101010010100110001000110101101;
        end
        6765: begin
            cosine_reg0 <= 36'sb100100101011000101110001000011100110;
            sine_reg0   <= 36'sb10000101001101001110110001111101001;
        end
        6766: begin
            cosine_reg0 <= 36'sb100100101010101011100111101010000110;
            sine_reg0   <= 36'sb10000101000111110111010101111100001;
        end
        6767: begin
            cosine_reg0 <= 36'sb100100101010010001011111010100000011;
            sine_reg0   <= 36'sb10000101000010011111110100110010100;
        end
        6768: begin
            cosine_reg0 <= 36'sb100100101001110111011000000001011100;
            sine_reg0   <= 36'sb10000100111101001000001110100000101;
        end
        6769: begin
            cosine_reg0 <= 36'sb100100101001011101010001110010010100;
            sine_reg0   <= 36'sb10000100110111110000100011000110110;
        end
        6770: begin
            cosine_reg0 <= 36'sb100100101001000011001100100110101100;
            sine_reg0   <= 36'sb10000100110010011000110010100101001;
        end
        6771: begin
            cosine_reg0 <= 36'sb100100101000101001001000011110100011;
            sine_reg0   <= 36'sb10000100101101000000111100111011110;
        end
        6772: begin
            cosine_reg0 <= 36'sb100100101000001111000101011001111100;
            sine_reg0   <= 36'sb10000100100111101001000010001010111;
        end
        6773: begin
            cosine_reg0 <= 36'sb100100100111110101000011011000111000;
            sine_reg0   <= 36'sb10000100100010010001000010010010111;
        end
        6774: begin
            cosine_reg0 <= 36'sb100100100111011011000010011011010110;
            sine_reg0   <= 36'sb10000100011100111000111101010011111;
        end
        6775: begin
            cosine_reg0 <= 36'sb100100100111000001000010100001011001;
            sine_reg0   <= 36'sb10000100010111100000110011001110000;
        end
        6776: begin
            cosine_reg0 <= 36'sb100100100110100111000011101011000001;
            sine_reg0   <= 36'sb10000100010010001000100100000001100;
        end
        6777: begin
            cosine_reg0 <= 36'sb100100100110001101000101111000010000;
            sine_reg0   <= 36'sb10000100001100110000001111101110101;
        end
        6778: begin
            cosine_reg0 <= 36'sb100100100101110011001001001001000110;
            sine_reg0   <= 36'sb10000100000111010111110110010101101;
        end
        6779: begin
            cosine_reg0 <= 36'sb100100100101011001001101011101100100;
            sine_reg0   <= 36'sb10000100000001111111010111110110101;
        end
        6780: begin
            cosine_reg0 <= 36'sb100100100100111111010010110101101011;
            sine_reg0   <= 36'sb10000011111100100110110100010001110;
        end
        6781: begin
            cosine_reg0 <= 36'sb100100100100100101011001010001011101;
            sine_reg0   <= 36'sb10000011110111001110001011100111100;
        end
        6782: begin
            cosine_reg0 <= 36'sb100100100100001011100000110000111010;
            sine_reg0   <= 36'sb10000011110001110101011101110111110;
        end
        6783: begin
            cosine_reg0 <= 36'sb100100100011110001101001010100000100;
            sine_reg0   <= 36'sb10000011101100011100101011000010111;
        end
        6784: begin
            cosine_reg0 <= 36'sb100100100011010111110010111010111011;
            sine_reg0   <= 36'sb10000011100111000011110011001001000;
        end
        6785: begin
            cosine_reg0 <= 36'sb100100100010111101111101100101100000;
            sine_reg0   <= 36'sb10000011100001101010110110001010100;
        end
        6786: begin
            cosine_reg0 <= 36'sb100100100010100100001001010011110100;
            sine_reg0   <= 36'sb10000011011100010001110100000111011;
        end
        6787: begin
            cosine_reg0 <= 36'sb100100100010001010010110000101111001;
            sine_reg0   <= 36'sb10000011010110111000101101000000000;
        end
        6788: begin
            cosine_reg0 <= 36'sb100100100001110000100011111011101110;
            sine_reg0   <= 36'sb10000011010001011111100000110100100;
        end
        6789: begin
            cosine_reg0 <= 36'sb100100100001010110110010110101010111;
            sine_reg0   <= 36'sb10000011001100000110001111100101001;
        end
        6790: begin
            cosine_reg0 <= 36'sb100100100000111101000010110010110010;
            sine_reg0   <= 36'sb10000011000110101100111001010010000;
        end
        6791: begin
            cosine_reg0 <= 36'sb100100100000100011010011110100000010;
            sine_reg0   <= 36'sb10000011000001010011011101111011011;
        end
        6792: begin
            cosine_reg0 <= 36'sb100100100000001001100101111001000111;
            sine_reg0   <= 36'sb10000010111011111001111101100001100;
        end
        6793: begin
            cosine_reg0 <= 36'sb100100011111101111111001000010000010;
            sine_reg0   <= 36'sb10000010110110100000011000000100100;
        end
        6794: begin
            cosine_reg0 <= 36'sb100100011111010110001101001110110101;
            sine_reg0   <= 36'sb10000010110001000110101101100100110;
        end
        6795: begin
            cosine_reg0 <= 36'sb100100011110111100100010011111100000;
            sine_reg0   <= 36'sb10000010101011101100111110000010010;
        end
        6796: begin
            cosine_reg0 <= 36'sb100100011110100010111000110100000100;
            sine_reg0   <= 36'sb10000010100110010011001001011101011;
        end
        6797: begin
            cosine_reg0 <= 36'sb100100011110001001010000001100100010;
            sine_reg0   <= 36'sb10000010100000111001001111110110010;
        end
        6798: begin
            cosine_reg0 <= 36'sb100100011101101111101000101000111011;
            sine_reg0   <= 36'sb10000010011011011111010001001101000;
        end
        6799: begin
            cosine_reg0 <= 36'sb100100011101010110000010001001010001;
            sine_reg0   <= 36'sb10000010010110000101001101100010000;
        end
        6800: begin
            cosine_reg0 <= 36'sb100100011100111100011100101101100100;
            sine_reg0   <= 36'sb10000010010000101011000100110101011;
        end
        6801: begin
            cosine_reg0 <= 36'sb100100011100100010111000010101110101;
            sine_reg0   <= 36'sb10000010001011010000110111000111011;
        end
        6802: begin
            cosine_reg0 <= 36'sb100100011100001001010101000010000101;
            sine_reg0   <= 36'sb10000010000101110110100100011000001;
        end
        6803: begin
            cosine_reg0 <= 36'sb100100011011101111110010110010010101;
            sine_reg0   <= 36'sb10000010000000011100001100100111111;
        end
        6804: begin
            cosine_reg0 <= 36'sb100100011011010110010001100110100110;
            sine_reg0   <= 36'sb10000001111011000001101111110110111;
        end
        6805: begin
            cosine_reg0 <= 36'sb100100011010111100110001011110111010;
            sine_reg0   <= 36'sb10000001110101100111001110000101011;
        end
        6806: begin
            cosine_reg0 <= 36'sb100100011010100011010010011011010000;
            sine_reg0   <= 36'sb10000001110000001100100111010011100;
        end
        6807: begin
            cosine_reg0 <= 36'sb100100011010001001110100011011101011;
            sine_reg0   <= 36'sb10000001101010110001111011100001011;
        end
        6808: begin
            cosine_reg0 <= 36'sb100100011001110000010111100000001011;
            sine_reg0   <= 36'sb10000001100101010111001010101111011;
        end
        6809: begin
            cosine_reg0 <= 36'sb100100011001010110111011101000110000;
            sine_reg0   <= 36'sb10000001011111111100010100111101101;
        end
        6810: begin
            cosine_reg0 <= 36'sb100100011000111101100000110101011101;
            sine_reg0   <= 36'sb10000001011010100001011010001100011;
        end
        6811: begin
            cosine_reg0 <= 36'sb100100011000100100000111000110010010;
            sine_reg0   <= 36'sb10000001010101000110011010011011110;
        end
        6812: begin
            cosine_reg0 <= 36'sb100100011000001010101110011011001111;
            sine_reg0   <= 36'sb10000001001111101011010101101100000;
        end
        6813: begin
            cosine_reg0 <= 36'sb100100010111110001010110110100010111;
            sine_reg0   <= 36'sb10000001001010010000001011111101011;
        end
        6814: begin
            cosine_reg0 <= 36'sb100100010111011000000000010001101010;
            sine_reg0   <= 36'sb10000001000100110100111101010000001;
        end
        6815: begin
            cosine_reg0 <= 36'sb100100010110111110101010110011001000;
            sine_reg0   <= 36'sb10000000111111011001101001100100011;
        end
        6816: begin
            cosine_reg0 <= 36'sb100100010110100101010110011000110011;
            sine_reg0   <= 36'sb10000000111001111110010000111010011;
        end
        6817: begin
            cosine_reg0 <= 36'sb100100010110001100000011000010101101;
            sine_reg0   <= 36'sb10000000110100100010110011010010010;
        end
        6818: begin
            cosine_reg0 <= 36'sb100100010101110010110000110000110101;
            sine_reg0   <= 36'sb10000000101111000111010000101100010;
        end
        6819: begin
            cosine_reg0 <= 36'sb100100010101011001011111100011001101;
            sine_reg0   <= 36'sb10000000101001101011101001001000101;
        end
        6820: begin
            cosine_reg0 <= 36'sb100100010101000000001111011001110101;
            sine_reg0   <= 36'sb10000000100100001111111100100111101;
        end
        6821: begin
            cosine_reg0 <= 36'sb100100010100100111000000010100110000;
            sine_reg0   <= 36'sb10000000011110110100001011001001011;
        end
        6822: begin
            cosine_reg0 <= 36'sb100100010100001101110010010011111101;
            sine_reg0   <= 36'sb10000000011001011000010100101110001;
        end
        6823: begin
            cosine_reg0 <= 36'sb100100010011110100100101010111011110;
            sine_reg0   <= 36'sb10000000010011111100011001010110000;
        end
        6824: begin
            cosine_reg0 <= 36'sb100100010011011011011001011111010011;
            sine_reg0   <= 36'sb10000000001110100000011001000001010;
        end
        6825: begin
            cosine_reg0 <= 36'sb100100010011000010001110101011011110;
            sine_reg0   <= 36'sb10000000001001000100010011110000010;
        end
        6826: begin
            cosine_reg0 <= 36'sb100100010010101001000100111100000000;
            sine_reg0   <= 36'sb10000000000011101000001001100011000;
        end
        6827: begin
            cosine_reg0 <= 36'sb100100010010001111111100010000111001;
            sine_reg0   <= 36'sb1111111111110001011111010011001110;
        end
        6828: begin
            cosine_reg0 <= 36'sb100100010001110110110100101010001011;
            sine_reg0   <= 36'sb1111111111000101111100110010100110;
        end
        6829: begin
            cosine_reg0 <= 36'sb100100010001011101101110000111110111;
            sine_reg0   <= 36'sb1111111110011010011001101010100010;
        end
        6830: begin
            cosine_reg0 <= 36'sb100100010001000100101000101001111101;
            sine_reg0   <= 36'sb1111111101101110110101111011000011;
        end
        6831: begin
            cosine_reg0 <= 36'sb100100010000101011100100010000011110;
            sine_reg0   <= 36'sb1111111101000011010001100100001100;
        end
        6832: begin
            cosine_reg0 <= 36'sb100100010000010010100000111011011100;
            sine_reg0   <= 36'sb1111111100010111101100100101111100;
        end
        6833: begin
            cosine_reg0 <= 36'sb100100001111111001011110101010110111;
            sine_reg0   <= 36'sb1111111011101100000111000000011000;
        end
        6834: begin
            cosine_reg0 <= 36'sb100100001111100000011101011110110001;
            sine_reg0   <= 36'sb1111111011000000100000110011011111;
        end
        6835: begin
            cosine_reg0 <= 36'sb100100001111000111011101010111001010;
            sine_reg0   <= 36'sb1111111010010100111001111111010100;
        end
        6836: begin
            cosine_reg0 <= 36'sb100100001110101110011110010100000011;
            sine_reg0   <= 36'sb1111111001101001010010100011111000;
        end
        6837: begin
            cosine_reg0 <= 36'sb100100001110010101100000010101011101;
            sine_reg0   <= 36'sb1111111000111101101010100001001101;
        end
        6838: begin
            cosine_reg0 <= 36'sb100100001101111100100011011011011010;
            sine_reg0   <= 36'sb1111111000010010000001110111010101;
        end
        6839: begin
            cosine_reg0 <= 36'sb100100001101100011100111100101111010;
            sine_reg0   <= 36'sb1111110111100110011000100110010010;
        end
        6840: begin
            cosine_reg0 <= 36'sb100100001101001010101100110100111110;
            sine_reg0   <= 36'sb1111110110111010101110101110000100;
        end
        6841: begin
            cosine_reg0 <= 36'sb100100001100110001110011001000100111;
            sine_reg0   <= 36'sb1111110110001111000100001110101110;
        end
        6842: begin
            cosine_reg0 <= 36'sb100100001100011000111010100000110110;
            sine_reg0   <= 36'sb1111110101100011011001001000010010;
        end
        6843: begin
            cosine_reg0 <= 36'sb100100001100000000000010111101101100;
            sine_reg0   <= 36'sb1111110100110111101101011010110001;
        end
        6844: begin
            cosine_reg0 <= 36'sb100100001011100111001100011111001010;
            sine_reg0   <= 36'sb1111110100001100000001000110001101;
        end
        6845: begin
            cosine_reg0 <= 36'sb100100001011001110010111000101010001;
            sine_reg0   <= 36'sb1111110011100000010100001010100111;
        end
        6846: begin
            cosine_reg0 <= 36'sb100100001010110101100010110000000010;
            sine_reg0   <= 36'sb1111110010110100100110101000000010;
        end
        6847: begin
            cosine_reg0 <= 36'sb100100001010011100101111011111011101;
            sine_reg0   <= 36'sb1111110010001000111000011110011111;
        end
        6848: begin
            cosine_reg0 <= 36'sb100100001010000011111101010011100101;
            sine_reg0   <= 36'sb1111110001011101001001101101111111;
        end
        6849: begin
            cosine_reg0 <= 36'sb100100001001101011001100001100011001;
            sine_reg0   <= 36'sb1111110000110001011010010110100100;
        end
        6850: begin
            cosine_reg0 <= 36'sb100100001001010010011100001001111011;
            sine_reg0   <= 36'sb1111110000000101101010011000010000;
        end
        6851: begin
            cosine_reg0 <= 36'sb100100001000111001101101001100001100;
            sine_reg0   <= 36'sb1111101111011001111001110011000101;
        end
        6852: begin
            cosine_reg0 <= 36'sb100100001000100000111111010011001100;
            sine_reg0   <= 36'sb1111101110101110001000100111000100;
        end
        6853: begin
            cosine_reg0 <= 36'sb100100001000001000010010011110111101;
            sine_reg0   <= 36'sb1111101110000010010110110100010000;
        end
        6854: begin
            cosine_reg0 <= 36'sb100100000111101111100110101111011111;
            sine_reg0   <= 36'sb1111101101010110100100011010101001;
        end
        6855: begin
            cosine_reg0 <= 36'sb100100000111010110111100000100110100;
            sine_reg0   <= 36'sb1111101100101010110001011010010001;
        end
        6856: begin
            cosine_reg0 <= 36'sb100100000110111110010010011110111101;
            sine_reg0   <= 36'sb1111101011111110111101110011001010;
        end
        6857: begin
            cosine_reg0 <= 36'sb100100000110100101101001111101111001;
            sine_reg0   <= 36'sb1111101011010011001001100101010111;
        end
        6858: begin
            cosine_reg0 <= 36'sb100100000110001101000010100001101011;
            sine_reg0   <= 36'sb1111101010100111010100110000110111;
        end
        6859: begin
            cosine_reg0 <= 36'sb100100000101110100011100001010010011;
            sine_reg0   <= 36'sb1111101001111011011111010101101110;
        end
        6860: begin
            cosine_reg0 <= 36'sb100100000101011011110110110111110011;
            sine_reg0   <= 36'sb1111101001001111101001010011111101;
        end
        6861: begin
            cosine_reg0 <= 36'sb100100000101000011010010101010001011;
            sine_reg0   <= 36'sb1111101000100011110010101011100101;
        end
        6862: begin
            cosine_reg0 <= 36'sb100100000100101010101111100001011011;
            sine_reg0   <= 36'sb1111100111110111111011011100101000;
        end
        6863: begin
            cosine_reg0 <= 36'sb100100000100010010001101011101100110;
            sine_reg0   <= 36'sb1111100111001100000011100111001001;
        end
        6864: begin
            cosine_reg0 <= 36'sb100100000011111001101100011110101100;
            sine_reg0   <= 36'sb1111100110100000001011001011000111;
        end
        6865: begin
            cosine_reg0 <= 36'sb100100000011100001001100100100101110;
            sine_reg0   <= 36'sb1111100101110100010010001000100111;
        end
        6866: begin
            cosine_reg0 <= 36'sb100100000011001000101101101111101101;
            sine_reg0   <= 36'sb1111100101001000011000011111101000;
        end
        6867: begin
            cosine_reg0 <= 36'sb100100000010110000001111111111101001;
            sine_reg0   <= 36'sb1111100100011100011110010000001101;
        end
        6868: begin
            cosine_reg0 <= 36'sb100100000010010111110011010100100100;
            sine_reg0   <= 36'sb1111100011110000100011011010010111;
        end
        6869: begin
            cosine_reg0 <= 36'sb100100000001111111010111101110011111;
            sine_reg0   <= 36'sb1111100011000100100111111110001000;
        end
        6870: begin
            cosine_reg0 <= 36'sb100100000001100110111101001101011011;
            sine_reg0   <= 36'sb1111100010011000101011111011100010;
        end
        6871: begin
            cosine_reg0 <= 36'sb100100000001001110100011110001011001;
            sine_reg0   <= 36'sb1111100001101100101111010010100111;
        end
        6872: begin
            cosine_reg0 <= 36'sb100100000000110110001011011010011000;
            sine_reg0   <= 36'sb1111100001000000110010000011011000;
        end
        6873: begin
            cosine_reg0 <= 36'sb100100000000011101110100001000011100;
            sine_reg0   <= 36'sb1111100000010100110100001101110110;
        end
        6874: begin
            cosine_reg0 <= 36'sb100100000000000101011101111011100100;
            sine_reg0   <= 36'sb1111011111101000110101110010000100;
        end
        6875: begin
            cosine_reg0 <= 36'sb100011111111101101001000110011110001;
            sine_reg0   <= 36'sb1111011110111100110110110000000011;
        end
        6876: begin
            cosine_reg0 <= 36'sb100011111111010100110100110001000100;
            sine_reg0   <= 36'sb1111011110010000110111000111110101;
        end
        6877: begin
            cosine_reg0 <= 36'sb100011111110111100100001110011011111;
            sine_reg0   <= 36'sb1111011101100100110110111001011100;
        end
        6878: begin
            cosine_reg0 <= 36'sb100011111110100100001111111011000010;
            sine_reg0   <= 36'sb1111011100111000110110000100111001;
        end
        6879: begin
            cosine_reg0 <= 36'sb100011111110001011111111000111101110;
            sine_reg0   <= 36'sb1111011100001100110100101010001111;
        end
        6880: begin
            cosine_reg0 <= 36'sb100011111101110011101111011001100100;
            sine_reg0   <= 36'sb1111011011100000110010101001011101;
        end
        6881: begin
            cosine_reg0 <= 36'sb100011111101011011100000110000100101;
            sine_reg0   <= 36'sb1111011010110100110000000010101000;
        end
        6882: begin
            cosine_reg0 <= 36'sb100011111101000011010011001100110010;
            sine_reg0   <= 36'sb1111011010001000101100110101101111;
        end
        6883: begin
            cosine_reg0 <= 36'sb100011111100101011000110101110001100;
            sine_reg0   <= 36'sb1111011001011100101001000010110101;
        end
        6884: begin
            cosine_reg0 <= 36'sb100011111100010010111011010100110100;
            sine_reg0   <= 36'sb1111011000110000100100101001111100;
        end
        6885: begin
            cosine_reg0 <= 36'sb100011111011111010110001000000101010;
            sine_reg0   <= 36'sb1111011000000100011111101011000101;
        end
        6886: begin
            cosine_reg0 <= 36'sb100011111011100010100111110001110000;
            sine_reg0   <= 36'sb1111010111011000011010000110010010;
        end
        6887: begin
            cosine_reg0 <= 36'sb100011111011001010011111101000000111;
            sine_reg0   <= 36'sb1111010110101100010011111011100100;
        end
        6888: begin
            cosine_reg0 <= 36'sb100011111010110010011000100011101111;
            sine_reg0   <= 36'sb1111010110000000001101001010111110;
        end
        6889: begin
            cosine_reg0 <= 36'sb100011111010011010010010100100101010;
            sine_reg0   <= 36'sb1111010101010100000101110100100001;
        end
        6890: begin
            cosine_reg0 <= 36'sb100011111010000010001101101010111000;
            sine_reg0   <= 36'sb1111010100100111111101111000001110;
        end
        6891: begin
            cosine_reg0 <= 36'sb100011111001101010001001110110011010;
            sine_reg0   <= 36'sb1111010011111011110101010110001000;
        end
        6892: begin
            cosine_reg0 <= 36'sb100011111001010010000111000111010010;
            sine_reg0   <= 36'sb1111010011001111101100001110010000;
        end
        6893: begin
            cosine_reg0 <= 36'sb100011111000111010000101011101011111;
            sine_reg0   <= 36'sb1111010010100011100010100000100111;
        end
        6894: begin
            cosine_reg0 <= 36'sb100011111000100010000100111001000100;
            sine_reg0   <= 36'sb1111010001110111011000001101010001;
        end
        6895: begin
            cosine_reg0 <= 36'sb100011111000001010000101011010000001;
            sine_reg0   <= 36'sb1111010001001011001101010100001101;
        end
        6896: begin
            cosine_reg0 <= 36'sb100011110111110010000111000000010111;
            sine_reg0   <= 36'sb1111010000011111000001110101011111;
        end
        6897: begin
            cosine_reg0 <= 36'sb100011110111011010001001101100000110;
            sine_reg0   <= 36'sb1111001111110010110101110001000111;
        end
        6898: begin
            cosine_reg0 <= 36'sb100011110111000010001101011101010000;
            sine_reg0   <= 36'sb1111001111000110101001000111000111;
        end
        6899: begin
            cosine_reg0 <= 36'sb100011110110101010010010010011110110;
            sine_reg0   <= 36'sb1111001110011010011011110111100001;
        end
        6900: begin
            cosine_reg0 <= 36'sb100011110110010010011000001111111001;
            sine_reg0   <= 36'sb1111001101101110001110000010010111;
        end
        6901: begin
            cosine_reg0 <= 36'sb100011110101111010011111010001011001;
            sine_reg0   <= 36'sb1111001101000001111111100111101011;
        end
        6902: begin
            cosine_reg0 <= 36'sb100011110101100010100111011000011000;
            sine_reg0   <= 36'sb1111001100010101110000100111011110;
        end
        6903: begin
            cosine_reg0 <= 36'sb100011110101001010110000100100110110;
            sine_reg0   <= 36'sb1111001011101001100001000001110001;
        end
        6904: begin
            cosine_reg0 <= 36'sb100011110100110010111010110110110100;
            sine_reg0   <= 36'sb1111001010111101010000110110100111;
        end
        6905: begin
            cosine_reg0 <= 36'sb100011110100011011000110001110010100;
            sine_reg0   <= 36'sb1111001010010001000000000110000001;
        end
        6906: begin
            cosine_reg0 <= 36'sb100011110100000011010010101011010110;
            sine_reg0   <= 36'sb1111001001100100101110110000000010;
        end
        6907: begin
            cosine_reg0 <= 36'sb100011110011101011100000001101111011;
            sine_reg0   <= 36'sb1111001000111000011100110100101010;
        end
        6908: begin
            cosine_reg0 <= 36'sb100011110011010011101110110110000011;
            sine_reg0   <= 36'sb1111001000001100001010010011111011;
        end
        6909: begin
            cosine_reg0 <= 36'sb100011110010111011111110100011110001;
            sine_reg0   <= 36'sb1111000111011111110111001101110111;
        end
        6910: begin
            cosine_reg0 <= 36'sb100011110010100100001111010111000101;
            sine_reg0   <= 36'sb1111000110110011100011100010100001;
        end
        6911: begin
            cosine_reg0 <= 36'sb100011110010001100100001001111111111;
            sine_reg0   <= 36'sb1111000110000111001111010001111000;
        end
        6912: begin
            cosine_reg0 <= 36'sb100011110001110100110100001110100001;
            sine_reg0   <= 36'sb1111000101011010111010011100000000;
        end
        6913: begin
            cosine_reg0 <= 36'sb100011110001011101001000010010101011;
            sine_reg0   <= 36'sb1111000100101110100101000000111010;
        end
        6914: begin
            cosine_reg0 <= 36'sb100011110001000101011101011100011111;
            sine_reg0   <= 36'sb1111000100000010001111000000101000;
        end
        6915: begin
            cosine_reg0 <= 36'sb100011110000101101110011101011111101;
            sine_reg0   <= 36'sb1111000011010101111000011011001011;
        end
        6916: begin
            cosine_reg0 <= 36'sb100011110000010110001011000001000111;
            sine_reg0   <= 36'sb1111000010101001100001010000100100;
        end
        6917: begin
            cosine_reg0 <= 36'sb100011101111111110100011011011111101;
            sine_reg0   <= 36'sb1111000001111101001001100000110111;
        end
        6918: begin
            cosine_reg0 <= 36'sb100011101111100110111100111100100000;
            sine_reg0   <= 36'sb1111000001010000110001001100000100;
        end
        6919: begin
            cosine_reg0 <= 36'sb100011101111001111010111100010110001;
            sine_reg0   <= 36'sb1111000000100100011000010010001110;
        end
        6920: begin
            cosine_reg0 <= 36'sb100011101110110111110011001110110000;
            sine_reg0   <= 36'sb1110111111110111111110110011010101;
        end
        6921: begin
            cosine_reg0 <= 36'sb100011101110100000010000000000100000;
            sine_reg0   <= 36'sb1110111111001011100100101111011011;
        end
        6922: begin
            cosine_reg0 <= 36'sb100011101110001000101101111000000001;
            sine_reg0   <= 36'sb1110111110011111001010000110100100;
        end
        6923: begin
            cosine_reg0 <= 36'sb100011101101110001001100110101010011;
            sine_reg0   <= 36'sb1110111101110010101110111000101111;
        end
        6924: begin
            cosine_reg0 <= 36'sb100011101101011001101100111000010111;
            sine_reg0   <= 36'sb1110111101000110010011000101111111;
        end
        6925: begin
            cosine_reg0 <= 36'sb100011101101000010001110000001010000;
            sine_reg0   <= 36'sb1110111100011001110110101110010101;
        end
        6926: begin
            cosine_reg0 <= 36'sb100011101100101010110000001111111100;
            sine_reg0   <= 36'sb1110111011101101011001110001110011;
        end
        6927: begin
            cosine_reg0 <= 36'sb100011101100010011010011100100011110;
            sine_reg0   <= 36'sb1110111011000000111100010000011100;
        end
        6928: begin
            cosine_reg0 <= 36'sb100011101011111011110111111110110110;
            sine_reg0   <= 36'sb1110111010010100011110001010010000;
        end
        6929: begin
            cosine_reg0 <= 36'sb100011101011100100011101011111000101;
            sine_reg0   <= 36'sb1110111001100111111111011111010001;
        end
        6930: begin
            cosine_reg0 <= 36'sb100011101011001101000100000101001100;
            sine_reg0   <= 36'sb1110111000111011100000001111100001;
        end
        6931: begin
            cosine_reg0 <= 36'sb100011101010110101101011110001001100;
            sine_reg0   <= 36'sb1110111000001111000000011011000010;
        end
        6932: begin
            cosine_reg0 <= 36'sb100011101010011110010100100011000110;
            sine_reg0   <= 36'sb1110110111100010100000000001110110;
        end
        6933: begin
            cosine_reg0 <= 36'sb100011101010000110111110011010111011;
            sine_reg0   <= 36'sb1110110110110101111111000011111110;
        end
        6934: begin
            cosine_reg0 <= 36'sb100011101001101111101001011000101011;
            sine_reg0   <= 36'sb1110110110001001011101100001011011;
        end
        6935: begin
            cosine_reg0 <= 36'sb100011101001011000010101011100010111;
            sine_reg0   <= 36'sb1110110101011100111011011010010000;
        end
        6936: begin
            cosine_reg0 <= 36'sb100011101001000001000010100110000001;
            sine_reg0   <= 36'sb1110110100110000011000101110011111;
        end
        6937: begin
            cosine_reg0 <= 36'sb100011101000101001110000110101101001;
            sine_reg0   <= 36'sb1110110100000011110101011110001000;
        end
        6938: begin
            cosine_reg0 <= 36'sb100011101000010010100000001011010001;
            sine_reg0   <= 36'sb1110110011010111010001101001001111;
        end
        6939: begin
            cosine_reg0 <= 36'sb100011100111111011010000100110111000;
            sine_reg0   <= 36'sb1110110010101010101101001111110011;
        end
        6940: begin
            cosine_reg0 <= 36'sb100011100111100100000010001000100001;
            sine_reg0   <= 36'sb1110110001111110001000010001111000;
        end
        6941: begin
            cosine_reg0 <= 36'sb100011100111001100110100110000001011;
            sine_reg0   <= 36'sb1110110001010001100010101111011111;
        end
        6942: begin
            cosine_reg0 <= 36'sb100011100110110101101000011101111001;
            sine_reg0   <= 36'sb1110110000100100111100101000101010;
        end
        6943: begin
            cosine_reg0 <= 36'sb100011100110011110011101010001101001;
            sine_reg0   <= 36'sb1110101111111000010101111101011001;
        end
        6944: begin
            cosine_reg0 <= 36'sb100011100110000111010011001011011111;
            sine_reg0   <= 36'sb1110101111001011101110101101110000;
        end
        6945: begin
            cosine_reg0 <= 36'sb100011100101110000001010001011011010;
            sine_reg0   <= 36'sb1110101110011111000110111001110000;
        end
        6946: begin
            cosine_reg0 <= 36'sb100011100101011001000010010001011011;
            sine_reg0   <= 36'sb1110101101110010011110100001011010;
        end
        6947: begin
            cosine_reg0 <= 36'sb100011100101000001111011011101100011;
            sine_reg0   <= 36'sb1110101101000101110101100100110001;
        end
        6948: begin
            cosine_reg0 <= 36'sb100011100100101010110101101111110100;
            sine_reg0   <= 36'sb1110101100011001001100000011110101;
        end
        6949: begin
            cosine_reg0 <= 36'sb100011100100010011110001001000001101;
            sine_reg0   <= 36'sb1110101011101100100001111110101001;
        end
        6950: begin
            cosine_reg0 <= 36'sb100011100011111100101101100110110001;
            sine_reg0   <= 36'sb1110101010111111110111010101001111;
        end
        6951: begin
            cosine_reg0 <= 36'sb100011100011100101101011001011011111;
            sine_reg0   <= 36'sb1110101010010011001100000111100111;
        end
        6952: begin
            cosine_reg0 <= 36'sb100011100011001110101001110110011001;
            sine_reg0   <= 36'sb1110101001100110100000010101110101;
        end
        6953: begin
            cosine_reg0 <= 36'sb100011100010110111101001100111100000;
            sine_reg0   <= 36'sb1110101000111001110011111111111001;
        end
        6954: begin
            cosine_reg0 <= 36'sb100011100010100000101010011110110100;
            sine_reg0   <= 36'sb1110101000001101000111000101110101;
        end
        6955: begin
            cosine_reg0 <= 36'sb100011100010001001101100011100010110;
            sine_reg0   <= 36'sb1110100111100000011001100111101011;
        end
        6956: begin
            cosine_reg0 <= 36'sb100011100001110010101111100000001000;
            sine_reg0   <= 36'sb1110100110110011101011100101011101;
        end
        6957: begin
            cosine_reg0 <= 36'sb100011100001011011110011101010001001;
            sine_reg0   <= 36'sb1110100110000110111100111111001100;
        end
        6958: begin
            cosine_reg0 <= 36'sb100011100001000100111000111010011100;
            sine_reg0   <= 36'sb1110100101011010001101110100111011;
        end
        6959: begin
            cosine_reg0 <= 36'sb100011100000101101111111010001000001;
            sine_reg0   <= 36'sb1110100100101101011110000110101011;
        end
        6960: begin
            cosine_reg0 <= 36'sb100011100000010111000110101101111000;
            sine_reg0   <= 36'sb1110100100000000101101110100011101;
        end
        6961: begin
            cosine_reg0 <= 36'sb100011100000000000001111010001000011;
            sine_reg0   <= 36'sb1110100011010011111100111110010011;
        end
        6962: begin
            cosine_reg0 <= 36'sb100011011111101001011000111010100011;
            sine_reg0   <= 36'sb1110100010100111001011100100010000;
        end
        6963: begin
            cosine_reg0 <= 36'sb100011011111010010100011101010011000;
            sine_reg0   <= 36'sb1110100001111010011001100110010100;
        end
        6964: begin
            cosine_reg0 <= 36'sb100011011110111011101111100000100011;
            sine_reg0   <= 36'sb1110100001001101100111000100100010;
        end
        6965: begin
            cosine_reg0 <= 36'sb100011011110100100111100011101000101;
            sine_reg0   <= 36'sb1110100000100000110011111110111011;
        end
        6966: begin
            cosine_reg0 <= 36'sb100011011110001110001010100000000000;
            sine_reg0   <= 36'sb1110011111110100000000010101100010;
        end
        6967: begin
            cosine_reg0 <= 36'sb100011011101110111011001101001010011;
            sine_reg0   <= 36'sb1110011111000111001100001000010110;
        end
        6968: begin
            cosine_reg0 <= 36'sb100011011101100000101001111001000000;
            sine_reg0   <= 36'sb1110011110011010010111010111011100;
        end
        6969: begin
            cosine_reg0 <= 36'sb100011011101001001111011001111001000;
            sine_reg0   <= 36'sb1110011101101101100010000010110011;
        end
        6970: begin
            cosine_reg0 <= 36'sb100011011100110011001101101011101100;
            sine_reg0   <= 36'sb1110011101000000101100001010011111;
        end
        6971: begin
            cosine_reg0 <= 36'sb100011011100011100100001001110101011;
            sine_reg0   <= 36'sb1110011100010011110101101110100000;
        end
        6972: begin
            cosine_reg0 <= 36'sb100011011100000101110101111000001001;
            sine_reg0   <= 36'sb1110011011100110111110101110111000;
        end
        6973: begin
            cosine_reg0 <= 36'sb100011011011101111001011101000000100;
            sine_reg0   <= 36'sb1110011010111010000111001011101010;
        end
        6974: begin
            cosine_reg0 <= 36'sb100011011011011000100010011110011110;
            sine_reg0   <= 36'sb1110011010001101001111000100110110;
        end
        6975: begin
            cosine_reg0 <= 36'sb100011011011000001111010011011011001;
            sine_reg0   <= 36'sb1110011001100000010110011010011111;
        end
        6976: begin
            cosine_reg0 <= 36'sb100011011010101011010011011110110100;
            sine_reg0   <= 36'sb1110011000110011011101001100100110;
        end
        6977: begin
            cosine_reg0 <= 36'sb100011011010010100101101101000110001;
            sine_reg0   <= 36'sb1110011000000110100011011011001101;
        end
        6978: begin
            cosine_reg0 <= 36'sb100011011001111110001000111001010000;
            sine_reg0   <= 36'sb1110010111011001101001000110010110;
        end
        6979: begin
            cosine_reg0 <= 36'sb100011011001100111100101010000010011;
            sine_reg0   <= 36'sb1110010110101100101110001110000010;
        end
        6980: begin
            cosine_reg0 <= 36'sb100011011001010001000010101101111010;
            sine_reg0   <= 36'sb1110010101111111110010110010010100;
        end
        6981: begin
            cosine_reg0 <= 36'sb100011011000111010100001010010000110;
            sine_reg0   <= 36'sb1110010101010010110110110011001100;
        end
        6982: begin
            cosine_reg0 <= 36'sb100011011000100100000000111100111000;
            sine_reg0   <= 36'sb1110010100100101111010010000101101;
        end
        6983: begin
            cosine_reg0 <= 36'sb100011011000001101100001101110010010;
            sine_reg0   <= 36'sb1110010011111000111101001010111001;
        end
        6984: begin
            cosine_reg0 <= 36'sb100011010111110111000011100110010010;
            sine_reg0   <= 36'sb1110010011001011111111100001110000;
        end
        6985: begin
            cosine_reg0 <= 36'sb100011010111100000100110100100111100;
            sine_reg0   <= 36'sb1110010010011111000001010101010110;
        end
        6986: begin
            cosine_reg0 <= 36'sb100011010111001010001010101010001111;
            sine_reg0   <= 36'sb1110010001110010000010100101101011;
        end
        6987: begin
            cosine_reg0 <= 36'sb100011010110110011101111110110001100;
            sine_reg0   <= 36'sb1110010001000101000011010010110001;
        end
        6988: begin
            cosine_reg0 <= 36'sb100011010110011101010110001000110101;
            sine_reg0   <= 36'sb1110010000011000000011011100101011;
        end
        6989: begin
            cosine_reg0 <= 36'sb100011010110000110111101100010001010;
            sine_reg0   <= 36'sb1110001111101011000011000011011001;
        end
        6990: begin
            cosine_reg0 <= 36'sb100011010101110000100110000010001011;
            sine_reg0   <= 36'sb1110001110111110000010000110111110;
        end
        6991: begin
            cosine_reg0 <= 36'sb100011010101011010001111101000111011;
            sine_reg0   <= 36'sb1110001110010001000000100111011011;
        end
        6992: begin
            cosine_reg0 <= 36'sb100011010101000011111010010110011001;
            sine_reg0   <= 36'sb1110001101100011111110100100110010;
        end
        6993: begin
            cosine_reg0 <= 36'sb100011010100101101100110001010100110;
            sine_reg0   <= 36'sb1110001100110110111011111111000101;
        end
        6994: begin
            cosine_reg0 <= 36'sb100011010100010111010011000101100100;
            sine_reg0   <= 36'sb1110001100001001111000110110010110;
        end
        6995: begin
            cosine_reg0 <= 36'sb100011010100000001000001000111010100;
            sine_reg0   <= 36'sb1110001011011100110101001010100101;
        end
        6996: begin
            cosine_reg0 <= 36'sb100011010011101010110000001111110101;
            sine_reg0   <= 36'sb1110001010101111110000111011110110;
        end
        6997: begin
            cosine_reg0 <= 36'sb100011010011010100100000011111001001;
            sine_reg0   <= 36'sb1110001010000010101100001010001001;
        end
        6998: begin
            cosine_reg0 <= 36'sb100011010010111110010001110101010001;
            sine_reg0   <= 36'sb1110001001010101100110110101100001;
        end
        6999: begin
            cosine_reg0 <= 36'sb100011010010101000000100010010001110;
            sine_reg0   <= 36'sb1110001000101000100000111101111111;
        end
        7000: begin
            cosine_reg0 <= 36'sb100011010010010001110111110110000001;
            sine_reg0   <= 36'sb1110000111111011011010100011100100;
        end
        7001: begin
            cosine_reg0 <= 36'sb100011010001111011101100100000101001;
            sine_reg0   <= 36'sb1110000111001110010011100110010100;
        end
        7002: begin
            cosine_reg0 <= 36'sb100011010001100101100010010010001001;
            sine_reg0   <= 36'sb1110000110100001001100000110001111;
        end
        7003: begin
            cosine_reg0 <= 36'sb100011010001001111011001001010100010;
            sine_reg0   <= 36'sb1110000101110100000100000011010110;
        end
        7004: begin
            cosine_reg0 <= 36'sb100011010000111001010001001001110011;
            sine_reg0   <= 36'sb1110000101000110111011011101101101;
        end
        7005: begin
            cosine_reg0 <= 36'sb100011010000100011001010001111111110;
            sine_reg0   <= 36'sb1110000100011001110010010101010101;
        end
        7006: begin
            cosine_reg0 <= 36'sb100011010000001101000100011101000011;
            sine_reg0   <= 36'sb1110000011101100101000101010001110;
        end
        7007: begin
            cosine_reg0 <= 36'sb100011001111110110111111110001000100;
            sine_reg0   <= 36'sb1110000010111111011110011100011100;
        end
        7008: begin
            cosine_reg0 <= 36'sb100011001111100000111100001100000010;
            sine_reg0   <= 36'sb1110000010010010010011101100000000;
        end
        7009: begin
            cosine_reg0 <= 36'sb100011001111001010111001101101111100;
            sine_reg0   <= 36'sb1110000001100101001000011000111011;
        end
        7010: begin
            cosine_reg0 <= 36'sb100011001110110100111000010110110101;
            sine_reg0   <= 36'sb1110000000110111111100100011001111;
        end
        7011: begin
            cosine_reg0 <= 36'sb100011001110011110111000000110101101;
            sine_reg0   <= 36'sb1110000000001010110000001010111111;
        end
        7012: begin
            cosine_reg0 <= 36'sb100011001110001000111000111101100100;
            sine_reg0   <= 36'sb1101111111011101100011010000001011;
        end
        7013: begin
            cosine_reg0 <= 36'sb100011001101110010111010111011011100;
            sine_reg0   <= 36'sb1101111110110000010101110010110110;
        end
        7014: begin
            cosine_reg0 <= 36'sb100011001101011100111110000000010110;
            sine_reg0   <= 36'sb1101111110000011000111110011000001;
        end
        7015: begin
            cosine_reg0 <= 36'sb100011001101000111000010001100010001;
            sine_reg0   <= 36'sb1101111101010101111001010000101111;
        end
        7016: begin
            cosine_reg0 <= 36'sb100011001100110001000111011111010000;
            sine_reg0   <= 36'sb1101111100101000101010001100000000;
        end
        7017: begin
            cosine_reg0 <= 36'sb100011001100011011001101111001010011;
            sine_reg0   <= 36'sb1101111011111011011010100100110110;
        end
        7018: begin
            cosine_reg0 <= 36'sb100011001100000101010101011010011011;
            sine_reg0   <= 36'sb1101111011001110001010011011010100;
        end
        7019: begin
            cosine_reg0 <= 36'sb100011001011101111011110000010101000;
            sine_reg0   <= 36'sb1101111010100000111001101111011010;
        end
        7020: begin
            cosine_reg0 <= 36'sb100011001011011001100111110001111100;
            sine_reg0   <= 36'sb1101111001110011101000100001001100;
        end
        7021: begin
            cosine_reg0 <= 36'sb100011001011000011110010101000011000;
            sine_reg0   <= 36'sb1101111001000110010110110000101010;
        end
        7022: begin
            cosine_reg0 <= 36'sb100011001010101101111110100101111011;
            sine_reg0   <= 36'sb1101111000011001000100011101110110;
        end
        7023: begin
            cosine_reg0 <= 36'sb100011001010011000001011101010101000;
            sine_reg0   <= 36'sb1101110111101011110001101000110010;
        end
        7024: begin
            cosine_reg0 <= 36'sb100011001010000010011001110110011110;
            sine_reg0   <= 36'sb1101110110111110011110010001100000;
        end
        7025: begin
            cosine_reg0 <= 36'sb100011001001101100101001001001011111;
            sine_reg0   <= 36'sb1101110110010001001010011000000010;
        end
        7026: begin
            cosine_reg0 <= 36'sb100011001001010110111001100011101100;
            sine_reg0   <= 36'sb1101110101100011110101111100011000;
        end
        7027: begin
            cosine_reg0 <= 36'sb100011001001000001001011000101000101;
            sine_reg0   <= 36'sb1101110100110110100000111110100110;
        end
        7028: begin
            cosine_reg0 <= 36'sb100011001000101011011101101101101100;
            sine_reg0   <= 36'sb1101110100001001001011011110101100;
        end
        7029: begin
            cosine_reg0 <= 36'sb100011001000010101110001011101100000;
            sine_reg0   <= 36'sb1101110011011011110101011100101101;
        end
        7030: begin
            cosine_reg0 <= 36'sb100011001000000000000110010100100100;
            sine_reg0   <= 36'sb1101110010101110011110111000101010;
        end
        7031: begin
            cosine_reg0 <= 36'sb100011000111101010011100010010110111;
            sine_reg0   <= 36'sb1101110010000001000111110010100101;
        end
        7032: begin
            cosine_reg0 <= 36'sb100011000111010100110011011000011010;
            sine_reg0   <= 36'sb1101110001010011110000001010011111;
        end
        7033: begin
            cosine_reg0 <= 36'sb100011000110111111001011100101010000;
            sine_reg0   <= 36'sb1101110000100110011000000000011011;
        end
        7034: begin
            cosine_reg0 <= 36'sb100011000110101001100100111001010111;
            sine_reg0   <= 36'sb1101101111111000111111010100011011;
        end
        7035: begin
            cosine_reg0 <= 36'sb100011000110010011111111010100110010;
            sine_reg0   <= 36'sb1101101111001011100110000110011111;
        end
        7036: begin
            cosine_reg0 <= 36'sb100011000101111110011010110111100000;
            sine_reg0   <= 36'sb1101101110011110001100010110101010;
        end
        7037: begin
            cosine_reg0 <= 36'sb100011000101101000110111100001100011;
            sine_reg0   <= 36'sb1101101101110000110010000100111101;
        end
        7038: begin
            cosine_reg0 <= 36'sb100011000101010011010101010010111100;
            sine_reg0   <= 36'sb1101101101000011010111010001011011;
        end
        7039: begin
            cosine_reg0 <= 36'sb100011000100111101110100001011101011;
            sine_reg0   <= 36'sb1101101100010101111011111100000100;
        end
        7040: begin
            cosine_reg0 <= 36'sb100011000100101000010100001011110010;
            sine_reg0   <= 36'sb1101101011101000100000000100111100;
        end
        7041: begin
            cosine_reg0 <= 36'sb100011000100010010110101010011010000;
            sine_reg0   <= 36'sb1101101010111011000011101100000011;
        end
        7042: begin
            cosine_reg0 <= 36'sb100011000011111101010111100010001000;
            sine_reg0   <= 36'sb1101101010001101100110110001011010;
        end
        7043: begin
            cosine_reg0 <= 36'sb100011000011100111111010111000011001;
            sine_reg0   <= 36'sb1101101001100000001001010101000101;
        end
        7044: begin
            cosine_reg0 <= 36'sb100011000011010010011111010110000100;
            sine_reg0   <= 36'sb1101101000110010101011010111000101;
        end
        7045: begin
            cosine_reg0 <= 36'sb100011000010111101000100111011001100;
            sine_reg0   <= 36'sb1101101000000101001100110111011011;
        end
        7046: begin
            cosine_reg0 <= 36'sb100011000010100111101011100111101111;
            sine_reg0   <= 36'sb1101100111010111101101110110001010;
        end
        7047: begin
            cosine_reg0 <= 36'sb100011000010010010010011011011101111;
            sine_reg0   <= 36'sb1101100110101010001110010011010010;
        end
        7048: begin
            cosine_reg0 <= 36'sb100011000001111100111100010111001101;
            sine_reg0   <= 36'sb1101100101111100101110001110110110;
        end
        7049: begin
            cosine_reg0 <= 36'sb100011000001100111100110011010001010;
            sine_reg0   <= 36'sb1101100101001111001101101000111000;
        end
        7050: begin
            cosine_reg0 <= 36'sb100011000001010010010001100100100111;
            sine_reg0   <= 36'sb1101100100100001101100100001011000;
        end
        7051: begin
            cosine_reg0 <= 36'sb100011000000111100111101110110100011;
            sine_reg0   <= 36'sb1101100011110100001010111000011010;
        end
        7052: begin
            cosine_reg0 <= 36'sb100011000000100111101011010000000001;
            sine_reg0   <= 36'sb1101100011000110101000101101111111;
        end
        7053: begin
            cosine_reg0 <= 36'sb100011000000010010011001110001000001;
            sine_reg0   <= 36'sb1101100010011001000110000010001000;
        end
        7054: begin
            cosine_reg0 <= 36'sb100010111111111101001001011001100011;
            sine_reg0   <= 36'sb1101100001101011100010110100110111;
        end
        7055: begin
            cosine_reg0 <= 36'sb100010111111100111111010001001101010;
            sine_reg0   <= 36'sb1101100000111101111111000110001110;
        end
        7056: begin
            cosine_reg0 <= 36'sb100010111111010010101100000001010100;
            sine_reg0   <= 36'sb1101100000010000011010110110001111;
        end
        7057: begin
            cosine_reg0 <= 36'sb100010111110111101011111000000100100;
            sine_reg0   <= 36'sb1101011111100010110110000100111100;
        end
        7058: begin
            cosine_reg0 <= 36'sb100010111110101000010011000111011010;
            sine_reg0   <= 36'sb1101011110110101010000110010010110;
        end
        7059: begin
            cosine_reg0 <= 36'sb100010111110010011001000010101110111;
            sine_reg0   <= 36'sb1101011110000111101010111110011111;
        end
        7060: begin
            cosine_reg0 <= 36'sb100010111101111101111110101011111011;
            sine_reg0   <= 36'sb1101011101011010000100101001011001;
        end
        7061: begin
            cosine_reg0 <= 36'sb100010111101101000110110001001101000;
            sine_reg0   <= 36'sb1101011100101100011101110011000101;
        end
        7062: begin
            cosine_reg0 <= 36'sb100010111101010011101110101110111111;
            sine_reg0   <= 36'sb1101011011111110110110011011100110;
        end
        7063: begin
            cosine_reg0 <= 36'sb100010111100111110101000011011111111;
            sine_reg0   <= 36'sb1101011011010001001110100010111101;
        end
        7064: begin
            cosine_reg0 <= 36'sb100010111100101001100011010000101010;
            sine_reg0   <= 36'sb1101011010100011100110001001001011;
        end
        7065: begin
            cosine_reg0 <= 36'sb100010111100010100011111001101000010;
            sine_reg0   <= 36'sb1101011001110101111101001110010011;
        end
        7066: begin
            cosine_reg0 <= 36'sb100010111011111111011100010001000101;
            sine_reg0   <= 36'sb1101011001001000010011110010010111;
        end
        7067: begin
            cosine_reg0 <= 36'sb100010111011101010011010011100110111;
            sine_reg0   <= 36'sb1101011000011010101001110101011000;
        end
        7068: begin
            cosine_reg0 <= 36'sb100010111011010101011001110000010110;
            sine_reg0   <= 36'sb1101010111101100111111010111010111;
        end
        7069: begin
            cosine_reg0 <= 36'sb100010111011000000011010001011100100;
            sine_reg0   <= 36'sb1101010110111111010100011000010111;
        end
        7070: begin
            cosine_reg0 <= 36'sb100010111010101011011011101110100010;
            sine_reg0   <= 36'sb1101010110010001101000111000011010;
        end
        7071: begin
            cosine_reg0 <= 36'sb100010111010010110011110011001010001;
            sine_reg0   <= 36'sb1101010101100011111100110111100001;
        end
        7072: begin
            cosine_reg0 <= 36'sb100010111010000001100010001011110001;
            sine_reg0   <= 36'sb1101010100110110010000010101101101;
        end
        7073: begin
            cosine_reg0 <= 36'sb100010111001101100100111000110000100;
            sine_reg0   <= 36'sb1101010100001000100011010011000010;
        end
        7074: begin
            cosine_reg0 <= 36'sb100010111001010111101101001000001001;
            sine_reg0   <= 36'sb1101010011011010110101101111011111;
        end
        7075: begin
            cosine_reg0 <= 36'sb100010111001000010110100010010000011;
            sine_reg0   <= 36'sb1101010010101101000111101011001000;
        end
        7076: begin
            cosine_reg0 <= 36'sb100010111000101101111100100011110001;
            sine_reg0   <= 36'sb1101010001111111011001000101111110;
        end
        7077: begin
            cosine_reg0 <= 36'sb100010111000011001000101111101010100;
            sine_reg0   <= 36'sb1101010001010001101010000000000011;
        end
        7078: begin
            cosine_reg0 <= 36'sb100010111000000100010000011110101110;
            sine_reg0   <= 36'sb1101010000100011111010011001011000;
        end
        7079: begin
            cosine_reg0 <= 36'sb100010110111101111011100000111111111;
            sine_reg0   <= 36'sb1101001111110110001010010010000000;
        end
        7080: begin
            cosine_reg0 <= 36'sb100010110111011010101000111001000111;
            sine_reg0   <= 36'sb1101001111001000011001101001111011;
        end
        7081: begin
            cosine_reg0 <= 36'sb100010110111000101110110110010001001;
            sine_reg0   <= 36'sb1101001110011010101000100001001100;
        end
        7082: begin
            cosine_reg0 <= 36'sb100010110110110001000101110011000100;
            sine_reg0   <= 36'sb1101001101101100110110110111110101;
        end
        7083: begin
            cosine_reg0 <= 36'sb100010110110011100010101111011111001;
            sine_reg0   <= 36'sb1101001100111111000100101101110111;
        end
        7084: begin
            cosine_reg0 <= 36'sb100010110110000111100111001100101001;
            sine_reg0   <= 36'sb1101001100010001010010000011010100;
        end
        7085: begin
            cosine_reg0 <= 36'sb100010110101110010111001100101010101;
            sine_reg0   <= 36'sb1101001011100011011110111000001111;
        end
        7086: begin
            cosine_reg0 <= 36'sb100010110101011110001101000101111110;
            sine_reg0   <= 36'sb1101001010110101101011001100100111;
        end
        7087: begin
            cosine_reg0 <= 36'sb100010110101001001100001101110100100;
            sine_reg0   <= 36'sb1101001010000111110111000000100000;
        end
        7088: begin
            cosine_reg0 <= 36'sb100010110100110100110111011111001001;
            sine_reg0   <= 36'sb1101001001011010000010010011111011;
        end
        7089: begin
            cosine_reg0 <= 36'sb100010110100100000001110010111101100;
            sine_reg0   <= 36'sb1101001000101100001101000110111011;
        end
        7090: begin
            cosine_reg0 <= 36'sb100010110100001011100110011000010000;
            sine_reg0   <= 36'sb1101000111111110010111011001011111;
        end
        7091: begin
            cosine_reg0 <= 36'sb100010110011110110111111100000110100;
            sine_reg0   <= 36'sb1101000111010000100001001011101100;
        end
        7092: begin
            cosine_reg0 <= 36'sb100010110011100010011001110001011001;
            sine_reg0   <= 36'sb1101000110100010101010011101100001;
        end
        7093: begin
            cosine_reg0 <= 36'sb100010110011001101110101001010000001;
            sine_reg0   <= 36'sb1101000101110100110011001111000001;
        end
        7094: begin
            cosine_reg0 <= 36'sb100010110010111001010001101010101100;
            sine_reg0   <= 36'sb1101000101000110111011100000001111;
        end
        7095: begin
            cosine_reg0 <= 36'sb100010110010100100101111010011011011;
            sine_reg0   <= 36'sb1101000100011001000011010001001010;
        end
        7096: begin
            cosine_reg0 <= 36'sb100010110010010000001110000100001110;
            sine_reg0   <= 36'sb1101000011101011001010100001110110;
        end
        7097: begin
            cosine_reg0 <= 36'sb100010110001111011101101111101000111;
            sine_reg0   <= 36'sb1101000010111101010001010010010100;
        end
        7098: begin
            cosine_reg0 <= 36'sb100010110001100111001110111110000110;
            sine_reg0   <= 36'sb1101000010001111010111100010100110;
        end
        7099: begin
            cosine_reg0 <= 36'sb100010110001010010110001000111001011;
            sine_reg0   <= 36'sb1101000001100001011101010010101110;
        end
        7100: begin
            cosine_reg0 <= 36'sb100010110000111110010100011000011001;
            sine_reg0   <= 36'sb1101000000110011100010100010101100;
        end
        7101: begin
            cosine_reg0 <= 36'sb100010110000101001111000110001101111;
            sine_reg0   <= 36'sb1101000000000101100111010010100100;
        end
        7102: begin
            cosine_reg0 <= 36'sb100010110000010101011110010011001111;
            sine_reg0   <= 36'sb1100111111010111101011100010010111;
        end
        7103: begin
            cosine_reg0 <= 36'sb100010110000000001000100111100111001;
            sine_reg0   <= 36'sb1100111110101001101111010010000111;
        end
        7104: begin
            cosine_reg0 <= 36'sb100010101111101100101100101110101101;
            sine_reg0   <= 36'sb1100111101111011110010100001110101;
        end
        7105: begin
            cosine_reg0 <= 36'sb100010101111011000010101101000101110;
            sine_reg0   <= 36'sb1100111101001101110101010001100011;
        end
        7106: begin
            cosine_reg0 <= 36'sb100010101111000011111111101010111011;
            sine_reg0   <= 36'sb1100111100011111110111100001010011;
        end
        7107: begin
            cosine_reg0 <= 36'sb100010101110101111101010110101010101;
            sine_reg0   <= 36'sb1100111011110001111001010001000111;
        end
        7108: begin
            cosine_reg0 <= 36'sb100010101110011011010111000111111101;
            sine_reg0   <= 36'sb1100111011000011111010100001000001;
        end
        7109: begin
            cosine_reg0 <= 36'sb100010101110000111000100100010110100;
            sine_reg0   <= 36'sb1100111010010101111011010001000001;
        end
        7110: begin
            cosine_reg0 <= 36'sb100010101101110010110011000101111011;
            sine_reg0   <= 36'sb1100111001100111111011100001001011;
        end
        7111: begin
            cosine_reg0 <= 36'sb100010101101011110100010110001010010;
            sine_reg0   <= 36'sb1100111000111001111011010001100000;
        end
        7112: begin
            cosine_reg0 <= 36'sb100010101101001010010011100100111011;
            sine_reg0   <= 36'sb1100111000001011111010100010000001;
        end
        7113: begin
            cosine_reg0 <= 36'sb100010101100110110000101100000110101;
            sine_reg0   <= 36'sb1100110111011101111001010010110001;
        end
        7114: begin
            cosine_reg0 <= 36'sb100010101100100001111000100101000010;
            sine_reg0   <= 36'sb1100110110101111110111100011110001;
        end
        7115: begin
            cosine_reg0 <= 36'sb100010101100001101101100110001100011;
            sine_reg0   <= 36'sb1100110110000001110101010101000011;
        end
        7116: begin
            cosine_reg0 <= 36'sb100010101011111001100010000110011000;
            sine_reg0   <= 36'sb1100110101010011110010100110101001;
        end
        7117: begin
            cosine_reg0 <= 36'sb100010101011100101011000100011100010;
            sine_reg0   <= 36'sb1100110100100101101111011000100100;
        end
        7118: begin
            cosine_reg0 <= 36'sb100010101011010001010000001001000010;
            sine_reg0   <= 36'sb1100110011110111101011101010110110;
        end
        7119: begin
            cosine_reg0 <= 36'sb100010101010111101001000110110111001;
            sine_reg0   <= 36'sb1100110011001001100111011101100010;
        end
        7120: begin
            cosine_reg0 <= 36'sb100010101010101001000010101101000111;
            sine_reg0   <= 36'sb1100110010011011100010110000101000;
        end
        7121: begin
            cosine_reg0 <= 36'sb100010101010010100111101101011101101;
            sine_reg0   <= 36'sb1100110001101101011101100100001011;
        end
        7122: begin
            cosine_reg0 <= 36'sb100010101010000000111001110010101100;
            sine_reg0   <= 36'sb1100110000111111010111111000001100;
        end
        7123: begin
            cosine_reg0 <= 36'sb100010101001101100110111000010000101;
            sine_reg0   <= 36'sb1100110000010001010001101100101101;
        end
        7124: begin
            cosine_reg0 <= 36'sb100010101001011000110101011001111000;
            sine_reg0   <= 36'sb1100101111100011001011000001110001;
        end
        7125: begin
            cosine_reg0 <= 36'sb100010101001000100110100111010000111;
            sine_reg0   <= 36'sb1100101110110101000011110111011000;
        end
        7126: begin
            cosine_reg0 <= 36'sb100010101000110000110101100010110010;
            sine_reg0   <= 36'sb1100101110000110111100001101100100;
        end
        7127: begin
            cosine_reg0 <= 36'sb100010101000011100110111010011111010;
            sine_reg0   <= 36'sb1100101101011000110100000100011000;
        end
        7128: begin
            cosine_reg0 <= 36'sb100010101000001000111010001101011111;
            sine_reg0   <= 36'sb1100101100101010101011011011110101;
        end
        7129: begin
            cosine_reg0 <= 36'sb100010100111110100111110001111100010;
            sine_reg0   <= 36'sb1100101011111100100010010011111101;
        end
        7130: begin
            cosine_reg0 <= 36'sb100010100111100001000011011010000101;
            sine_reg0   <= 36'sb1100101011001110011000101100110001;
        end
        7131: begin
            cosine_reg0 <= 36'sb100010100111001101001001101101001000;
            sine_reg0   <= 36'sb1100101010100000001110100110010100;
        end
        7132: begin
            cosine_reg0 <= 36'sb100010100110111001010001001000101011;
            sine_reg0   <= 36'sb1100101001110010000100000000100111;
        end
        7133: begin
            cosine_reg0 <= 36'sb100010100110100101011001101100110000;
            sine_reg0   <= 36'sb1100101001000011111000111011101011;
        end
        7134: begin
            cosine_reg0 <= 36'sb100010100110010001100011011001010111;
            sine_reg0   <= 36'sb1100101000010101101101010111100100;
        end
        7135: begin
            cosine_reg0 <= 36'sb100010100101111101101110001110100001;
            sine_reg0   <= 36'sb1100100111100111100001010100010010;
        end
        7136: begin
            cosine_reg0 <= 36'sb100010100101101001111010001100001110;
            sine_reg0   <= 36'sb1100100110111001010100110001110111;
        end
        7137: begin
            cosine_reg0 <= 36'sb100010100101010110000111010010100001;
            sine_reg0   <= 36'sb1100100110001011000111110000010110;
        end
        7138: begin
            cosine_reg0 <= 36'sb100010100101000010010101100001011000;
            sine_reg0   <= 36'sb1100100101011100111010001111101111;
        end
        7139: begin
            cosine_reg0 <= 36'sb100010100100101110100100111000110110;
            sine_reg0   <= 36'sb1100100100101110101100010000000101;
        end
        7140: begin
            cosine_reg0 <= 36'sb100010100100011010110101011000111010;
            sine_reg0   <= 36'sb1100100100000000011101110001011001;
        end
        7141: begin
            cosine_reg0 <= 36'sb100010100100000111000111000001100110;
            sine_reg0   <= 36'sb1100100011010010001110110011101101;
        end
        7142: begin
            cosine_reg0 <= 36'sb100010100011110011011001110010111010;
            sine_reg0   <= 36'sb1100100010100011111111010111000100;
        end
        7143: begin
            cosine_reg0 <= 36'sb100010100011011111101101101100110111;
            sine_reg0   <= 36'sb1100100001110101101111011011011110;
        end
        7144: begin
            cosine_reg0 <= 36'sb100010100011001100000010101111011110;
            sine_reg0   <= 36'sb1100100001000111011111000000111110;
        end
        7145: begin
            cosine_reg0 <= 36'sb100010100010111000011000111010110000;
            sine_reg0   <= 36'sb1100100000011001001110000111100101;
        end
        7146: begin
            cosine_reg0 <= 36'sb100010100010100100110000001110101100;
            sine_reg0   <= 36'sb1100011111101010111100101111010101;
        end
        7147: begin
            cosine_reg0 <= 36'sb100010100010010001001000101011010101;
            sine_reg0   <= 36'sb1100011110111100101010111000010000;
        end
        7148: begin
            cosine_reg0 <= 36'sb100010100001111101100010010000101011;
            sine_reg0   <= 36'sb1100011110001110011000100010010111;
        end
        7149: begin
            cosine_reg0 <= 36'sb100010100001101001111100111110101111;
            sine_reg0   <= 36'sb1100011101100000000101101101101110;
        end
        7150: begin
            cosine_reg0 <= 36'sb100010100001010110011000110101100001;
            sine_reg0   <= 36'sb1100011100110001110010011010010100;
        end
        7151: begin
            cosine_reg0 <= 36'sb100010100001000010110101110101000010;
            sine_reg0   <= 36'sb1100011100000011011110101000001100;
        end
        7152: begin
            cosine_reg0 <= 36'sb100010100000101111010011111101010011;
            sine_reg0   <= 36'sb1100011011010101001010010111011001;
        end
        7153: begin
            cosine_reg0 <= 36'sb100010100000011011110011001110010100;
            sine_reg0   <= 36'sb1100011010100110110101100111111011;
        end
        7154: begin
            cosine_reg0 <= 36'sb100010100000001000010011101000000111;
            sine_reg0   <= 36'sb1100011001111000100000011001110100;
        end
        7155: begin
            cosine_reg0 <= 36'sb100010011111110100110101001010101100;
            sine_reg0   <= 36'sb1100011001001010001010101101000110;
        end
        7156: begin
            cosine_reg0 <= 36'sb100010011111100001010111110110000100;
            sine_reg0   <= 36'sb1100011000011011110100100001110100;
        end
        7157: begin
            cosine_reg0 <= 36'sb100010011111001101111011101010010000;
            sine_reg0   <= 36'sb1100010111101101011101110111111110;
        end
        7158: begin
            cosine_reg0 <= 36'sb100010011110111010100000100111010000;
            sine_reg0   <= 36'sb1100010110111111000110101111100110;
        end
        7159: begin
            cosine_reg0 <= 36'sb100010011110100111000110101101000101;
            sine_reg0   <= 36'sb1100010110010000101111001000101111;
        end
        7160: begin
            cosine_reg0 <= 36'sb100010011110010011101101111011110000;
            sine_reg0   <= 36'sb1100010101100010010111000011011010;
        end
        7161: begin
            cosine_reg0 <= 36'sb100010011110000000010110010011010001;
            sine_reg0   <= 36'sb1100010100110011111110011111101001;
        end
        7162: begin
            cosine_reg0 <= 36'sb100010011101101100111111110011101010;
            sine_reg0   <= 36'sb1100010100000101100101011101011110;
        end
        7163: begin
            cosine_reg0 <= 36'sb100010011101011001101010011100111011;
            sine_reg0   <= 36'sb1100010011010111001011111100111010;
        end
        7164: begin
            cosine_reg0 <= 36'sb100010011101000110010110001111000101;
            sine_reg0   <= 36'sb1100010010101000110001111101111111;
        end
        7165: begin
            cosine_reg0 <= 36'sb100010011100110011000011001010001001;
            sine_reg0   <= 36'sb1100010001111010010111100000110000;
        end
        7166: begin
            cosine_reg0 <= 36'sb100010011100011111110001001110000110;
            sine_reg0   <= 36'sb1100010001001011111100100101001101;
        end
        7167: begin
            cosine_reg0 <= 36'sb100010011100001100100000011010111111;
            sine_reg0   <= 36'sb1100010000011101100001001011011001;
        end
        7168: begin
            cosine_reg0 <= 36'sb100010011011111001010000110000110100;
            sine_reg0   <= 36'sb1100001111101111000101010011010101;
        end
        7169: begin
            cosine_reg0 <= 36'sb100010011011100110000010001111100110;
            sine_reg0   <= 36'sb1100001111000000101000111101000100;
        end
        7170: begin
            cosine_reg0 <= 36'sb100010011011010010110100110111010100;
            sine_reg0   <= 36'sb1100001110010010001100001000100111;
        end
        7171: begin
            cosine_reg0 <= 36'sb100010011010111111101000101000000001;
            sine_reg0   <= 36'sb1100001101100011101110110101111111;
        end
        7172: begin
            cosine_reg0 <= 36'sb100010011010101100011101100001101101;
            sine_reg0   <= 36'sb1100001100110101010001000101001111;
        end
        7173: begin
            cosine_reg0 <= 36'sb100010011010011001010011100100011000;
            sine_reg0   <= 36'sb1100001100000110110010110110011000;
        end
        7174: begin
            cosine_reg0 <= 36'sb100010011010000110001010110000000011;
            sine_reg0   <= 36'sb1100001011011000010100001001011101;
        end
        7175: begin
            cosine_reg0 <= 36'sb100010011001110011000011000100110000;
            sine_reg0   <= 36'sb1100001010101001110100111110011110;
        end
        7176: begin
            cosine_reg0 <= 36'sb100010011001011111111100100010011110;
            sine_reg0   <= 36'sb1100001001111011010101010101011110;
        end
        7177: begin
            cosine_reg0 <= 36'sb100010011001001100110111001001001111;
            sine_reg0   <= 36'sb1100001001001100110101001110011111;
        end
        7178: begin
            cosine_reg0 <= 36'sb100010011000111001110010111001000011;
            sine_reg0   <= 36'sb1100001000011110010100101001100010;
        end
        7179: begin
            cosine_reg0 <= 36'sb100010011000100110101111110001111011;
            sine_reg0   <= 36'sb1100000111101111110011100110101001;
        end
        7180: begin
            cosine_reg0 <= 36'sb100010011000010011101101110011110111;
            sine_reg0   <= 36'sb1100000111000001010010000101110110;
        end
        7181: begin
            cosine_reg0 <= 36'sb100010011000000000101100111110111001;
            sine_reg0   <= 36'sb1100000110010010110000000111001011;
        end
        7182: begin
            cosine_reg0 <= 36'sb100010010111101101101101010011000001;
            sine_reg0   <= 36'sb1100000101100100001101101010101001;
        end
        7183: begin
            cosine_reg0 <= 36'sb100010010111011010101110110000010001;
            sine_reg0   <= 36'sb1100000100110101101010110000010011;
        end
        7184: begin
            cosine_reg0 <= 36'sb100010010111000111110001010110100111;
            sine_reg0   <= 36'sb1100000100000111000111011000001001;
        end
        7185: begin
            cosine_reg0 <= 36'sb100010010110110100110101000110000110;
            sine_reg0   <= 36'sb1100000011011000100011100010001111;
        end
        7186: begin
            cosine_reg0 <= 36'sb100010010110100001111001111110101111;
            sine_reg0   <= 36'sb1100000010101001111111001110100101;
        end
        7187: begin
            cosine_reg0 <= 36'sb100010010110001111000000000000100001;
            sine_reg0   <= 36'sb1100000001111011011010011101001110;
        end
        7188: begin
            cosine_reg0 <= 36'sb100010010101111100000111001011011101;
            sine_reg0   <= 36'sb1100000001001100110101001110001011;
        end
        7189: begin
            cosine_reg0 <= 36'sb100010010101101001001111011111100101;
            sine_reg0   <= 36'sb1100000000011110001111100001011110;
        end
        7190: begin
            cosine_reg0 <= 36'sb100010010101010110011000111100111001;
            sine_reg0   <= 36'sb1011111111101111101001010111001001;
        end
        7191: begin
            cosine_reg0 <= 36'sb100010010101000011100011100011011001;
            sine_reg0   <= 36'sb1011111111000001000010101111001110;
        end
        7192: begin
            cosine_reg0 <= 36'sb100010010100110000101111010011000111;
            sine_reg0   <= 36'sb1011111110010010011011101001101110;
        end
        7193: begin
            cosine_reg0 <= 36'sb100010010100011101111100001100000011;
            sine_reg0   <= 36'sb1011111101100011110100000110101011;
        end
        7194: begin
            cosine_reg0 <= 36'sb100010010100001011001010001110001111;
            sine_reg0   <= 36'sb1011111100110101001100000110001000;
        end
        7195: begin
            cosine_reg0 <= 36'sb100010010011111000011001011001101001;
            sine_reg0   <= 36'sb1011111100000110100011101000000101;
        end
        7196: begin
            cosine_reg0 <= 36'sb100010010011100101101001101110010100;
            sine_reg0   <= 36'sb1011111011010111111010101100100101;
        end
        7197: begin
            cosine_reg0 <= 36'sb100010010011010010111011001100010001;
            sine_reg0   <= 36'sb1011111010101001010001010011101001;
        end
        7198: begin
            cosine_reg0 <= 36'sb100010010011000000001101110011011111;
            sine_reg0   <= 36'sb1011111001111010100111011101010100;
        end
        7199: begin
            cosine_reg0 <= 36'sb100010010010101101100001100011111111;
            sine_reg0   <= 36'sb1011111001001011111101001001100111;
        end
        7200: begin
            cosine_reg0 <= 36'sb100010010010011010110110011101110011;
            sine_reg0   <= 36'sb1011111000011101010010011000100011;
        end
        7201: begin
            cosine_reg0 <= 36'sb100010010010001000001100100000111010;
            sine_reg0   <= 36'sb1011110111101110100111001010001100;
        end
        7202: begin
            cosine_reg0 <= 36'sb100010010001110101100011101101010111;
            sine_reg0   <= 36'sb1011110110111111111011011110100001;
        end
        7203: begin
            cosine_reg0 <= 36'sb100010010001100010111100000011001001;
            sine_reg0   <= 36'sb1011110110010001001111010101100110;
        end
        7204: begin
            cosine_reg0 <= 36'sb100010010001010000010101100010010000;
            sine_reg0   <= 36'sb1011110101100010100010101111011100;
        end
        7205: begin
            cosine_reg0 <= 36'sb100010010000111101110000001010101111;
            sine_reg0   <= 36'sb1011110100110011110101101100000101;
        end
        7206: begin
            cosine_reg0 <= 36'sb100010010000101011001011111100100101;
            sine_reg0   <= 36'sb1011110100000101001000001011100010;
        end
        7207: begin
            cosine_reg0 <= 36'sb100010010000011000101000110111110100;
            sine_reg0   <= 36'sb1011110011010110011010001101110110;
        end
        7208: begin
            cosine_reg0 <= 36'sb100010010000000110000110111100011100;
            sine_reg0   <= 36'sb1011110010100111101011110011000010;
        end
        7209: begin
            cosine_reg0 <= 36'sb100010001111110011100110001010011101;
            sine_reg0   <= 36'sb1011110001111000111100111011001000;
        end
        7210: begin
            cosine_reg0 <= 36'sb100010001111100001000110100001111000;
            sine_reg0   <= 36'sb1011110001001010001101100110001010;
        end
        7211: begin
            cosine_reg0 <= 36'sb100010001111001110101000000010101111;
            sine_reg0   <= 36'sb1011110000011011011101110100001010;
        end
        7212: begin
            cosine_reg0 <= 36'sb100010001110111100001010101101000010;
            sine_reg0   <= 36'sb1011101111101100101101100101001001;
        end
        7213: begin
            cosine_reg0 <= 36'sb100010001110101001101110100000110001;
            sine_reg0   <= 36'sb1011101110111101111100111001001001;
        end
        7214: begin
            cosine_reg0 <= 36'sb100010001110010111010011011101111101;
            sine_reg0   <= 36'sb1011101110001111001011110000001101;
        end
        7215: begin
            cosine_reg0 <= 36'sb100010001110000100111001100100101000;
            sine_reg0   <= 36'sb1011101101100000011010001010010101;
        end
        7216: begin
            cosine_reg0 <= 36'sb100010001101110010100000110100110001;
            sine_reg0   <= 36'sb1011101100110001101000000111100100;
        end
        7217: begin
            cosine_reg0 <= 36'sb100010001101100000001001001110011001;
            sine_reg0   <= 36'sb1011101100000010110101100111111100;
        end
        7218: begin
            cosine_reg0 <= 36'sb100010001101001101110010110001100010;
            sine_reg0   <= 36'sb1011101011010100000010101011011101;
        end
        7219: begin
            cosine_reg0 <= 36'sb100010001100111011011101011110001011;
            sine_reg0   <= 36'sb1011101010100101001111010010001011;
        end
        7220: begin
            cosine_reg0 <= 36'sb100010001100101001001001010100010110;
            sine_reg0   <= 36'sb1011101001110110011011011100000111;
        end
        7221: begin
            cosine_reg0 <= 36'sb100010001100010110110110010100000011;
            sine_reg0   <= 36'sb1011101001000111100111001001010010;
        end
        7222: begin
            cosine_reg0 <= 36'sb100010001100000100100100011101010011;
            sine_reg0   <= 36'sb1011101000011000110010011001101111;
        end
        7223: begin
            cosine_reg0 <= 36'sb100010001011110010010011110000000110;
            sine_reg0   <= 36'sb1011100111101001111101001101011111;
        end
        7224: begin
            cosine_reg0 <= 36'sb100010001011100000000100001100011110;
            sine_reg0   <= 36'sb1011100110111011000111100100100100;
        end
        7225: begin
            cosine_reg0 <= 36'sb100010001011001101110101110010011011;
            sine_reg0   <= 36'sb1011100110001100010001011111000001;
        end
        7226: begin
            cosine_reg0 <= 36'sb100010001010111011101000100001111110;
            sine_reg0   <= 36'sb1011100101011101011010111100110101;
        end
        7227: begin
            cosine_reg0 <= 36'sb100010001010101001011100011011000111;
            sine_reg0   <= 36'sb1011100100101110100011111110000101;
        end
        7228: begin
            cosine_reg0 <= 36'sb100010001010010111010001011101110111;
            sine_reg0   <= 36'sb1011100011111111101100100010110001;
        end
        7229: begin
            cosine_reg0 <= 36'sb100010001010000101000111101010001111;
            sine_reg0   <= 36'sb1011100011010000110100101010111010;
        end
        7230: begin
            cosine_reg0 <= 36'sb100010001001110010111111000000010000;
            sine_reg0   <= 36'sb1011100010100001111100010110100100;
        end
        7231: begin
            cosine_reg0 <= 36'sb100010001001100000110111011111111010;
            sine_reg0   <= 36'sb1011100001110011000011100101110000;
        end
        7232: begin
            cosine_reg0 <= 36'sb100010001001001110110001001001001110;
            sine_reg0   <= 36'sb1011100001000100001010011000011111;
        end
        7233: begin
            cosine_reg0 <= 36'sb100010001000111100101011111100001100;
            sine_reg0   <= 36'sb1011100000010101010000101110110011;
        end
        7234: begin
            cosine_reg0 <= 36'sb100010001000101010100111111000110110;
            sine_reg0   <= 36'sb1011011111100110010110101000101111;
        end
        7235: begin
            cosine_reg0 <= 36'sb100010001000011000100100111111001100;
            sine_reg0   <= 36'sb1011011110110111011100000110010100;
        end
        7236: begin
            cosine_reg0 <= 36'sb100010001000000110100011001111001110;
            sine_reg0   <= 36'sb1011011110001000100001000111100011;
        end
        7237: begin
            cosine_reg0 <= 36'sb100010000111110100100010101000111110;
            sine_reg0   <= 36'sb1011011101011001100101101100011111;
        end
        7238: begin
            cosine_reg0 <= 36'sb100010000111100010100011001100011100;
            sine_reg0   <= 36'sb1011011100101010101001110101001010;
        end
        7239: begin
            cosine_reg0 <= 36'sb100010000111010000100100111001101001;
            sine_reg0   <= 36'sb1011011011111011101101100001100100;
        end
        7240: begin
            cosine_reg0 <= 36'sb100010000110111110100111110000100110;
            sine_reg0   <= 36'sb1011011011001100110000110001110001;
        end
        7241: begin
            cosine_reg0 <= 36'sb100010000110101100101011110001010010;
            sine_reg0   <= 36'sb1011011010011101110011100101110001;
        end
        7242: begin
            cosine_reg0 <= 36'sb100010000110011010110000111011110000;
            sine_reg0   <= 36'sb1011011001101110110101111101101000;
        end
        7243: begin
            cosine_reg0 <= 36'sb100010000110001000110111001111111111;
            sine_reg0   <= 36'sb1011011000111111110111111001010101;
        end
        7244: begin
            cosine_reg0 <= 36'sb100010000101110110111110101110000000;
            sine_reg0   <= 36'sb1011011000010000111001011000111100;
        end
        7245: begin
            cosine_reg0 <= 36'sb100010000101100101000111010101110100;
            sine_reg0   <= 36'sb1011010111100001111010011100011110;
        end
        7246: begin
            cosine_reg0 <= 36'sb100010000101010011010001000111011100;
            sine_reg0   <= 36'sb1011010110110010111011000011111101;
        end
        7247: begin
            cosine_reg0 <= 36'sb100010000101000001011100000010111000;
            sine_reg0   <= 36'sb1011010110000011111011001111011010;
        end
        7248: begin
            cosine_reg0 <= 36'sb100010000100101111101000001000001001;
            sine_reg0   <= 36'sb1011010101010100111010111110111001;
        end
        7249: begin
            cosine_reg0 <= 36'sb100010000100011101110101010111010000;
            sine_reg0   <= 36'sb1011010100100101111010010010011001;
        end
        7250: begin
            cosine_reg0 <= 36'sb100010000100001100000011110000001110;
            sine_reg0   <= 36'sb1011010011110110111001001001111110;
        end
        7251: begin
            cosine_reg0 <= 36'sb100010000011111010010011010011000010;
            sine_reg0   <= 36'sb1011010011000111110111100101101000;
        end
        7252: begin
            cosine_reg0 <= 36'sb100010000011101000100011111111101110;
            sine_reg0   <= 36'sb1011010010011000110101100101011010;
        end
        7253: begin
            cosine_reg0 <= 36'sb100010000011010110110101110110010011;
            sine_reg0   <= 36'sb1011010001101001110011001001010110;
        end
        7254: begin
            cosine_reg0 <= 36'sb100010000011000101001000110110110000;
            sine_reg0   <= 36'sb1011010000111010110000010001011101;
        end
        7255: begin
            cosine_reg0 <= 36'sb100010000010110011011101000001001000;
            sine_reg0   <= 36'sb1011010000001011101100111101110010;
        end
        7256: begin
            cosine_reg0 <= 36'sb100010000010100001110010010101011010;
            sine_reg0   <= 36'sb1011001111011100101001001110010101;
        end
        7257: begin
            cosine_reg0 <= 36'sb100010000010010000001000110011100111;
            sine_reg0   <= 36'sb1011001110101101100101000011001010;
        end
        7258: begin
            cosine_reg0 <= 36'sb100010000001111110100000011011110000;
            sine_reg0   <= 36'sb1011001101111110100000011100010001;
        end
        7259: begin
            cosine_reg0 <= 36'sb100010000001101100111001001101110110;
            sine_reg0   <= 36'sb1011001101001111011011011001101100;
        end
        7260: begin
            cosine_reg0 <= 36'sb100010000001011011010011001001111001;
            sine_reg0   <= 36'sb1011001100100000010101111011011110;
        end
        7261: begin
            cosine_reg0 <= 36'sb100010000001001001101110001111111001;
            sine_reg0   <= 36'sb1011001011110001010000000001100111;
        end
        7262: begin
            cosine_reg0 <= 36'sb100010000000111000001010011111111001;
            sine_reg0   <= 36'sb1011001011000010001001101100001011;
        end
        7263: begin
            cosine_reg0 <= 36'sb100010000000100110100111111001110111;
            sine_reg0   <= 36'sb1011001010010011000010111011001011;
        end
        7264: begin
            cosine_reg0 <= 36'sb100010000000010101000110011101110110;
            sine_reg0   <= 36'sb1011001001100011111011101110101000;
        end
        7265: begin
            cosine_reg0 <= 36'sb100010000000000011100110001011110101;
            sine_reg0   <= 36'sb1011001000110100110100000110100100;
        end
        7266: begin
            cosine_reg0 <= 36'sb100001111111110010000111000011110101;
            sine_reg0   <= 36'sb1011001000000101101100000011000001;
        end
        7267: begin
            cosine_reg0 <= 36'sb100001111111100000101001000101110111;
            sine_reg0   <= 36'sb1011000111010110100011100100000010;
        end
        7268: begin
            cosine_reg0 <= 36'sb100001111111001111001100010001111100;
            sine_reg0   <= 36'sb1011000110100111011010101001100111;
        end
        7269: begin
            cosine_reg0 <= 36'sb100001111110111101110000101000000100;
            sine_reg0   <= 36'sb1011000101111000010001010011110011;
        end
        7270: begin
            cosine_reg0 <= 36'sb100001111110101100010110001000010000;
            sine_reg0   <= 36'sb1011000101001001000111100010100111;
        end
        7271: begin
            cosine_reg0 <= 36'sb100001111110011010111100110010100001;
            sine_reg0   <= 36'sb1011000100011001111101010110000110;
        end
        7272: begin
            cosine_reg0 <= 36'sb100001111110001001100100100110110111;
            sine_reg0   <= 36'sb1011000011101010110010101110010001;
        end
        7273: begin
            cosine_reg0 <= 36'sb100001111101111000001101100101010011;
            sine_reg0   <= 36'sb1011000010111011100111101011001001;
        end
        7274: begin
            cosine_reg0 <= 36'sb100001111101100110110111101101110110;
            sine_reg0   <= 36'sb1011000010001100011100001100110010;
        end
        7275: begin
            cosine_reg0 <= 36'sb100001111101010101100011000000100000;
            sine_reg0   <= 36'sb1011000001011101010000010011001100;
        end
        7276: begin
            cosine_reg0 <= 36'sb100001111101000100001111011101010010;
            sine_reg0   <= 36'sb1011000000101110000011111110011001;
        end
        7277: begin
            cosine_reg0 <= 36'sb100001111100110010111101000100001100;
            sine_reg0   <= 36'sb1010111111111110110111001110011011;
        end
        7278: begin
            cosine_reg0 <= 36'sb100001111100100001101011110101010000;
            sine_reg0   <= 36'sb1010111111001111101010000011010100;
        end
        7279: begin
            cosine_reg0 <= 36'sb100001111100010000011011110000011110;
            sine_reg0   <= 36'sb1010111110100000011100011101000111;
        end
        7280: begin
            cosine_reg0 <= 36'sb100001111011111111001100110101110111;
            sine_reg0   <= 36'sb1010111101110001001110011011110011;
        end
        7281: begin
            cosine_reg0 <= 36'sb100001111011101101111111000101011010;
            sine_reg0   <= 36'sb1010111101000001111111111111011101;
        end
        7282: begin
            cosine_reg0 <= 36'sb100001111011011100110010011111001010;
            sine_reg0   <= 36'sb1010111100010010110001001000000100;
        end
        7283: begin
            cosine_reg0 <= 36'sb100001111011001011100111000011000111;
            sine_reg0   <= 36'sb1010111011100011100001110101101100;
        end
        7284: begin
            cosine_reg0 <= 36'sb100001111010111010011100110001010001;
            sine_reg0   <= 36'sb1010111010110100010010001000010110;
        end
        7285: begin
            cosine_reg0 <= 36'sb100001111010101001010011101001101000;
            sine_reg0   <= 36'sb1010111010000101000010000000000011;
        end
        7286: begin
            cosine_reg0 <= 36'sb100001111010011000001011101100001111;
            sine_reg0   <= 36'sb1010111001010101110001011100110110;
        end
        7287: begin
            cosine_reg0 <= 36'sb100001111010000111000100111001000100;
            sine_reg0   <= 36'sb1010111000100110100000011110110000;
        end
        7288: begin
            cosine_reg0 <= 36'sb100001111001110101111111010000001010;
            sine_reg0   <= 36'sb1010110111110111001111000101110011;
        end
        7289: begin
            cosine_reg0 <= 36'sb100001111001100100111010110001100000;
            sine_reg0   <= 36'sb1010110111000111111101010010000010;
        end
        7290: begin
            cosine_reg0 <= 36'sb100001111001010011110111011101000111;
            sine_reg0   <= 36'sb1010110110011000101011000011011101;
        end
        7291: begin
            cosine_reg0 <= 36'sb100001111001000010110101010011000001;
            sine_reg0   <= 36'sb1010110101101001011000011010000111;
        end
        7292: begin
            cosine_reg0 <= 36'sb100001111000110001110100010011001101;
            sine_reg0   <= 36'sb1010110100111010000101010110000010;
        end
        7293: begin
            cosine_reg0 <= 36'sb100001111000100000110100011101101100;
            sine_reg0   <= 36'sb1010110100001010110001110111001110;
        end
        7294: begin
            cosine_reg0 <= 36'sb100001111000001111110101110010011111;
            sine_reg0   <= 36'sb1010110011011011011101111101101111;
        end
        7295: begin
            cosine_reg0 <= 36'sb100001110111111110111000010001100111;
            sine_reg0   <= 36'sb1010110010101100001001101001100110;
        end
        7296: begin
            cosine_reg0 <= 36'sb100001110111101101111011111011000011;
            sine_reg0   <= 36'sb1010110001111100110100111010110101;
        end
        7297: begin
            cosine_reg0 <= 36'sb100001110111011101000000101110110110;
            sine_reg0   <= 36'sb1010110001001101011111110001011101;
        end
        7298: begin
            cosine_reg0 <= 36'sb100001110111001100000110101100111111;
            sine_reg0   <= 36'sb1010110000011110001010001101100001;
        end
        7299: begin
            cosine_reg0 <= 36'sb100001110110111011001101110101011111;
            sine_reg0   <= 36'sb1010101111101110110100001111000010;
        end
        7300: begin
            cosine_reg0 <= 36'sb100001110110101010010110001000010111;
            sine_reg0   <= 36'sb1010101110111111011101110110000010;
        end
        7301: begin
            cosine_reg0 <= 36'sb100001110110011001011111100101101000;
            sine_reg0   <= 36'sb1010101110010000000111000010100011;
        end
        7302: begin
            cosine_reg0 <= 36'sb100001110110001000101010001101010010;
            sine_reg0   <= 36'sb1010101101100000101111110100100111;
        end
        7303: begin
            cosine_reg0 <= 36'sb100001110101110111110101111111010101;
            sine_reg0   <= 36'sb1010101100110001011000001100001111;
        end
        7304: begin
            cosine_reg0 <= 36'sb100001110101100111000010111011110011;
            sine_reg0   <= 36'sb1010101100000010000000001001011110;
        end
        7305: begin
            cosine_reg0 <= 36'sb100001110101010110010001000010101011;
            sine_reg0   <= 36'sb1010101011010010100111101100010101;
        end
        7306: begin
            cosine_reg0 <= 36'sb100001110101000101100000010100000000;
            sine_reg0   <= 36'sb1010101010100011001110110100110110;
        end
        7307: begin
            cosine_reg0 <= 36'sb100001110100110100110000101111110001;
            sine_reg0   <= 36'sb1010101001110011110101100011000011;
        end
        7308: begin
            cosine_reg0 <= 36'sb100001110100100100000010010101111111;
            sine_reg0   <= 36'sb1010101001000100011011110110111110;
        end
        7309: begin
            cosine_reg0 <= 36'sb100001110100010011010101000110101010;
            sine_reg0   <= 36'sb1010101000010101000001110000101000;
        end
        7310: begin
            cosine_reg0 <= 36'sb100001110100000010101001000001110100;
            sine_reg0   <= 36'sb1010100111100101100111010000000011;
        end
        7311: begin
            cosine_reg0 <= 36'sb100001110011110001111110000111011101;
            sine_reg0   <= 36'sb1010100110110110001100010101010010;
        end
        7312: begin
            cosine_reg0 <= 36'sb100001110011100001010100010111100101;
            sine_reg0   <= 36'sb1010100110000110110001000000010110;
        end
        7313: begin
            cosine_reg0 <= 36'sb100001110011010000101011110010001101;
            sine_reg0   <= 36'sb1010100101010111010101010001010000;
        end
        7314: begin
            cosine_reg0 <= 36'sb100001110011000000000100010111010110;
            sine_reg0   <= 36'sb1010100100100111111001001000000011;
        end
        7315: begin
            cosine_reg0 <= 36'sb100001110010101111011110000111000001;
            sine_reg0   <= 36'sb1010100011111000011100100100110001;
        end
        7316: begin
            cosine_reg0 <= 36'sb100001110010011110111001000001001110;
            sine_reg0   <= 36'sb1010100011001000111111100111011011;
        end
        7317: begin
            cosine_reg0 <= 36'sb100001110010001110010101000101111110;
            sine_reg0   <= 36'sb1010100010011001100010010000000011;
        end
        7318: begin
            cosine_reg0 <= 36'sb100001110001111101110010010101010001;
            sine_reg0   <= 36'sb1010100001101010000100011110101011;
        end
        7319: begin
            cosine_reg0 <= 36'sb100001110001101101010000101111001000;
            sine_reg0   <= 36'sb1010100000111010100110010011010101;
        end
        7320: begin
            cosine_reg0 <= 36'sb100001110001011100110000010011100011;
            sine_reg0   <= 36'sb1010100000001011000111101110000011;
        end
        7321: begin
            cosine_reg0 <= 36'sb100001110001001100010001000010100101;
            sine_reg0   <= 36'sb1010011111011011101000101110110110;
        end
        7322: begin
            cosine_reg0 <= 36'sb100001110000111011110010111100001100;
            sine_reg0   <= 36'sb1010011110101100001001010101110000;
        end
        7323: begin
            cosine_reg0 <= 36'sb100001110000101011010110000000011001;
            sine_reg0   <= 36'sb1010011101111100101001100010110100;
        end
        7324: begin
            cosine_reg0 <= 36'sb100001110000011010111010001111001110;
            sine_reg0   <= 36'sb1010011101001101001001010110000010;
        end
        7325: begin
            cosine_reg0 <= 36'sb100001110000001010011111101000101011;
            sine_reg0   <= 36'sb1010011100011101101000101111011110;
        end
        7326: begin
            cosine_reg0 <= 36'sb100001101111111010000110001100110000;
            sine_reg0   <= 36'sb1010011011101110000111101111001000;
        end
        7327: begin
            cosine_reg0 <= 36'sb100001101111101001101101111011011110;
            sine_reg0   <= 36'sb1010011010111110100110010101000010;
        end
        7328: begin
            cosine_reg0 <= 36'sb100001101111011001010110110100110110;
            sine_reg0   <= 36'sb1010011010001111000100100001001111;
        end
        7329: begin
            cosine_reg0 <= 36'sb100001101111001001000000111000111000;
            sine_reg0   <= 36'sb1010011001011111100010010011110000;
        end
        7330: begin
            cosine_reg0 <= 36'sb100001101110111000101100000111100110;
            sine_reg0   <= 36'sb1010011000101111111111101100100110;
        end
        7331: begin
            cosine_reg0 <= 36'sb100001101110101000011000100000111111;
            sine_reg0   <= 36'sb1010011000000000011100101011110101;
        end
        7332: begin
            cosine_reg0 <= 36'sb100001101110011000000110000101000100;
            sine_reg0   <= 36'sb1010010111010000111001010001011101;
        end
        7333: begin
            cosine_reg0 <= 36'sb100001101110000111110100110011110110;
            sine_reg0   <= 36'sb1010010110100001010101011101100001;
        end
        7334: begin
            cosine_reg0 <= 36'sb100001101101110111100100101101010110;
            sine_reg0   <= 36'sb1010010101110001110001010000000010;
        end
        7335: begin
            cosine_reg0 <= 36'sb100001101101100111010101110001100100;
            sine_reg0   <= 36'sb1010010101000010001100101001000010;
        end
        7336: begin
            cosine_reg0 <= 36'sb100001101101010111001000000000100000;
            sine_reg0   <= 36'sb1010010100010010100111101000100011;
        end
        7337: begin
            cosine_reg0 <= 36'sb100001101101000110111011011010001101;
            sine_reg0   <= 36'sb1010010011100011000010001110100111;
        end
        7338: begin
            cosine_reg0 <= 36'sb100001101100110110101111111110101001;
            sine_reg0   <= 36'sb1010010010110011011100011011001111;
        end
        7339: begin
            cosine_reg0 <= 36'sb100001101100100110100101101101110101;
            sine_reg0   <= 36'sb1010010010000011110110001110011110;
        end
        7340: begin
            cosine_reg0 <= 36'sb100001101100010110011100100111110011;
            sine_reg0   <= 36'sb1010010001010100001111101000010110;
        end
        7341: begin
            cosine_reg0 <= 36'sb100001101100000110010100101100100011;
            sine_reg0   <= 36'sb1010010000100100101000101000110111;
        end
        7342: begin
            cosine_reg0 <= 36'sb100001101011110110001101111100000110;
            sine_reg0   <= 36'sb1010001111110101000001010000000101;
        end
        7343: begin
            cosine_reg0 <= 36'sb100001101011100110001000010110011011;
            sine_reg0   <= 36'sb1010001111000101011001011110000000;
        end
        7344: begin
            cosine_reg0 <= 36'sb100001101011010110000011111011100100;
            sine_reg0   <= 36'sb1010001110010101110001010010101011;
        end
        7345: begin
            cosine_reg0 <= 36'sb100001101011000110000000101011100010;
            sine_reg0   <= 36'sb1010001101100110001000101110000111;
        end
        7346: begin
            cosine_reg0 <= 36'sb100001101010110101111110100110010101;
            sine_reg0   <= 36'sb1010001100110110011111110000010111;
        end
        7347: begin
            cosine_reg0 <= 36'sb100001101010100101111101101011111101;
            sine_reg0   <= 36'sb1010001100000110110110011001011011;
        end
        7348: begin
            cosine_reg0 <= 36'sb100001101010010101111101111100011011;
            sine_reg0   <= 36'sb1010001011010111001100101001010111;
        end
        7349: begin
            cosine_reg0 <= 36'sb100001101010000101111111010111110001;
            sine_reg0   <= 36'sb1010001010100111100010100000001100;
        end
        7350: begin
            cosine_reg0 <= 36'sb100001101001110110000001111101111101;
            sine_reg0   <= 36'sb1010001001110111110111111101111011;
        end
        7351: begin
            cosine_reg0 <= 36'sb100001101001100110000101101111000010;
            sine_reg0   <= 36'sb1010001001001000001101000010100111;
        end
        7352: begin
            cosine_reg0 <= 36'sb100001101001010110001010101011000000;
            sine_reg0   <= 36'sb1010001000011000100001101110010001;
        end
        7353: begin
            cosine_reg0 <= 36'sb100001101001000110010000110001110111;
            sine_reg0   <= 36'sb1010000111101000110110000000111011;
        end
        7354: begin
            cosine_reg0 <= 36'sb100001101000110110011000000011100111;
            sine_reg0   <= 36'sb1010000110111001001001111010100111;
        end
        7355: begin
            cosine_reg0 <= 36'sb100001101000100110100000100000010011;
            sine_reg0   <= 36'sb1010000110001001011101011011011000;
        end
        7356: begin
            cosine_reg0 <= 36'sb100001101000010110101010000111111001;
            sine_reg0   <= 36'sb1010000101011001110000100011001101;
        end
        7357: begin
            cosine_reg0 <= 36'sb100001101000000110110100111010011011;
            sine_reg0   <= 36'sb1010000100101010000011010010001011;
        end
        7358: begin
            cosine_reg0 <= 36'sb100001100111110111000000110111111010;
            sine_reg0   <= 36'sb1010000011111010010101101000010010;
        end
        7359: begin
            cosine_reg0 <= 36'sb100001100111100111001110000000010110;
            sine_reg0   <= 36'sb1010000011001010100111100101100100;
        end
        7360: begin
            cosine_reg0 <= 36'sb100001100111010111011100010011101111;
            sine_reg0   <= 36'sb1010000010011010111001001010000011;
        end
        7361: begin
            cosine_reg0 <= 36'sb100001100111000111101011110010000110;
            sine_reg0   <= 36'sb1010000001101011001010010101110001;
        end
        7362: begin
            cosine_reg0 <= 36'sb100001100110110111111100011011011100;
            sine_reg0   <= 36'sb1010000000111011011011001000101111;
        end
        7363: begin
            cosine_reg0 <= 36'sb100001100110101000001110001111110010;
            sine_reg0   <= 36'sb1010000000001011101011100011000000;
        end
        7364: begin
            cosine_reg0 <= 36'sb100001100110011000100001001111000111;
            sine_reg0   <= 36'sb1001111111011011111011100100100110;
        end
        7365: begin
            cosine_reg0 <= 36'sb100001100110001000110101011001011101;
            sine_reg0   <= 36'sb1001111110101100001011001101100010;
        end
        7366: begin
            cosine_reg0 <= 36'sb100001100101111001001010101110110101;
            sine_reg0   <= 36'sb1001111101111100011010011101110110;
        end
        7367: begin
            cosine_reg0 <= 36'sb100001100101101001100001001111001110;
            sine_reg0   <= 36'sb1001111101001100101001010101100100;
        end
        7368: begin
            cosine_reg0 <= 36'sb100001100101011001111000111010101010;
            sine_reg0   <= 36'sb1001111100011100110111110100101110;
        end
        7369: begin
            cosine_reg0 <= 36'sb100001100101001010010001110001001000;
            sine_reg0   <= 36'sb1001111011101101000101111011010101;
        end
        7370: begin
            cosine_reg0 <= 36'sb100001100100111010101011110010101011;
            sine_reg0   <= 36'sb1001111010111101010011101001011100;
        end
        7371: begin
            cosine_reg0 <= 36'sb100001100100101011000110111111010001;
            sine_reg0   <= 36'sb1001111010001101100000111111000100;
        end
        7372: begin
            cosine_reg0 <= 36'sb100001100100011011100011010110111100;
            sine_reg0   <= 36'sb1001111001011101101101111100001111;
        end
        7373: begin
            cosine_reg0 <= 36'sb100001100100001100000000111001101101;
            sine_reg0   <= 36'sb1001111000101101111010100000111111;
        end
        7374: begin
            cosine_reg0 <= 36'sb100001100011111100011111100111100100;
            sine_reg0   <= 36'sb1001110111111110000110101101010110;
        end
        7375: begin
            cosine_reg0 <= 36'sb100001100011101100111111100000100010;
            sine_reg0   <= 36'sb1001110111001110010010100001010110;
        end
        7376: begin
            cosine_reg0 <= 36'sb100001100011011101100000100100100110;
            sine_reg0   <= 36'sb1001110110011110011101111101000000;
        end
        7377: begin
            cosine_reg0 <= 36'sb100001100011001110000010110011110011;
            sine_reg0   <= 36'sb1001110101101110101001000000010111;
        end
        7378: begin
            cosine_reg0 <= 36'sb100001100010111110100110001110001000;
            sine_reg0   <= 36'sb1001110100111110110011101011011100;
        end
        7379: begin
            cosine_reg0 <= 36'sb100001100010101111001010110011100110;
            sine_reg0   <= 36'sb1001110100001110111101111110010000;
        end
        7380: begin
            cosine_reg0 <= 36'sb100001100010011111110000100100001101;
            sine_reg0   <= 36'sb1001110011011111000111111000110111;
        end
        7381: begin
            cosine_reg0 <= 36'sb100001100010010000010111011111111111;
            sine_reg0   <= 36'sb1001110010101111010001011011010010;
        end
        7382: begin
            cosine_reg0 <= 36'sb100001100010000000111111100110111100;
            sine_reg0   <= 36'sb1001110001111111011010100101100010;
        end
        7383: begin
            cosine_reg0 <= 36'sb100001100001110001101000111001000100;
            sine_reg0   <= 36'sb1001110001001111100011010111101001;
        end
        7384: begin
            cosine_reg0 <= 36'sb100001100001100010010011010110011000;
            sine_reg0   <= 36'sb1001110000011111101011110001101010;
        end
        7385: begin
            cosine_reg0 <= 36'sb100001100001010010111110111110111000;
            sine_reg0   <= 36'sb1001101111101111110011110011100110;
        end
        7386: begin
            cosine_reg0 <= 36'sb100001100001000011101011110010100110;
            sine_reg0   <= 36'sb1001101110111111111011011101011111;
        end
        7387: begin
            cosine_reg0 <= 36'sb100001100000110100011001110001100001;
            sine_reg0   <= 36'sb1001101110010000000010101111010111;
        end
        7388: begin
            cosine_reg0 <= 36'sb100001100000100101001000111011101011;
            sine_reg0   <= 36'sb1001101101100000001001101001001111;
        end
        7389: begin
            cosine_reg0 <= 36'sb100001100000010101111001010001000100;
            sine_reg0   <= 36'sb1001101100110000010000001011001010;
        end
        7390: begin
            cosine_reg0 <= 36'sb100001100000000110101010110001101100;
            sine_reg0   <= 36'sb1001101100000000010110010101001001;
        end
        7391: begin
            cosine_reg0 <= 36'sb100001011111110111011101011101100101;
            sine_reg0   <= 36'sb1001101011010000011100000111001110;
        end
        7392: begin
            cosine_reg0 <= 36'sb100001011111101000010001010100101110;
            sine_reg0   <= 36'sb1001101010100000100001100001011100;
        end
        7393: begin
            cosine_reg0 <= 36'sb100001011111011001000110010111001000;
            sine_reg0   <= 36'sb1001101001110000100110100011110011;
        end
        7394: begin
            cosine_reg0 <= 36'sb100001011111001001111100100100110100;
            sine_reg0   <= 36'sb1001101001000000101011001110010110;
        end
        7395: begin
            cosine_reg0 <= 36'sb100001011110111010110011111101110011;
            sine_reg0   <= 36'sb1001101000010000101111100001000111;
        end
        7396: begin
            cosine_reg0 <= 36'sb100001011110101011101100100010000101;
            sine_reg0   <= 36'sb1001100111100000110011011100000111;
        end
        7397: begin
            cosine_reg0 <= 36'sb100001011110011100100110010001101010;
            sine_reg0   <= 36'sb1001100110110000110110111111011000;
        end
        7398: begin
            cosine_reg0 <= 36'sb100001011110001101100001001100100100;
            sine_reg0   <= 36'sb1001100110000000111010001010111101;
        end
        7399: begin
            cosine_reg0 <= 36'sb100001011101111110011101010010110010;
            sine_reg0   <= 36'sb1001100101010000111100111110110110;
        end
        7400: begin
            cosine_reg0 <= 36'sb100001011101101111011010100100010110;
            sine_reg0   <= 36'sb1001100100100000111111011011000111;
        end
        7401: begin
            cosine_reg0 <= 36'sb100001011101100000011001000001001111;
            sine_reg0   <= 36'sb1001100011110001000001011111110000;
        end
        7402: begin
            cosine_reg0 <= 36'sb100001011101010001011000101001011111;
            sine_reg0   <= 36'sb1001100011000001000011001100110011;
        end
        7403: begin
            cosine_reg0 <= 36'sb100001011101000010011001011101000111;
            sine_reg0   <= 36'sb1001100010010001000100100010010011;
        end
        7404: begin
            cosine_reg0 <= 36'sb100001011100110011011011011100000110;
            sine_reg0   <= 36'sb1001100001100001000101100000010001;
        end
        7405: begin
            cosine_reg0 <= 36'sb100001011100100100011110100110011101;
            sine_reg0   <= 36'sb1001100000110001000110000110110000;
        end
        7406: begin
            cosine_reg0 <= 36'sb100001011100010101100010111100001101;
            sine_reg0   <= 36'sb1001100000000001000110010101110000;
        end
        7407: begin
            cosine_reg0 <= 36'sb100001011100000110101000011101010110;
            sine_reg0   <= 36'sb1001011111010001000110001101010100;
        end
        7408: begin
            cosine_reg0 <= 36'sb100001011011110111101111001001111001;
            sine_reg0   <= 36'sb1001011110100001000101101101011101;
        end
        7409: begin
            cosine_reg0 <= 36'sb100001011011101000110111000001110111;
            sine_reg0   <= 36'sb1001011101110001000100110110001110;
        end
        7410: begin
            cosine_reg0 <= 36'sb100001011011011010000000000101010000;
            sine_reg0   <= 36'sb1001011101000001000011100111101001;
        end
        7411: begin
            cosine_reg0 <= 36'sb100001011011001011001010010100000101;
            sine_reg0   <= 36'sb1001011100010001000010000001101110;
        end
        7412: begin
            cosine_reg0 <= 36'sb100001011010111100010101101110010110;
            sine_reg0   <= 36'sb1001011011100001000000000100100001;
        end
        7413: begin
            cosine_reg0 <= 36'sb100001011010101101100010010100000100;
            sine_reg0   <= 36'sb1001011010110000111101110000000010;
        end
        7414: begin
            cosine_reg0 <= 36'sb100001011010011110110000000101001111;
            sine_reg0   <= 36'sb1001011010000000111011000100010100;
        end
        7415: begin
            cosine_reg0 <= 36'sb100001011010001111111111000001111001;
            sine_reg0   <= 36'sb1001011001010000111000000001011001;
        end
        7416: begin
            cosine_reg0 <= 36'sb100001011010000001001111001010000001;
            sine_reg0   <= 36'sb1001011000100000110100100111010010;
        end
        7417: begin
            cosine_reg0 <= 36'sb100001011001110010100000011101101000;
            sine_reg0   <= 36'sb1001010111110000110000110110000010;
        end
        7418: begin
            cosine_reg0 <= 36'sb100001011001100011110010111100101110;
            sine_reg0   <= 36'sb1001010111000000101100101101101010;
        end
        7419: begin
            cosine_reg0 <= 36'sb100001011001010101000110100111010101;
            sine_reg0   <= 36'sb1001010110010000101000001110001011;
        end
        7420: begin
            cosine_reg0 <= 36'sb100001011001000110011011011101011101;
            sine_reg0   <= 36'sb1001010101100000100011010111101001;
        end
        7421: begin
            cosine_reg0 <= 36'sb100001011000110111110001011111000110;
            sine_reg0   <= 36'sb1001010100110000011110001010000100;
        end
        7422: begin
            cosine_reg0 <= 36'sb100001011000101001001000101100010001;
            sine_reg0   <= 36'sb1001010100000000011000100101011111;
        end
        7423: begin
            cosine_reg0 <= 36'sb100001011000011010100001000100111111;
            sine_reg0   <= 36'sb1001010011010000010010101001111011;
        end
        7424: begin
            cosine_reg0 <= 36'sb100001011000001011111010101001001111;
            sine_reg0   <= 36'sb1001010010100000001100010111011010;
        end
        7425: begin
            cosine_reg0 <= 36'sb100001010111111101010101011001000100;
            sine_reg0   <= 36'sb1001010001110000000101101101111111;
        end
        7426: begin
            cosine_reg0 <= 36'sb100001010111101110110001010100011100;
            sine_reg0   <= 36'sb1001010000111111111110101101101011;
        end
        7427: begin
            cosine_reg0 <= 36'sb100001010111100000001110011011011010;
            sine_reg0   <= 36'sb1001010000001111110111010110011111;
        end
        7428: begin
            cosine_reg0 <= 36'sb100001010111010001101100101101111100;
            sine_reg0   <= 36'sb1001001111011111101111101000011110;
        end
        7429: begin
            cosine_reg0 <= 36'sb100001010111000011001100001100000101;
            sine_reg0   <= 36'sb1001001110101111100111100011101010;
        end
        7430: begin
            cosine_reg0 <= 36'sb100001010110110100101100110101110100;
            sine_reg0   <= 36'sb1001001101111111011111001000000100;
        end
        7431: begin
            cosine_reg0 <= 36'sb100001010110100110001110101011001010;
            sine_reg0   <= 36'sb1001001101001111010110010101101110;
        end
        7432: begin
            cosine_reg0 <= 36'sb100001010110010111110001101100000111;
            sine_reg0   <= 36'sb1001001100011111001101001100101010;
        end
        7433: begin
            cosine_reg0 <= 36'sb100001010110001001010101111000101101;
            sine_reg0   <= 36'sb1001001011101111000011101100111011;
        end
        7434: begin
            cosine_reg0 <= 36'sb100001010101111010111011010000111011;
            sine_reg0   <= 36'sb1001001010111110111001110110100001;
        end
        7435: begin
            cosine_reg0 <= 36'sb100001010101101100100001110100110011;
            sine_reg0   <= 36'sb1001001010001110101111101001011111;
        end
        7436: begin
            cosine_reg0 <= 36'sb100001010101011110001001100100010100;
            sine_reg0   <= 36'sb1001001001011110100101000101110110;
        end
        7437: begin
            cosine_reg0 <= 36'sb100001010101001111110010011111100000;
            sine_reg0   <= 36'sb1001001000101110011010001011101001;
        end
        7438: begin
            cosine_reg0 <= 36'sb100001010101000001011100100110010111;
            sine_reg0   <= 36'sb1001000111111110001110111010111001;
        end
        7439: begin
            cosine_reg0 <= 36'sb100001010100110011000111111000111001;
            sine_reg0   <= 36'sb1001000111001110000011010011101000;
        end
        7440: begin
            cosine_reg0 <= 36'sb100001010100100100110100010111000111;
            sine_reg0   <= 36'sb1001000110011101110111010101111000;
        end
        7441: begin
            cosine_reg0 <= 36'sb100001010100010110100010000001000010;
            sine_reg0   <= 36'sb1001000101101101101011000001101011;
        end
        7442: begin
            cosine_reg0 <= 36'sb100001010100001000010000110110101001;
            sine_reg0   <= 36'sb1001000100111101011110010111000011;
        end
        7443: begin
            cosine_reg0 <= 36'sb100001010011111010000000110111111111;
            sine_reg0   <= 36'sb1001000100001101010001010110000001;
        end
        7444: begin
            cosine_reg0 <= 36'sb100001010011101011110010000101000011;
            sine_reg0   <= 36'sb1001000011011101000011111110100111;
        end
        7445: begin
            cosine_reg0 <= 36'sb100001010011011101100100011101110101;
            sine_reg0   <= 36'sb1001000010101100110110010000111000;
        end
        7446: begin
            cosine_reg0 <= 36'sb100001010011001111011000000010010111;
            sine_reg0   <= 36'sb1001000001111100101000001100110101;
        end
        7447: begin
            cosine_reg0 <= 36'sb100001010011000001001100110010101000;
            sine_reg0   <= 36'sb1001000001001100011001110010100000;
        end
        7448: begin
            cosine_reg0 <= 36'sb100001010010110011000010101110101010;
            sine_reg0   <= 36'sb1001000000011100001011000001111011;
        end
        7449: begin
            cosine_reg0 <= 36'sb100001010010100100111001110110011101;
            sine_reg0   <= 36'sb1000111111101011111011111011000111;
        end
        7450: begin
            cosine_reg0 <= 36'sb100001010010010110110010001010000001;
            sine_reg0   <= 36'sb1000111110111011101100011110000111;
        end
        7451: begin
            cosine_reg0 <= 36'sb100001010010001000101011101001011000;
            sine_reg0   <= 36'sb1000111110001011011100101010111100;
        end
        7452: begin
            cosine_reg0 <= 36'sb100001010001111010100110010100100001;
            sine_reg0   <= 36'sb1000111101011011001100100001101001;
        end
        7453: begin
            cosine_reg0 <= 36'sb100001010001101100100010001011011101;
            sine_reg0   <= 36'sb1000111100101010111100000010001111;
        end
        7454: begin
            cosine_reg0 <= 36'sb100001010001011110011111001110001101;
            sine_reg0   <= 36'sb1000111011111010101011001100101111;
        end
        7455: begin
            cosine_reg0 <= 36'sb100001010001010000011101011100110000;
            sine_reg0   <= 36'sb1000111011001010011010000001001101;
        end
        7456: begin
            cosine_reg0 <= 36'sb100001010001000010011100110111001001;
            sine_reg0   <= 36'sb1000111010011010001000011111101001;
        end
        7457: begin
            cosine_reg0 <= 36'sb100001010000110100011101011101010111;
            sine_reg0   <= 36'sb1000111001101001110110101000000110;
        end
        7458: begin
            cosine_reg0 <= 36'sb100001010000100110011111001111011011;
            sine_reg0   <= 36'sb1000111000111001100100011010100110;
        end
        7459: begin
            cosine_reg0 <= 36'sb100001010000011000100010001101010101;
            sine_reg0   <= 36'sb1000111000001001010001110111001001;
        end
        7460: begin
            cosine_reg0 <= 36'sb100001010000001010100110010111000110;
            sine_reg0   <= 36'sb1000110111011000111110111101110011;
        end
        7461: begin
            cosine_reg0 <= 36'sb100001001111111100101011101100101111;
            sine_reg0   <= 36'sb1000110110101000101011101110100101;
        end
        7462: begin
            cosine_reg0 <= 36'sb100001001111101110110010001110001111;
            sine_reg0   <= 36'sb1000110101111000011000001001100000;
        end
        7463: begin
            cosine_reg0 <= 36'sb100001001111100000111001111011101000;
            sine_reg0   <= 36'sb1000110101001000000100001110101000;
        end
        7464: begin
            cosine_reg0 <= 36'sb100001001111010011000010110100111010;
            sine_reg0   <= 36'sb1000110100010111101111111101111101;
        end
        7465: begin
            cosine_reg0 <= 36'sb100001001111000101001100111010000110;
            sine_reg0   <= 36'sb1000110011100111011011010111100001;
        end
        7466: begin
            cosine_reg0 <= 36'sb100001001110110111011000001011001100;
            sine_reg0   <= 36'sb1000110010110111000110011011010111;
        end
        7467: begin
            cosine_reg0 <= 36'sb100001001110101001100100101000001100;
            sine_reg0   <= 36'sb1000110010000110110001001001100000;
        end
        7468: begin
            cosine_reg0 <= 36'sb100001001110011011110010010001000111;
            sine_reg0   <= 36'sb1000110001010110011011100001111110;
        end
        7469: begin
            cosine_reg0 <= 36'sb100001001110001110000001000101111111;
            sine_reg0   <= 36'sb1000110000100110000101100100110011;
        end
        7470: begin
            cosine_reg0 <= 36'sb100001001110000000010001000110110010;
            sine_reg0   <= 36'sb1000101111110101101111010010000001;
        end
        7471: begin
            cosine_reg0 <= 36'sb100001001101110010100010010011100010;
            sine_reg0   <= 36'sb1000101111000101011000101001101010;
        end
        7472: begin
            cosine_reg0 <= 36'sb100001001101100100110100101100010000;
            sine_reg0   <= 36'sb1000101110010101000001101011101111;
        end
        7473: begin
            cosine_reg0 <= 36'sb100001001101010111001000010000111011;
            sine_reg0   <= 36'sb1000101101100100101010011000010010;
        end
        7474: begin
            cosine_reg0 <= 36'sb100001001101001001011101000001100101;
            sine_reg0   <= 36'sb1000101100110100010010101111010101;
        end
        7475: begin
            cosine_reg0 <= 36'sb100001001100111011110010111110001110;
            sine_reg0   <= 36'sb1000101100000011111010110000111011;
        end
        7476: begin
            cosine_reg0 <= 36'sb100001001100101110001010000110110110;
            sine_reg0   <= 36'sb1000101011010011100010011101000101;
        end
        7477: begin
            cosine_reg0 <= 36'sb100001001100100000100010011011011110;
            sine_reg0   <= 36'sb1000101010100011001001110011110100;
        end
        7478: begin
            cosine_reg0 <= 36'sb100001001100010010111011111100000110;
            sine_reg0   <= 36'sb1000101001110010110000110101001100;
        end
        7479: begin
            cosine_reg0 <= 36'sb100001001100000101010110101000110000;
            sine_reg0   <= 36'sb1000101001000010010111100001001100;
        end
        7480: begin
            cosine_reg0 <= 36'sb100001001011110111110010100001011011;
            sine_reg0   <= 36'sb1000101000010001111101110111111001;
        end
        7481: begin
            cosine_reg0 <= 36'sb100001001011101010001111100110001000;
            sine_reg0   <= 36'sb1000100111100001100011111001010010;
        end
        7482: begin
            cosine_reg0 <= 36'sb100001001011011100101101110110110111;
            sine_reg0   <= 36'sb1000100110110001001001100101011011;
        end
        7483: begin
            cosine_reg0 <= 36'sb100001001011001111001101010011101010;
            sine_reg0   <= 36'sb1000100110000000101110111100010100;
        end
        7484: begin
            cosine_reg0 <= 36'sb100001001011000001101101111100100000;
            sine_reg0   <= 36'sb1000100101010000010011111110000001;
        end
        7485: begin
            cosine_reg0 <= 36'sb100001001010110100001111110001011010;
            sine_reg0   <= 36'sb1000100100011111111000101010100011;
        end
        7486: begin
            cosine_reg0 <= 36'sb100001001010100110110010110010011001;
            sine_reg0   <= 36'sb1000100011101111011101000001111011;
        end
        7487: begin
            cosine_reg0 <= 36'sb100001001010011001010110111111011101;
            sine_reg0   <= 36'sb1000100010111111000001000100001011;
        end
        7488: begin
            cosine_reg0 <= 36'sb100001001010001011111100011000100111;
            sine_reg0   <= 36'sb1000100010001110100100110001010110;
        end
        7489: begin
            cosine_reg0 <= 36'sb100001001001111110100010111101110111;
            sine_reg0   <= 36'sb1000100001011110001000001001011101;
        end
        7490: begin
            cosine_reg0 <= 36'sb100001001001110001001010101111001101;
            sine_reg0   <= 36'sb1000100000101101101011001100100010;
        end
        7491: begin
            cosine_reg0 <= 36'sb100001001001100011110011101100101011;
            sine_reg0   <= 36'sb1000011111111101001101111010101000;
        end
        7492: begin
            cosine_reg0 <= 36'sb100001001001010110011101110110010001;
            sine_reg0   <= 36'sb1000011111001100110000010011101111;
        end
        7493: begin
            cosine_reg0 <= 36'sb100001001001001001001001001011111111;
            sine_reg0   <= 36'sb1000011110011100010010010111111001;
        end
        7494: begin
            cosine_reg0 <= 36'sb100001001000111011110101101101110101;
            sine_reg0   <= 36'sb1000011101101011110100000111001010;
        end
        7495: begin
            cosine_reg0 <= 36'sb100001001000101110100011011011110101;
            sine_reg0   <= 36'sb1000011100111011010101100001100010;
        end
        7496: begin
            cosine_reg0 <= 36'sb100001001000100001010010010101111111;
            sine_reg0   <= 36'sb1000011100001010110110100111000011;
        end
        7497: begin
            cosine_reg0 <= 36'sb100001001000010100000010011100010011;
            sine_reg0   <= 36'sb1000011011011010010111010111101111;
        end
        7498: begin
            cosine_reg0 <= 36'sb100001001000000110110011101110110010;
            sine_reg0   <= 36'sb1000011010101001110111110011101000;
        end
        7499: begin
            cosine_reg0 <= 36'sb100001000111111001100110001101011100;
            sine_reg0   <= 36'sb1000011001111001010111111010110001;
        end
        7500: begin
            cosine_reg0 <= 36'sb100001000111101100011001111000010010;
            sine_reg0   <= 36'sb1000011001001000110111101101001010;
        end
        7501: begin
            cosine_reg0 <= 36'sb100001000111011111001110101111010100;
            sine_reg0   <= 36'sb1000011000011000010111001010110101;
        end
        7502: begin
            cosine_reg0 <= 36'sb100001000111010010000100110010100011;
            sine_reg0   <= 36'sb1000010111100111110110010011110110;
        end
        7503: begin
            cosine_reg0 <= 36'sb100001000111000100111100000010000000;
            sine_reg0   <= 36'sb1000010110110111010101001000001100;
        end
        7504: begin
            cosine_reg0 <= 36'sb100001000110110111110100011101101010;
            sine_reg0   <= 36'sb1000010110000110110011100111111011;
        end
        7505: begin
            cosine_reg0 <= 36'sb100001000110101010101110000101100011;
            sine_reg0   <= 36'sb1000010101010110010001110011000100;
        end
        7506: begin
            cosine_reg0 <= 36'sb100001000110011101101000111001101011;
            sine_reg0   <= 36'sb1000010100100101101111101001101001;
        end
        7507: begin
            cosine_reg0 <= 36'sb100001000110010000100100111010000010;
            sine_reg0   <= 36'sb1000010011110101001101001011101100;
        end
        7508: begin
            cosine_reg0 <= 36'sb100001000110000011100010000110101001;
            sine_reg0   <= 36'sb1000010011000100101010011001001111;
        end
        7509: begin
            cosine_reg0 <= 36'sb100001000101110110100000011111100000;
            sine_reg0   <= 36'sb1000010010010100000111010010010100;
        end
        7510: begin
            cosine_reg0 <= 36'sb100001000101101001100000000100101000;
            sine_reg0   <= 36'sb1000010001100011100011110110111011;
        end
        7511: begin
            cosine_reg0 <= 36'sb100001000101011100100000110110000001;
            sine_reg0   <= 36'sb1000010000110011000000000111001001;
        end
        7512: begin
            cosine_reg0 <= 36'sb100001000101001111100010110011101101;
            sine_reg0   <= 36'sb1000010000000010011100000010111101;
        end
        7513: begin
            cosine_reg0 <= 36'sb100001000101000010100101111101101011;
            sine_reg0   <= 36'sb1000001111010001110111101010011011;
        end
        7514: begin
            cosine_reg0 <= 36'sb100001000100110101101010010011111011;
            sine_reg0   <= 36'sb1000001110100001010010111101100011;
        end
        7515: begin
            cosine_reg0 <= 36'sb100001000100101000101111110110011111;
            sine_reg0   <= 36'sb1000001101110000101101111100011001;
        end
        7516: begin
            cosine_reg0 <= 36'sb100001000100011011110110100101010111;
            sine_reg0   <= 36'sb1000001101000000001000100110111101;
        end
        7517: begin
            cosine_reg0 <= 36'sb100001000100001110111110100000100100;
            sine_reg0   <= 36'sb1000001100001111100010111101010010;
        end
        7518: begin
            cosine_reg0 <= 36'sb100001000100000010000111101000000101;
            sine_reg0   <= 36'sb1000001011011110111100111111011001;
        end
        7519: begin
            cosine_reg0 <= 36'sb100001000011110101010001111011111011;
            sine_reg0   <= 36'sb1000001010101110010110101101010101;
        end
        7520: begin
            cosine_reg0 <= 36'sb100001000011101000011101011100001000;
            sine_reg0   <= 36'sb1000001001111101110000000111000111;
        end
        7521: begin
            cosine_reg0 <= 36'sb100001000011011011101010001000101011;
            sine_reg0   <= 36'sb1000001001001101001001001100110001;
        end
        7522: begin
            cosine_reg0 <= 36'sb100001000011001110111000000001100100;
            sine_reg0   <= 36'sb1000001000011100100001111110010101;
        end
        7523: begin
            cosine_reg0 <= 36'sb100001000011000010000111000110110101;
            sine_reg0   <= 36'sb1000000111101011111010011011110101;
        end
        7524: begin
            cosine_reg0 <= 36'sb100001000010110101010111011000011110;
            sine_reg0   <= 36'sb1000000110111011010010100101010010;
        end
        7525: begin
            cosine_reg0 <= 36'sb100001000010101000101000110110011111;
            sine_reg0   <= 36'sb1000000110001010101010011010101111;
        end
        7526: begin
            cosine_reg0 <= 36'sb100001000010011011111011100000111001;
            sine_reg0   <= 36'sb1000000101011010000001111100001110;
        end
        7527: begin
            cosine_reg0 <= 36'sb100001000010001111001111010111101101;
            sine_reg0   <= 36'sb1000000100101001011001001001110000;
        end
        7528: begin
            cosine_reg0 <= 36'sb100001000010000010100100011010111010;
            sine_reg0   <= 36'sb1000000011111000110000000011010111;
        end
        7529: begin
            cosine_reg0 <= 36'sb100001000001110101111010101010100001;
            sine_reg0   <= 36'sb1000000011001000000110101001000101;
        end
        7530: begin
            cosine_reg0 <= 36'sb100001000001101001010010000110100011;
            sine_reg0   <= 36'sb1000000010010111011100111010111101;
        end
        7531: begin
            cosine_reg0 <= 36'sb100001000001011100101010101111000001;
            sine_reg0   <= 36'sb1000000001100110110010111000111111;
        end
        7532: begin
            cosine_reg0 <= 36'sb100001000001010000000100100011111010;
            sine_reg0   <= 36'sb1000000000110110001000100011001110;
        end
        7533: begin
            cosine_reg0 <= 36'sb100001000001000011011111100101001111;
            sine_reg0   <= 36'sb1000000000000101011101111001101011;
        end
        7534: begin
            cosine_reg0 <= 36'sb100001000000110110111011110011000010;
            sine_reg0   <= 36'sb111111111010100110010111100011001;
        end
        7535: begin
            cosine_reg0 <= 36'sb100001000000101010011001001101010001;
            sine_reg0   <= 36'sb111111110100100000111101011011001;
        end
        7536: begin
            cosine_reg0 <= 36'sb100001000000011101110111110011111110;
            sine_reg0   <= 36'sb111111101110011011100000110101110;
        end
        7537: begin
            cosine_reg0 <= 36'sb100001000000010001010111100111001001;
            sine_reg0   <= 36'sb111111101000010110000001110011000;
        end
        7538: begin
            cosine_reg0 <= 36'sb100001000000000100111000100110110011;
            sine_reg0   <= 36'sb111111100010010000100000010011011;
        end
        7539: begin
            cosine_reg0 <= 36'sb100000111111111000011010110010111100;
            sine_reg0   <= 36'sb111111011100001010111100010110111;
        end
        7540: begin
            cosine_reg0 <= 36'sb100000111111101011111110001011100101;
            sine_reg0   <= 36'sb111111010110000101010101111110000;
        end
        7541: begin
            cosine_reg0 <= 36'sb100000111111011111100010110000101110;
            sine_reg0   <= 36'sb111111001111111111101101001000110;
        end
        7542: begin
            cosine_reg0 <= 36'sb100000111111010011001000100010010111;
            sine_reg0   <= 36'sb111111001001111010000001110111011;
        end
        7543: begin
            cosine_reg0 <= 36'sb100000111111000110101111100000100001;
            sine_reg0   <= 36'sb111111000011110100010100001010010;
        end
        7544: begin
            cosine_reg0 <= 36'sb100000111110111010010111101011001101;
            sine_reg0   <= 36'sb111110111101101110100100000001100;
        end
        7545: begin
            cosine_reg0 <= 36'sb100000111110101110000001000010011011;
            sine_reg0   <= 36'sb111110110111101000110001011101011;
        end
        7546: begin
            cosine_reg0 <= 36'sb100000111110100001101011100110001011;
            sine_reg0   <= 36'sb111110110001100010111100011110001;
        end
        7547: begin
            cosine_reg0 <= 36'sb100000111110010101010111010110011111;
            sine_reg0   <= 36'sb111110101011011101000101000100000;
        end
        7548: begin
            cosine_reg0 <= 36'sb100000111110001001000100010011010101;
            sine_reg0   <= 36'sb111110100101010111001011001111010;
        end
        7549: begin
            cosine_reg0 <= 36'sb100000111101111100110010011100110000;
            sine_reg0   <= 36'sb111110011111010001001111000000000;
        end
        7550: begin
            cosine_reg0 <= 36'sb100000111101110000100001110010101111;
            sine_reg0   <= 36'sb111110011001001011010000010110101;
        end
        7551: begin
            cosine_reg0 <= 36'sb100000111101100100010010010101010011;
            sine_reg0   <= 36'sb111110010011000101001111010011010;
        end
        7552: begin
            cosine_reg0 <= 36'sb100000111101011000000100000100011100;
            sine_reg0   <= 36'sb111110001100111111001011110110010;
        end
        7553: begin
            cosine_reg0 <= 36'sb100000111101001011110111000000001011;
            sine_reg0   <= 36'sb111110000110111001000101111111110;
        end
        7554: begin
            cosine_reg0 <= 36'sb100000111100111111101011001000100001;
            sine_reg0   <= 36'sb111110000000110010111101101111111;
        end
        7555: begin
            cosine_reg0 <= 36'sb100000111100110011100000011101011101;
            sine_reg0   <= 36'sb111101111010101100110011000111001;
        end
        7556: begin
            cosine_reg0 <= 36'sb100000111100100111010110111111000000;
            sine_reg0   <= 36'sb111101110100100110100110000101101;
        end
        7557: begin
            cosine_reg0 <= 36'sb100000111100011011001110101101001011;
            sine_reg0   <= 36'sb111101101110100000010110101011100;
        end
        7558: begin
            cosine_reg0 <= 36'sb100000111100001111000111100111111110;
            sine_reg0   <= 36'sb111101101000011010000100111001001;
        end
        7559: begin
            cosine_reg0 <= 36'sb100000111100000011000001101111011010;
            sine_reg0   <= 36'sb111101100010010011110000101110101;
        end
        7560: begin
            cosine_reg0 <= 36'sb100000111011110110111101000011011111;
            sine_reg0   <= 36'sb111101011100001101011010001100011;
        end
        7561: begin
            cosine_reg0 <= 36'sb100000111011101010111001100100001101;
            sine_reg0   <= 36'sb111101010110000111000001010010011;
        end
        7562: begin
            cosine_reg0 <= 36'sb100000111011011110110111010001100101;
            sine_reg0   <= 36'sb111101010000000000100110000001001;
        end
        7563: begin
            cosine_reg0 <= 36'sb100000111011010010110110001011101000;
            sine_reg0   <= 36'sb111101001001111010001000011000110;
        end
        7564: begin
            cosine_reg0 <= 36'sb100000111011000110110110010010010110;
            sine_reg0   <= 36'sb111101000011110011101000011001100;
        end
        7565: begin
            cosine_reg0 <= 36'sb100000111010111010110111100101101111;
            sine_reg0   <= 36'sb111100111101101101000110000011100;
        end
        7566: begin
            cosine_reg0 <= 36'sb100000111010101110111010000101110100;
            sine_reg0   <= 36'sb111100110111100110100001010111001;
        end
        7567: begin
            cosine_reg0 <= 36'sb100000111010100010111101110010100101;
            sine_reg0   <= 36'sb111100110001011111111010010100101;
        end
        7568: begin
            cosine_reg0 <= 36'sb100000111010010111000010101100000011;
            sine_reg0   <= 36'sb111100101011011001010000111100001;
        end
        7569: begin
            cosine_reg0 <= 36'sb100000111010001011001000110010001111;
            sine_reg0   <= 36'sb111100100101010010100101001101111;
        end
        7570: begin
            cosine_reg0 <= 36'sb100000111001111111010000000101001000;
            sine_reg0   <= 36'sb111100011111001011110111001010001;
        end
        7571: begin
            cosine_reg0 <= 36'sb100000111001110011011000100100101111;
            sine_reg0   <= 36'sb111100011001000101000110110001010;
        end
        7572: begin
            cosine_reg0 <= 36'sb100000111001100111100010010001000100;
            sine_reg0   <= 36'sb111100010010111110010100000011010;
        end
        7573: begin
            cosine_reg0 <= 36'sb100000111001011011101101001010001001;
            sine_reg0   <= 36'sb111100001100110111011111000000100;
        end
        7574: begin
            cosine_reg0 <= 36'sb100000111001001111111001001111111110;
            sine_reg0   <= 36'sb111100000110110000100111101001010;
        end
        7575: begin
            cosine_reg0 <= 36'sb100000111001000100000110100010100010;
            sine_reg0   <= 36'sb111100000000101001101101111101101;
        end
        7576: begin
            cosine_reg0 <= 36'sb100000111000111000010101000001110111;
            sine_reg0   <= 36'sb111011111010100010110001111110000;
        end
        7577: begin
            cosine_reg0 <= 36'sb100000111000101100100100101101111101;
            sine_reg0   <= 36'sb111011110100011011110011101010100;
        end
        7578: begin
            cosine_reg0 <= 36'sb100000111000100000110101100110110100;
            sine_reg0   <= 36'sb111011101110010100110011000011011;
        end
        7579: begin
            cosine_reg0 <= 36'sb100000111000010101000111101100011100;
            sine_reg0   <= 36'sb111011101000001101110000001001000;
        end
        7580: begin
            cosine_reg0 <= 36'sb100000111000001001011010111110111000;
            sine_reg0   <= 36'sb111011100010000110101010111011011;
        end
        7581: begin
            cosine_reg0 <= 36'sb100000110111111101101111011110000101;
            sine_reg0   <= 36'sb111011011011111111100011011010111;
        end
        7582: begin
            cosine_reg0 <= 36'sb100000110111110010000101001010000110;
            sine_reg0   <= 36'sb111011010101111000011001100111110;
        end
        7583: begin
            cosine_reg0 <= 36'sb100000110111100110011100000010111011;
            sine_reg0   <= 36'sb111011001111110001001101100010010;
        end
        7584: begin
            cosine_reg0 <= 36'sb100000110111011010110100001000100011;
            sine_reg0   <= 36'sb111011001001101001111111001010100;
        end
        7585: begin
            cosine_reg0 <= 36'sb100000110111001111001101011011000000;
            sine_reg0   <= 36'sb111011000011100010101110100000111;
        end
        7586: begin
            cosine_reg0 <= 36'sb100000110111000011100111111010010011;
            sine_reg0   <= 36'sb111010111101011011011011100101100;
        end
        7587: begin
            cosine_reg0 <= 36'sb100000110110111000000011100110011010;
            sine_reg0   <= 36'sb111010110111010100000110011000101;
        end
        7588: begin
            cosine_reg0 <= 36'sb100000110110101100100000011111010111;
            sine_reg0   <= 36'sb111010110001001100101110111010100;
        end
        7589: begin
            cosine_reg0 <= 36'sb100000110110100000111110100101001011;
            sine_reg0   <= 36'sb111010101011000101010101001011011;
        end
        7590: begin
            cosine_reg0 <= 36'sb100000110110010101011101110111110101;
            sine_reg0   <= 36'sb111010100100111101111001001011100;
        end
        7591: begin
            cosine_reg0 <= 36'sb100000110110001001111110010111010110;
            sine_reg0   <= 36'sb111010011110110110011010111011000;
        end
        7592: begin
            cosine_reg0 <= 36'sb100000110101111110100000000011101111;
            sine_reg0   <= 36'sb111010011000101110111010011010011;
        end
        7593: begin
            cosine_reg0 <= 36'sb100000110101110011000010111101000001;
            sine_reg0   <= 36'sb111010010010100111010111101001100;
        end
        7594: begin
            cosine_reg0 <= 36'sb100000110101100111100111000011001010;
            sine_reg0   <= 36'sb111010001100011111110010101000111;
        end
        7595: begin
            cosine_reg0 <= 36'sb100000110101011100001100010110001101;
            sine_reg0   <= 36'sb111010000110011000001011011000110;
        end
        7596: begin
            cosine_reg0 <= 36'sb100000110101010000110010110110001001;
            sine_reg0   <= 36'sb111010000000010000100001111001001;
        end
        7597: begin
            cosine_reg0 <= 36'sb100000110101000101011010100010111110;
            sine_reg0   <= 36'sb111001111010001000110110001010100;
        end
        7598: begin
            cosine_reg0 <= 36'sb100000110100111010000011011100101110;
            sine_reg0   <= 36'sb111001110100000001001000001101000;
        end
        7599: begin
            cosine_reg0 <= 36'sb100000110100101110101101100011011001;
            sine_reg0   <= 36'sb111001101101111001011000000000110;
        end
        7600: begin
            cosine_reg0 <= 36'sb100000110100100011011000110110111111;
            sine_reg0   <= 36'sb111001100111110001100101100110001;
        end
        7601: begin
            cosine_reg0 <= 36'sb100000110100011000000101010111100000;
            sine_reg0   <= 36'sb111001100001101001110000111101011;
        end
        7602: begin
            cosine_reg0 <= 36'sb100000110100001100110011000100111110;
            sine_reg0   <= 36'sb111001011011100001111010000110101;
        end
        7603: begin
            cosine_reg0 <= 36'sb100000110100000001100001111111010111;
            sine_reg0   <= 36'sb111001010101011010000001000010001;
        end
        7604: begin
            cosine_reg0 <= 36'sb100000110011110110010010000110101110;
            sine_reg0   <= 36'sb111001001111010010000101110000010;
        end
        7605: begin
            cosine_reg0 <= 36'sb100000110011101011000011011011000010;
            sine_reg0   <= 36'sb111001001001001010001000010001001;
        end
        7606: begin
            cosine_reg0 <= 36'sb100000110011011111110101111100010100;
            sine_reg0   <= 36'sb111001000011000010001000100101000;
        end
        7607: begin
            cosine_reg0 <= 36'sb100000110011010100101001101010100100;
            sine_reg0   <= 36'sb111000111100111010000110101100001;
        end
        7608: begin
            cosine_reg0 <= 36'sb100000110011001001011110100101110010;
            sine_reg0   <= 36'sb111000110110110010000010100110110;
        end
        7609: begin
            cosine_reg0 <= 36'sb100000110010111110010100101110000000;
            sine_reg0   <= 36'sb111000110000101001111100010101000;
        end
        7610: begin
            cosine_reg0 <= 36'sb100000110010110011001100000011001101;
            sine_reg0   <= 36'sb111000101010100001110011110111010;
        end
        7611: begin
            cosine_reg0 <= 36'sb100000110010101000000100100101011010;
            sine_reg0   <= 36'sb111000100100011001101001001101110;
        end
        7612: begin
            cosine_reg0 <= 36'sb100000110010011100111110010100100111;
            sine_reg0   <= 36'sb111000011110010001011100011000101;
        end
        7613: begin
            cosine_reg0 <= 36'sb100000110010010001111001010000110101;
            sine_reg0   <= 36'sb111000011000001001001101011000001;
        end
        7614: begin
            cosine_reg0 <= 36'sb100000110010000110110101011010000100;
            sine_reg0   <= 36'sb111000010010000000111100001100100;
        end
        7615: begin
            cosine_reg0 <= 36'sb100000110001111011110010110000010101;
            sine_reg0   <= 36'sb111000001011111000101000110110000;
        end
        7616: begin
            cosine_reg0 <= 36'sb100000110001110000110001010011101000;
            sine_reg0   <= 36'sb111000000101110000010011010101000;
        end
        7617: begin
            cosine_reg0 <= 36'sb100000110001100101110001000011111101;
            sine_reg0   <= 36'sb110111111111100111111011101001100;
        end
        7618: begin
            cosine_reg0 <= 36'sb100000110001011010110010000001010101;
            sine_reg0   <= 36'sb110111111001011111100001110011111;
        end
        7619: begin
            cosine_reg0 <= 36'sb100000110001001111110100001011110001;
            sine_reg0   <= 36'sb110111110011010111000101110100010;
        end
        7620: begin
            cosine_reg0 <= 36'sb100000110001000100110111100011010000;
            sine_reg0   <= 36'sb110111101101001110100111101011000;
        end
        7621: begin
            cosine_reg0 <= 36'sb100000110000111001111100000111110011;
            sine_reg0   <= 36'sb110111100111000110000111011000010;
        end
        7622: begin
            cosine_reg0 <= 36'sb100000110000101111000001111001011011;
            sine_reg0   <= 36'sb110111100000111101100100111100011;
        end
        7623: begin
            cosine_reg0 <= 36'sb100000110000100100001000111000001000;
            sine_reg0   <= 36'sb110111011010110101000000010111100;
        end
        7624: begin
            cosine_reg0 <= 36'sb100000110000011001010001000011111010;
            sine_reg0   <= 36'sb110111010100101100011001101001111;
        end
        7625: begin
            cosine_reg0 <= 36'sb100000110000001110011010011100110010;
            sine_reg0   <= 36'sb110111001110100011110000110011110;
        end
        7626: begin
            cosine_reg0 <= 36'sb100000110000000011100101000010110000;
            sine_reg0   <= 36'sb110111001000011011000101110101010;
        end
        7627: begin
            cosine_reg0 <= 36'sb100000101111111000110000110101110101;
            sine_reg0   <= 36'sb110111000010010010011000101110111;
        end
        7628: begin
            cosine_reg0 <= 36'sb100000101111101101111101110110000010;
            sine_reg0   <= 36'sb110110111100001001101001100000101;
        end
        7629: begin
            cosine_reg0 <= 36'sb100000101111100011001100000011010101;
            sine_reg0   <= 36'sb110110110110000000111000001010111;
        end
        7630: begin
            cosine_reg0 <= 36'sb100000101111011000011011011101110001;
            sine_reg0   <= 36'sb110110101111111000000100101101110;
        end
        7631: begin
            cosine_reg0 <= 36'sb100000101111001101101100000101010101;
            sine_reg0   <= 36'sb110110101001101111001111001001100;
        end
        7632: begin
            cosine_reg0 <= 36'sb100000101111000010111101111010000001;
            sine_reg0   <= 36'sb110110100011100110010111011110100;
        end
        7633: begin
            cosine_reg0 <= 36'sb100000101110111000010000111011110111;
            sine_reg0   <= 36'sb110110011101011101011101101100110;
        end
        7634: begin
            cosine_reg0 <= 36'sb100000101110101101100101001010110110;
            sine_reg0   <= 36'sb110110010111010100100001110100110;
        end
        7635: begin
            cosine_reg0 <= 36'sb100000101110100010111010100110111111;
            sine_reg0   <= 36'sb110110010001001011100011110110101;
        end
        7636: begin
            cosine_reg0 <= 36'sb100000101110011000010001010000010011;
            sine_reg0   <= 36'sb110110001011000010100011110010100;
        end
        7637: begin
            cosine_reg0 <= 36'sb100000101110001101101001000110110010;
            sine_reg0   <= 36'sb110110000100111001100001101000110;
        end
        7638: begin
            cosine_reg0 <= 36'sb100000101110000011000010001010011011;
            sine_reg0   <= 36'sb110101111110110000011101011001101;
        end
        7639: begin
            cosine_reg0 <= 36'sb100000101101111000011100011011010000;
            sine_reg0   <= 36'sb110101111000100111010111000101010;
        end
        7640: begin
            cosine_reg0 <= 36'sb100000101101101101110111111001010010;
            sine_reg0   <= 36'sb110101110010011110001110101011111;
        end
        7641: begin
            cosine_reg0 <= 36'sb100000101101100011010100100100100000;
            sine_reg0   <= 36'sb110101101100010101000100001101111;
        end
        7642: begin
            cosine_reg0 <= 36'sb100000101101011000110010011100111010;
            sine_reg0   <= 36'sb110101100110001011110111101011011;
        end
        7643: begin
            cosine_reg0 <= 36'sb100000101101001110010001100010100010;
            sine_reg0   <= 36'sb110101100000000010101001000100100;
        end
        7644: begin
            cosine_reg0 <= 36'sb100000101101000011110001110101011000;
            sine_reg0   <= 36'sb110101011001111001011000011001110;
        end
        7645: begin
            cosine_reg0 <= 36'sb100000101100111001010011010101011011;
            sine_reg0   <= 36'sb110101010011110000000101101011010;
        end
        7646: begin
            cosine_reg0 <= 36'sb100000101100101110110110000010101101;
            sine_reg0   <= 36'sb110101001101100110110000111001001;
        end
        7647: begin
            cosine_reg0 <= 36'sb100000101100100100011001111101001110;
            sine_reg0   <= 36'sb110101000111011101011010000011110;
        end
        7648: begin
            cosine_reg0 <= 36'sb100000101100011001111111000100111110;
            sine_reg0   <= 36'sb110101000001010100000001001011011;
        end
        7649: begin
            cosine_reg0 <= 36'sb100000101100001111100101011001111110;
            sine_reg0   <= 36'sb110100111011001010100110010000001;
        end
        7650: begin
            cosine_reg0 <= 36'sb100000101100000101001100111100001110;
            sine_reg0   <= 36'sb110100110101000001001001010010010;
        end
        7651: begin
            cosine_reg0 <= 36'sb100000101011111010110101101011101110;
            sine_reg0   <= 36'sb110100101110110111101010010010000;
        end
        7652: begin
            cosine_reg0 <= 36'sb100000101011110000011111101000100000;
            sine_reg0   <= 36'sb110100101000101110001001001111110;
        end
        7653: begin
            cosine_reg0 <= 36'sb100000101011100110001010110010100010;
            sine_reg0   <= 36'sb110100100010100100100110001011101;
        end
        7654: begin
            cosine_reg0 <= 36'sb100000101011011011110111001001110110;
            sine_reg0   <= 36'sb110100011100011011000001000101110;
        end
        7655: begin
            cosine_reg0 <= 36'sb100000101011010001100100101110011100;
            sine_reg0   <= 36'sb110100010110010001011001111110100;
        end
        7656: begin
            cosine_reg0 <= 36'sb100000101011000111010011100000010101;
            sine_reg0   <= 36'sb110100010000000111110000110110001;
        end
        7657: begin
            cosine_reg0 <= 36'sb100000101010111101000011011111100001;
            sine_reg0   <= 36'sb110100001001111110000101101100111;
        end
        7658: begin
            cosine_reg0 <= 36'sb100000101010110010110100101100000000;
            sine_reg0   <= 36'sb110100000011110100011000100010111;
        end
        7659: begin
            cosine_reg0 <= 36'sb100000101010101000100111000101110010;
            sine_reg0   <= 36'sb110011111101101010101001011000011;
        end
        7660: begin
            cosine_reg0 <= 36'sb100000101010011110011010101100111001;
            sine_reg0   <= 36'sb110011110111100000111000001101110;
        end
        7661: begin
            cosine_reg0 <= 36'sb100000101010010100001111100001010011;
            sine_reg0   <= 36'sb110011110001010111000101000011001;
        end
        7662: begin
            cosine_reg0 <= 36'sb100000101010001010000101100011000011;
            sine_reg0   <= 36'sb110011101011001101001111111000110;
        end
        7663: begin
            cosine_reg0 <= 36'sb100000101001111111111100110010001000;
            sine_reg0   <= 36'sb110011100101000011011000101110111;
        end
        7664: begin
            cosine_reg0 <= 36'sb100000101001110101110101001110100011;
            sine_reg0   <= 36'sb110011011110111001011111100101110;
        end
        7665: begin
            cosine_reg0 <= 36'sb100000101001101011101110111000010011;
            sine_reg0   <= 36'sb110011011000101111100100011101100;
        end
        7666: begin
            cosine_reg0 <= 36'sb100000101001100001101001101111011010;
            sine_reg0   <= 36'sb110011010010100101100111010110100;
        end
        7667: begin
            cosine_reg0 <= 36'sb100000101001010111100101110011111000;
            sine_reg0   <= 36'sb110011001100011011101000010001000;
        end
        7668: begin
            cosine_reg0 <= 36'sb100000101001001101100011000101101101;
            sine_reg0   <= 36'sb110011000110010001100111001101001;
        end
        7669: begin
            cosine_reg0 <= 36'sb100000101001000011100001100100111010;
            sine_reg0   <= 36'sb110011000000000111100100001011010;
        end
        7670: begin
            cosine_reg0 <= 36'sb100000101000111001100001010001011110;
            sine_reg0   <= 36'sb110010111001111101011111001011100;
        end
        7671: begin
            cosine_reg0 <= 36'sb100000101000101111100010001011011011;
            sine_reg0   <= 36'sb110010110011110011011000001110001;
        end
        7672: begin
            cosine_reg0 <= 36'sb100000101000100101100100010010110000;
            sine_reg0   <= 36'sb110010101101101001001111010011011;
        end
        7673: begin
            cosine_reg0 <= 36'sb100000101000011011100111100111011111;
            sine_reg0   <= 36'sb110010100111011111000100011011100;
        end
        7674: begin
            cosine_reg0 <= 36'sb100000101000010001101100001001100111;
            sine_reg0   <= 36'sb110010100001010100110111100110110;
        end
        7675: begin
            cosine_reg0 <= 36'sb100000101000000111110001111001001001;
            sine_reg0   <= 36'sb110010011011001010101000110101011;
        end
        7676: begin
            cosine_reg0 <= 36'sb100000100111111101111000110110000101;
            sine_reg0   <= 36'sb110010010101000000011000000111100;
        end
        7677: begin
            cosine_reg0 <= 36'sb100000100111110100000001000000011011;
            sine_reg0   <= 36'sb110010001110110110000101011101100;
        end
        7678: begin
            cosine_reg0 <= 36'sb100000100111101010001010011000001101;
            sine_reg0   <= 36'sb110010001000101011110000110111101;
        end
        7679: begin
            cosine_reg0 <= 36'sb100000100111100000010100111101011010;
            sine_reg0   <= 36'sb110010000010100001011010010101111;
        end
        7680: begin
            cosine_reg0 <= 36'sb100000100111010110100000110000000011;
            sine_reg0   <= 36'sb110001111100010111000001111000110;
        end
        7681: begin
            cosine_reg0 <= 36'sb100000100111001100101101110000001000;
            sine_reg0   <= 36'sb110001110110001100100111100000100;
        end
        7682: begin
            cosine_reg0 <= 36'sb100000100111000010111011111101101010;
            sine_reg0   <= 36'sb110001110000000010001011001101001;
        end
        7683: begin
            cosine_reg0 <= 36'sb100000100110111001001011011000101000;
            sine_reg0   <= 36'sb110001101001110111101100111111000;
        end
        7684: begin
            cosine_reg0 <= 36'sb100000100110101111011100000001000100;
            sine_reg0   <= 36'sb110001100011101101001100110110011;
        end
        7685: begin
            cosine_reg0 <= 36'sb100000100110100101101101110110111101;
            sine_reg0   <= 36'sb110001011101100010101010110011100;
        end
        7686: begin
            cosine_reg0 <= 36'sb100000100110011100000000111010010101;
            sine_reg0   <= 36'sb110001010111011000000110110110100;
        end
        7687: begin
            cosine_reg0 <= 36'sb100000100110010010010101001011001010;
            sine_reg0   <= 36'sb110001010001001101100000111111111;
        end
        7688: begin
            cosine_reg0 <= 36'sb100000100110001000101010101001011111;
            sine_reg0   <= 36'sb110001001011000010111001001111100;
        end
        7689: begin
            cosine_reg0 <= 36'sb100000100101111111000001010101010011;
            sine_reg0   <= 36'sb110001000100111000001111100101111;
        end
        7690: begin
            cosine_reg0 <= 36'sb100000100101110101011001001110100110;
            sine_reg0   <= 36'sb110000111110101101100100000011001;
        end
        7691: begin
            cosine_reg0 <= 36'sb100000100101101011110010010101011001;
            sine_reg0   <= 36'sb110000111000100010110110100111101;
        end
        7692: begin
            cosine_reg0 <= 36'sb100000100101100010001100101001101100;
            sine_reg0   <= 36'sb110000110010011000000111010011011;
        end
        7693: begin
            cosine_reg0 <= 36'sb100000100101011000101000001011100000;
            sine_reg0   <= 36'sb110000101100001101010110000110110;
        end
        7694: begin
            cosine_reg0 <= 36'sb100000100101001111000100111010110101;
            sine_reg0   <= 36'sb110000100110000010100011000010001;
        end
        7695: begin
            cosine_reg0 <= 36'sb100000100101000101100010110111101011;
            sine_reg0   <= 36'sb110000011111110111101110000101100;
        end
        7696: begin
            cosine_reg0 <= 36'sb100000100100111100000010000010000100;
            sine_reg0   <= 36'sb110000011001101100110111010001010;
        end
        7697: begin
            cosine_reg0 <= 36'sb100000100100110010100010011001111110;
            sine_reg0   <= 36'sb110000010011100001111110100101100;
        end
        7698: begin
            cosine_reg0 <= 36'sb100000100100101001000011111111011010;
            sine_reg0   <= 36'sb110000001101010111000100000010101;
        end
        7699: begin
            cosine_reg0 <= 36'sb100000100100011111100110110010011010;
            sine_reg0   <= 36'sb110000000111001100000111101000110;
        end
        7700: begin
            cosine_reg0 <= 36'sb100000100100010110001010110010111100;
            sine_reg0   <= 36'sb110000000001000001001001011000010;
        end
        7701: begin
            cosine_reg0 <= 36'sb100000100100001100110000000001000011;
            sine_reg0   <= 36'sb101111111010110110001001010001001;
        end
        7702: begin
            cosine_reg0 <= 36'sb100000100100000011010110011100101101;
            sine_reg0   <= 36'sb101111110100101011000111010011111;
        end
        7703: begin
            cosine_reg0 <= 36'sb100000100011111001111110000101111011;
            sine_reg0   <= 36'sb101111101110100000000011100000101;
        end
        7704: begin
            cosine_reg0 <= 36'sb100000100011110000100110111100101110;
            sine_reg0   <= 36'sb101111101000010100111101110111101;
        end
        7705: begin
            cosine_reg0 <= 36'sb100000100011100111010001000001000110;
            sine_reg0   <= 36'sb101111100010001001110110011001001;
        end
        7706: begin
            cosine_reg0 <= 36'sb100000100011011101111100010011000100;
            sine_reg0   <= 36'sb101111011011111110101101000101010;
        end
        7707: begin
            cosine_reg0 <= 36'sb100000100011010100101000110010100111;
            sine_reg0   <= 36'sb101111010101110011100001111100011;
        end
        7708: begin
            cosine_reg0 <= 36'sb100000100011001011010110011111110000;
            sine_reg0   <= 36'sb101111001111101000010100111110101;
        end
        7709: begin
            cosine_reg0 <= 36'sb100000100011000010000101011010100000;
            sine_reg0   <= 36'sb101111001001011101000110001100011;
        end
        7710: begin
            cosine_reg0 <= 36'sb100000100010111000110101100010110110;
            sine_reg0   <= 36'sb101111000011010001110101100101111;
        end
        7711: begin
            cosine_reg0 <= 36'sb100000100010101111100110111000110100;
            sine_reg0   <= 36'sb101110111101000110100011001011001;
        end
        7712: begin
            cosine_reg0 <= 36'sb100000100010100110011001011100011001;
            sine_reg0   <= 36'sb101110110110111011001110111100101;
        end
        7713: begin
            cosine_reg0 <= 36'sb100000100010011101001101001101100110;
            sine_reg0   <= 36'sb101110110000101111111000111010100;
        end
        7714: begin
            cosine_reg0 <= 36'sb100000100010010100000010001100011011;
            sine_reg0   <= 36'sb101110101010100100100001000100111;
        end
        7715: begin
            cosine_reg0 <= 36'sb100000100010001010111000011000111001;
            sine_reg0   <= 36'sb101110100100011001000111011100010;
        end
        7716: begin
            cosine_reg0 <= 36'sb100000100010000001101111110010111111;
            sine_reg0   <= 36'sb101110011110001101101100000000101;
        end
        7717: begin
            cosine_reg0 <= 36'sb100000100001111000101000011010101111;
            sine_reg0   <= 36'sb101110011000000010001110110010011;
        end
        7718: begin
            cosine_reg0 <= 36'sb100000100001101111100010010000001001;
            sine_reg0   <= 36'sb101110010001110110101111110001110;
        end
        7719: begin
            cosine_reg0 <= 36'sb100000100001100110011101010011001101;
            sine_reg0   <= 36'sb101110001011101011001110111110111;
        end
        7720: begin
            cosine_reg0 <= 36'sb100000100001011101011001100011111010;
            sine_reg0   <= 36'sb101110000101011111101100011010000;
        end
        7721: begin
            cosine_reg0 <= 36'sb100000100001010100010111000010010011;
            sine_reg0   <= 36'sb101101111111010100001000000011100;
        end
        7722: begin
            cosine_reg0 <= 36'sb100000100001001011010101101110010111;
            sine_reg0   <= 36'sb101101111001001000100001111011100;
        end
        7723: begin
            cosine_reg0 <= 36'sb100000100001000010010101101000000110;
            sine_reg0   <= 36'sb101101110010111100111010000010010;
        end
        7724: begin
            cosine_reg0 <= 36'sb100000100000111001010110101111100000;
            sine_reg0   <= 36'sb101101101100110001010000011000000;
        end
        7725: begin
            cosine_reg0 <= 36'sb100000100000110000011001000100100111;
            sine_reg0   <= 36'sb101101100110100101100100111101000;
        end
        7726: begin
            cosine_reg0 <= 36'sb100000100000100111011100100111011010;
            sine_reg0   <= 36'sb101101100000011001110111110001100;
        end
        7727: begin
            cosine_reg0 <= 36'sb100000100000011110100001010111111010;
            sine_reg0   <= 36'sb101101011010001110001000110101110;
        end
        7728: begin
            cosine_reg0 <= 36'sb100000100000010101100111010110000111;
            sine_reg0   <= 36'sb101101010100000010011000001001111;
        end
        7729: begin
            cosine_reg0 <= 36'sb100000100000001100101110100010000010;
            sine_reg0   <= 36'sb101101001101110110100101101110010;
        end
        7730: begin
            cosine_reg0 <= 36'sb100000100000000011110110111011101010;
            sine_reg0   <= 36'sb101101000111101010110001100011000;
        end
        7731: begin
            cosine_reg0 <= 36'sb100000011111111011000000100011000001;
            sine_reg0   <= 36'sb101101000001011110111011101000100;
        end
        7732: begin
            cosine_reg0 <= 36'sb100000011111110010001011011000000110;
            sine_reg0   <= 36'sb101100111011010011000011111110111;
        end
        7733: begin
            cosine_reg0 <= 36'sb100000011111101001010111011010111001;
            sine_reg0   <= 36'sb101100110101000111001010100110011;
        end
        7734: begin
            cosine_reg0 <= 36'sb100000011111100000100100101011011100;
            sine_reg0   <= 36'sb101100101110111011001111011111010;
        end
        7735: begin
            cosine_reg0 <= 36'sb100000011111010111110011001001101111;
            sine_reg0   <= 36'sb101100101000101111010010101001111;
        end
        7736: begin
            cosine_reg0 <= 36'sb100000011111001111000010110101110001;
            sine_reg0   <= 36'sb101100100010100011010100000110010;
        end
        7737: begin
            cosine_reg0 <= 36'sb100000011111000110010011101111100011;
            sine_reg0   <= 36'sb101100011100010111010011110100110;
        end
        7738: begin
            cosine_reg0 <= 36'sb100000011110111101100101110111000110;
            sine_reg0   <= 36'sb101100010110001011010001110101100;
        end
        7739: begin
            cosine_reg0 <= 36'sb100000011110110100111001001100011010;
            sine_reg0   <= 36'sb101100001111111111001110001001000;
        end
        7740: begin
            cosine_reg0 <= 36'sb100000011110101100001101101111011111;
            sine_reg0   <= 36'sb101100001001110011001000101111001;
        end
        7741: begin
            cosine_reg0 <= 36'sb100000011110100011100011100000010101;
            sine_reg0   <= 36'sb101100000011100111000001101000100;
        end
        7742: begin
            cosine_reg0 <= 36'sb100000011110011010111010011110111101;
            sine_reg0   <= 36'sb101011111101011010111000110101000;
        end
        7743: begin
            cosine_reg0 <= 36'sb100000011110010010010010101011011000;
            sine_reg0   <= 36'sb101011110111001110101110010101001;
        end
        7744: begin
            cosine_reg0 <= 36'sb100000011110001001101100000101100101;
            sine_reg0   <= 36'sb101011110001000010100010001001001;
        end
        7745: begin
            cosine_reg0 <= 36'sb100000011110000001000110101101100100;
            sine_reg0   <= 36'sb101011101010110110010100010001000;
        end
        7746: begin
            cosine_reg0 <= 36'sb100000011101111000100010100011010111;
            sine_reg0   <= 36'sb101011100100101010000100101101001;
        end
        7747: begin
            cosine_reg0 <= 36'sb100000011101101111111111100110111110;
            sine_reg0   <= 36'sb101011011110011101110011011101110;
        end
        7748: begin
            cosine_reg0 <= 36'sb100000011101100111011101111000011000;
            sine_reg0   <= 36'sb101011011000010001100000100011001;
        end
        7749: begin
            cosine_reg0 <= 36'sb100000011101011110111101010111100111;
            sine_reg0   <= 36'sb101011010010000101001011111101100;
        end
        7750: begin
            cosine_reg0 <= 36'sb100000011101010110011110000100101010;
            sine_reg0   <= 36'sb101011001011111000110101101101000;
        end
        7751: begin
            cosine_reg0 <= 36'sb100000011101001101111111111111100001;
            sine_reg0   <= 36'sb101011000101101100011101110010000;
        end
        7752: begin
            cosine_reg0 <= 36'sb100000011101000101100011001000001110;
            sine_reg0   <= 36'sb101010111111100000000100001100101;
        end
        7753: begin
            cosine_reg0 <= 36'sb100000011100111101000111011110110001;
            sine_reg0   <= 36'sb101010111001010011101000111101010;
        end
        7754: begin
            cosine_reg0 <= 36'sb100000011100110100101101000011001001;
            sine_reg0   <= 36'sb101010110011000111001100000100000;
        end
        7755: begin
            cosine_reg0 <= 36'sb100000011100101100010011110101010111;
            sine_reg0   <= 36'sb101010101100111010101101100001001;
        end
        7756: begin
            cosine_reg0 <= 36'sb100000011100100011111011110101011100;
            sine_reg0   <= 36'sb101010100110101110001101010100111;
        end
        7757: begin
            cosine_reg0 <= 36'sb100000011100011011100101000011010111;
            sine_reg0   <= 36'sb101010100000100001101011011111100;
        end
        7758: begin
            cosine_reg0 <= 36'sb100000011100010011001111011111001010;
            sine_reg0   <= 36'sb101010011010010101001000000001011;
        end
        7759: begin
            cosine_reg0 <= 36'sb100000011100001010111011001000110100;
            sine_reg0   <= 36'sb101010010100001000100010111010100;
        end
        7760: begin
            cosine_reg0 <= 36'sb100000011100000010101000000000010101;
            sine_reg0   <= 36'sb101010001101111011111100001011001;
        end
        7761: begin
            cosine_reg0 <= 36'sb100000011011111010010110000101101111;
            sine_reg0   <= 36'sb101010000111101111010011110011110;
        end
        7762: begin
            cosine_reg0 <= 36'sb100000011011110010000101011001000001;
            sine_reg0   <= 36'sb101010000001100010101001110100011;
        end
        7763: begin
            cosine_reg0 <= 36'sb100000011011101001110101111010001100;
            sine_reg0   <= 36'sb101001111011010101111110001101010;
        end
        7764: begin
            cosine_reg0 <= 36'sb100000011011100001100111101001010000;
            sine_reg0   <= 36'sb101001110101001001010000111110110;
        end
        7765: begin
            cosine_reg0 <= 36'sb100000011011011001011010100110001101;
            sine_reg0   <= 36'sb101001101110111100100010001001000;
        end
        7766: begin
            cosine_reg0 <= 36'sb100000011011010001001110110001000100;
            sine_reg0   <= 36'sb101001101000101111110001101100010;
        end
        7767: begin
            cosine_reg0 <= 36'sb100000011011001001000100001001110101;
            sine_reg0   <= 36'sb101001100010100010111111101000111;
        end
        7768: begin
            cosine_reg0 <= 36'sb100000011011000000111010110000100000;
            sine_reg0   <= 36'sb101001011100010110001011111110111;
        end
        7769: begin
            cosine_reg0 <= 36'sb100000011010111000110010100101000101;
            sine_reg0   <= 36'sb101001010110001001010110101110110;
        end
        7770: begin
            cosine_reg0 <= 36'sb100000011010110000101011100111100110;
            sine_reg0   <= 36'sb101001001111111100011111111000100;
        end
        7771: begin
            cosine_reg0 <= 36'sb100000011010101000100101111000000001;
            sine_reg0   <= 36'sb101001001001101111100111011100100;
        end
        7772: begin
            cosine_reg0 <= 36'sb100000011010100000100001010110011001;
            sine_reg0   <= 36'sb101001000011100010101101011011000;
        end
        7773: begin
            cosine_reg0 <= 36'sb100000011010011000011110000010101100;
            sine_reg0   <= 36'sb101000111101010101110001110100010;
        end
        7774: begin
            cosine_reg0 <= 36'sb100000011010010000011011111100111011;
            sine_reg0   <= 36'sb101000110111001000110100101000010;
        end
        7775: begin
            cosine_reg0 <= 36'sb100000011010001000011011000101000110;
            sine_reg0   <= 36'sb101000110000111011110101110111101;
        end
        7776: begin
            cosine_reg0 <= 36'sb100000011010000000011011011011001111;
            sine_reg0   <= 36'sb101000101010101110110101100010010;
        end
        7777: begin
            cosine_reg0 <= 36'sb100000011001111000011100111111010100;
            sine_reg0   <= 36'sb101000100100100001110011101000101;
        end
        7778: begin
            cosine_reg0 <= 36'sb100000011001110000011111110001010111;
            sine_reg0   <= 36'sb101000011110010100110000001010111;
        end
        7779: begin
            cosine_reg0 <= 36'sb100000011001101000100011110001011000;
            sine_reg0   <= 36'sb101000011000000111101011001001011;
        end
        7780: begin
            cosine_reg0 <= 36'sb100000011001100000101000111111010110;
            sine_reg0   <= 36'sb101000010001111010100100100100001;
        end
        7781: begin
            cosine_reg0 <= 36'sb100000011001011000101111011011010011;
            sine_reg0   <= 36'sb101000001011101101011100011011100;
        end
        7782: begin
            cosine_reg0 <= 36'sb100000011001010000110111000101001110;
            sine_reg0   <= 36'sb101000000101100000010010101111110;
        end
        7783: begin
            cosine_reg0 <= 36'sb100000011001001000111111111101001001;
            sine_reg0   <= 36'sb100111111111010011000111100001000;
        end
        7784: begin
            cosine_reg0 <= 36'sb100000011001000001001010000011000010;
            sine_reg0   <= 36'sb100111111001000101111010101111110;
        end
        7785: begin
            cosine_reg0 <= 36'sb100000011000111001010101010110111011;
            sine_reg0   <= 36'sb100111110010111000101100011011111;
        end
        7786: begin
            cosine_reg0 <= 36'sb100000011000110001100001111000110100;
            sine_reg0   <= 36'sb100111101100101011011100100110000;
        end
        7787: begin
            cosine_reg0 <= 36'sb100000011000101001101111101000101101;
            sine_reg0   <= 36'sb100111100110011110001011001110000;
        end
        7788: begin
            cosine_reg0 <= 36'sb100000011000100001111110100110100110;
            sine_reg0   <= 36'sb100111100000010000111000010100011;
        end
        7789: begin
            cosine_reg0 <= 36'sb100000011000011010001110110010100000;
            sine_reg0   <= 36'sb100111011010000011100011111001011;
        end
        7790: begin
            cosine_reg0 <= 36'sb100000011000010010100000001100011011;
            sine_reg0   <= 36'sb100111010011110110001101111101000;
        end
        7791: begin
            cosine_reg0 <= 36'sb100000011000001010110010110100011000;
            sine_reg0   <= 36'sb100111001101101000110110011111101;
        end
        7792: begin
            cosine_reg0 <= 36'sb100000011000000011000110101010010110;
            sine_reg0   <= 36'sb100111000111011011011101100001101;
        end
        7793: begin
            cosine_reg0 <= 36'sb100000010111111011011011101110010101;
            sine_reg0   <= 36'sb100111000001001110000011000011000;
        end
        7794: begin
            cosine_reg0 <= 36'sb100000010111110011110010000000010111;
            sine_reg0   <= 36'sb100110111011000000100111000100001;
        end
        7795: begin
            cosine_reg0 <= 36'sb100000010111101100001001100000011100;
            sine_reg0   <= 36'sb100110110100110011001001100101010;
        end
        7796: begin
            cosine_reg0 <= 36'sb100000010111100100100010001110100011;
            sine_reg0   <= 36'sb100110101110100101101010100110100;
        end
        7797: begin
            cosine_reg0 <= 36'sb100000010111011100111100001010101110;
            sine_reg0   <= 36'sb100110101000011000001010001000010;
        end
        7798: begin
            cosine_reg0 <= 36'sb100000010111010101010111010100111100;
            sine_reg0   <= 36'sb100110100010001010101000001010101;
        end
        7799: begin
            cosine_reg0 <= 36'sb100000010111001101110011101101001101;
            sine_reg0   <= 36'sb100110011011111101000100101110000;
        end
        7800: begin
            cosine_reg0 <= 36'sb100000010111000110010001010011100010;
            sine_reg0   <= 36'sb100110010101101111011111110010100;
        end
        7801: begin
            cosine_reg0 <= 36'sb100000010110111110110000000111111100;
            sine_reg0   <= 36'sb100110001111100001111001011000011;
        end
        7802: begin
            cosine_reg0 <= 36'sb100000010110110111010000001010011010;
            sine_reg0   <= 36'sb100110001001010100010001100000000;
        end
        7803: begin
            cosine_reg0 <= 36'sb100000010110101111110001011010111101;
            sine_reg0   <= 36'sb100110000011000110101000001001011;
        end
        7804: begin
            cosine_reg0 <= 36'sb100000010110101000010011111001100101;
            sine_reg0   <= 36'sb100101111100111000111101010101000;
        end
        7805: begin
            cosine_reg0 <= 36'sb100000010110100000110111100110010011;
            sine_reg0   <= 36'sb100101110110101011010001000010111;
        end
        7806: begin
            cosine_reg0 <= 36'sb100000010110011001011100100001000110;
            sine_reg0   <= 36'sb100101110000011101100011010011011;
        end
        7807: begin
            cosine_reg0 <= 36'sb100000010110010010000010101001111111;
            sine_reg0   <= 36'sb100101101010001111110100000110101;
        end
        7808: begin
            cosine_reg0 <= 36'sb100000010110001010101010000000111111;
            sine_reg0   <= 36'sb100101100100000010000011011101001;
        end
        7809: begin
            cosine_reg0 <= 36'sb100000010110000011010010100110000101;
            sine_reg0   <= 36'sb100101011101110100010001010110111;
        end
        7810: begin
            cosine_reg0 <= 36'sb100000010101111011111100011001010010;
            sine_reg0   <= 36'sb100101010111100110011101110100001;
        end
        7811: begin
            cosine_reg0 <= 36'sb100000010101110100100111011010100110;
            sine_reg0   <= 36'sb100101010001011000101000110101010;
        end
        7812: begin
            cosine_reg0 <= 36'sb100000010101101101010011101010000001;
            sine_reg0   <= 36'sb100101001011001010110010011010011;
        end
        7813: begin
            cosine_reg0 <= 36'sb100000010101100110000001000111100100;
            sine_reg0   <= 36'sb100101000100111100111010100011110;
        end
        7814: begin
            cosine_reg0 <= 36'sb100000010101011110101111110011001111;
            sine_reg0   <= 36'sb100100111110101111000001010001101;
        end
        7815: begin
            cosine_reg0 <= 36'sb100000010101010111011111101101000010;
            sine_reg0   <= 36'sb100100111000100001000110100100010;
        end
        7816: begin
            cosine_reg0 <= 36'sb100000010101010000010000110100111110;
            sine_reg0   <= 36'sb100100110010010011001010011100000;
        end
        7817: begin
            cosine_reg0 <= 36'sb100000010101001001000011001011000010;
            sine_reg0   <= 36'sb100100101100000101001100111000111;
        end
        7818: begin
            cosine_reg0 <= 36'sb100000010101000001110110101111010000;
            sine_reg0   <= 36'sb100100100101110111001101111011010;
        end
        7819: begin
            cosine_reg0 <= 36'sb100000010100111010101011100001100111;
            sine_reg0   <= 36'sb100100011111101001001101100011010;
        end
        7820: begin
            cosine_reg0 <= 36'sb100000010100110011100001100010000111;
            sine_reg0   <= 36'sb100100011001011011001011110001011;
        end
        7821: begin
            cosine_reg0 <= 36'sb100000010100101100011000110000110010;
            sine_reg0   <= 36'sb100100010011001101001000100101101;
        end
        7822: begin
            cosine_reg0 <= 36'sb100000010100100101010001001101100110;
            sine_reg0   <= 36'sb100100001100111111000100000000010;
        end
        7823: begin
            cosine_reg0 <= 36'sb100000010100011110001010111000100101;
            sine_reg0   <= 36'sb100100000110110000111110000001101;
        end
        7824: begin
            cosine_reg0 <= 36'sb100000010100010111000101110001101111;
            sine_reg0   <= 36'sb100100000000100010110110101001111;
        end
        7825: begin
            cosine_reg0 <= 36'sb100000010100010000000001111001000100;
            sine_reg0   <= 36'sb100011111010010100101101111001010;
        end
        7826: begin
            cosine_reg0 <= 36'sb100000010100001000111111001110100100;
            sine_reg0   <= 36'sb100011110100000110100011110000000;
        end
        7827: begin
            cosine_reg0 <= 36'sb100000010100000001111101110010010000;
            sine_reg0   <= 36'sb100011101101111000011000001110100;
        end
        7828: begin
            cosine_reg0 <= 36'sb100000010011111010111101100100000111;
            sine_reg0   <= 36'sb100011100111101010001011010100110;
        end
        7829: begin
            cosine_reg0 <= 36'sb100000010011110011111110100100001011;
            sine_reg0   <= 36'sb100011100001011011111101000011001;
        end
        7830: begin
            cosine_reg0 <= 36'sb100000010011101101000000110010011011;
            sine_reg0   <= 36'sb100011011011001101101101011001111;
        end
        7831: begin
            cosine_reg0 <= 36'sb100000010011100110000100001110110111;
            sine_reg0   <= 36'sb100011010100111111011100011001010;
        end
        7832: begin
            cosine_reg0 <= 36'sb100000010011011111001000111001100001;
            sine_reg0   <= 36'sb100011001110110001001010000001100;
        end
        7833: begin
            cosine_reg0 <= 36'sb100000010011011000001110110010010111;
            sine_reg0   <= 36'sb100011001000100010110110010010110;
        end
        7834: begin
            cosine_reg0 <= 36'sb100000010011010001010101111001011011;
            sine_reg0   <= 36'sb100011000010010100100001001101010;
        end
        7835: begin
            cosine_reg0 <= 36'sb100000010011001010011110001110101101;
            sine_reg0   <= 36'sb100010111100000110001010110001011;
        end
        7836: begin
            cosine_reg0 <= 36'sb100000010011000011100111110010001100;
            sine_reg0   <= 36'sb100010110101110111110010111111011;
        end
        7837: begin
            cosine_reg0 <= 36'sb100000010010111100110010100011111010;
            sine_reg0   <= 36'sb100010101111101001011001110111010;
        end
        7838: begin
            cosine_reg0 <= 36'sb100000010010110101111110100011110110;
            sine_reg0   <= 36'sb100010101001011010111111011001100;
        end
        7839: begin
            cosine_reg0 <= 36'sb100000010010101111001011110010000001;
            sine_reg0   <= 36'sb100010100011001100100011100110010;
        end
        7840: begin
            cosine_reg0 <= 36'sb100000010010101000011010001110011100;
            sine_reg0   <= 36'sb100010011100111110000110011101110;
        end
        7841: begin
            cosine_reg0 <= 36'sb100000010010100001101001111001000101;
            sine_reg0   <= 36'sb100010010110101111101000000000001;
        end
        7842: begin
            cosine_reg0 <= 36'sb100000010010011010111010110001111110;
            sine_reg0   <= 36'sb100010010000100001001000001101111;
        end
        7843: begin
            cosine_reg0 <= 36'sb100000010010010100001100111001000110;
            sine_reg0   <= 36'sb100010001010010010100111000111000;
        end
        7844: begin
            cosine_reg0 <= 36'sb100000010010001101100000001110011111;
            sine_reg0   <= 36'sb100010000100000100000100101011111;
        end
        7845: begin
            cosine_reg0 <= 36'sb100000010010000110110100110010001000;
            sine_reg0   <= 36'sb100001111101110101100000111100110;
        end
        7846: begin
            cosine_reg0 <= 36'sb100000010010000000001010100100000010;
            sine_reg0   <= 36'sb100001110111100110111011111001110;
        end
        7847: begin
            cosine_reg0 <= 36'sb100000010001111001100001100100001100;
            sine_reg0   <= 36'sb100001110001011000010101100011010;
        end
        7848: begin
            cosine_reg0 <= 36'sb100000010001110010111001110010100111;
            sine_reg0   <= 36'sb100001101011001001101101111001011;
        end
        7849: begin
            cosine_reg0 <= 36'sb100000010001101100010011001111010100;
            sine_reg0   <= 36'sb100001100100111011000100111100011;
        end
        7850: begin
            cosine_reg0 <= 36'sb100000010001100101101101111010010010;
            sine_reg0   <= 36'sb100001011110101100011010101100101;
        end
        7851: begin
            cosine_reg0 <= 36'sb100000010001011111001001110011100011;
            sine_reg0   <= 36'sb100001011000011101101111001010010;
        end
        7852: begin
            cosine_reg0 <= 36'sb100000010001011000100110111011000101;
            sine_reg0   <= 36'sb100001010010001111000010010101011;
        end
        7853: begin
            cosine_reg0 <= 36'sb100000010001010010000101010000111010;
            sine_reg0   <= 36'sb100001001100000000010100001110100;
        end
        7854: begin
            cosine_reg0 <= 36'sb100000010001001011100100110101000001;
            sine_reg0   <= 36'sb100001000101110001100100110101110;
        end
        7855: begin
            cosine_reg0 <= 36'sb100000010001000101000101100111011011;
            sine_reg0   <= 36'sb100000111111100010110100001011010;
        end
        7856: begin
            cosine_reg0 <= 36'sb100000010000111110100111101000001000;
            sine_reg0   <= 36'sb100000111001010100000010001111100;
        end
        7857: begin
            cosine_reg0 <= 36'sb100000010000111000001010110111001000;
            sine_reg0   <= 36'sb100000110011000101001111000010011;
        end
        7858: begin
            cosine_reg0 <= 36'sb100000010000110001101111010100011101;
            sine_reg0   <= 36'sb100000101100110110011010100100100;
        end
        7859: begin
            cosine_reg0 <= 36'sb100000010000101011010101000000000100;
            sine_reg0   <= 36'sb100000100110100111100100110101111;
        end
        7860: begin
            cosine_reg0 <= 36'sb100000010000100100111011111010000000;
            sine_reg0   <= 36'sb100000100000011000101101110110110;
        end
        7861: begin
            cosine_reg0 <= 36'sb100000010000011110100100000010010001;
            sine_reg0   <= 36'sb100000011010001001110101100111100;
        end
        7862: begin
            cosine_reg0 <= 36'sb100000010000011000001101011000110110;
            sine_reg0   <= 36'sb100000010011111010111100001000010;
        end
        7863: begin
            cosine_reg0 <= 36'sb100000010000010001110111111101110000;
            sine_reg0   <= 36'sb100000001101101100000001011001010;
        end
        7864: begin
            cosine_reg0 <= 36'sb100000010000001011100011110000111110;
            sine_reg0   <= 36'sb100000000111011101000101011010111;
        end
        7865: begin
            cosine_reg0 <= 36'sb100000010000000101010000110010100010;
            sine_reg0   <= 36'sb100000000001001110001000001101001;
        end
        7866: begin
            cosine_reg0 <= 36'sb100000001111111110111111000010011100;
            sine_reg0   <= 36'sb11111111010111111001001110000100;
        end
        7867: begin
            cosine_reg0 <= 36'sb100000001111111000101110100000101100;
            sine_reg0   <= 36'sb11111110100110000001010000101000;
        end
        7868: begin
            cosine_reg0 <= 36'sb100000001111110010011111001101010001;
            sine_reg0   <= 36'sb11111101110100001001001001011000;
        end
        7869: begin
            cosine_reg0 <= 36'sb100000001111101100010001001000001101;
            sine_reg0   <= 36'sb11111101000010010000111000010110;
        end
        7870: begin
            cosine_reg0 <= 36'sb100000001111100110000100010001011111;
            sine_reg0   <= 36'sb11111100010000011000011101100011;
        end
        7871: begin
            cosine_reg0 <= 36'sb100000001111011111111000101001001000;
            sine_reg0   <= 36'sb11111011011110011111111001000011;
        end
        7872: begin
            cosine_reg0 <= 36'sb100000001111011001101110001111001001;
            sine_reg0   <= 36'sb11111010101100100111001010110101;
        end
        7873: begin
            cosine_reg0 <= 36'sb100000001111010011100101000011100000;
            sine_reg0   <= 36'sb11111001111010101110010010111101;
        end
        7874: begin
            cosine_reg0 <= 36'sb100000001111001101011101000110001111;
            sine_reg0   <= 36'sb11111001001000110101010001011101;
        end
        7875: begin
            cosine_reg0 <= 36'sb100000001111000111010110010111010101;
            sine_reg0   <= 36'sb11111000010110111100000110010101;
        end
        7876: begin
            cosine_reg0 <= 36'sb100000001111000001010000110110110100;
            sine_reg0   <= 36'sb11110111100101000010110001101001;
        end
        7877: begin
            cosine_reg0 <= 36'sb100000001110111011001100100100101010;
            sine_reg0   <= 36'sb11110110110011001001010011011010;
        end
        7878: begin
            cosine_reg0 <= 36'sb100000001110110101001001100000111001;
            sine_reg0   <= 36'sb11110110000001001111101011101010;
        end
        7879: begin
            cosine_reg0 <= 36'sb100000001110101111000111101011100001;
            sine_reg0   <= 36'sb11110101001111010101111010011011;
        end
        7880: begin
            cosine_reg0 <= 36'sb100000001110101001000111000100100010;
            sine_reg0   <= 36'sb11110100011101011011111111101111;
        end
        7881: begin
            cosine_reg0 <= 36'sb100000001110100011000111101011111011;
            sine_reg0   <= 36'sb11110011101011100001111011101000;
        end
        7882: begin
            cosine_reg0 <= 36'sb100000001110011101001001100001101110;
            sine_reg0   <= 36'sb11110010111001100111101110000111;
        end
        7883: begin
            cosine_reg0 <= 36'sb100000001110010111001100100101111011;
            sine_reg0   <= 36'sb11110010000111101101010111001111;
        end
        7884: begin
            cosine_reg0 <= 36'sb100000001110010001010000111000100001;
            sine_reg0   <= 36'sb11110001010101110010110111000010;
        end
        7885: begin
            cosine_reg0 <= 36'sb100000001110001011010110011001100010;
            sine_reg0   <= 36'sb11110000100011111000001101100001;
        end
        7886: begin
            cosine_reg0 <= 36'sb100000001110000101011101001000111100;
            sine_reg0   <= 36'sb11101111110001111101011010101111;
        end
        7887: begin
            cosine_reg0 <= 36'sb100000001101111111100101000110110001;
            sine_reg0   <= 36'sb11101111000000000010011110101101;
        end
        7888: begin
            cosine_reg0 <= 36'sb100000001101111001101110010011000001;
            sine_reg0   <= 36'sb11101110001110000111011001011101;
        end
        7889: begin
            cosine_reg0 <= 36'sb100000001101110011111000101101101100;
            sine_reg0   <= 36'sb11101101011100001100001011000010;
        end
        7890: begin
            cosine_reg0 <= 36'sb100000001101101110000100010110110010;
            sine_reg0   <= 36'sb11101100101010010000110011011101;
        end
        7891: begin
            cosine_reg0 <= 36'sb100000001101101000010001001110010011;
            sine_reg0   <= 36'sb11101011111000010101010010101111;
        end
        7892: begin
            cosine_reg0 <= 36'sb100000001101100010011111010100010000;
            sine_reg0   <= 36'sb11101011000110011001101000111100;
        end
        7893: begin
            cosine_reg0 <= 36'sb100000001101011100101110101000101001;
            sine_reg0   <= 36'sb11101010010100011101110110000101;
        end
        7894: begin
            cosine_reg0 <= 36'sb100000001101010110111111001011011110;
            sine_reg0   <= 36'sb11101001100010100001111010001011;
        end
        7895: begin
            cosine_reg0 <= 36'sb100000001101010001010000111100101111;
            sine_reg0   <= 36'sb11101000110000100101110101010001;
        end
        7896: begin
            cosine_reg0 <= 36'sb100000001101001011100011111100011101;
            sine_reg0   <= 36'sb11100111111110101001100111011001;
        end
        7897: begin
            cosine_reg0 <= 36'sb100000001101000101111000001010100111;
            sine_reg0   <= 36'sb11100111001100101101010000100101;
        end
        7898: begin
            cosine_reg0 <= 36'sb100000001101000000001101100111001110;
            sine_reg0   <= 36'sb11100110011010110000110000110110;
        end
        7899: begin
            cosine_reg0 <= 36'sb100000001100111010100100010010010011;
            sine_reg0   <= 36'sb11100101101000110100001000001111;
        end
        7900: begin
            cosine_reg0 <= 36'sb100000001100110100111100001011110100;
            sine_reg0   <= 36'sb11100100110110110111010110110001;
        end
        7901: begin
            cosine_reg0 <= 36'sb100000001100101111010101010011110100;
            sine_reg0   <= 36'sb11100100000100111010011100011110;
        end
        7902: begin
            cosine_reg0 <= 36'sb100000001100101001101111101010010001;
            sine_reg0   <= 36'sb11100011010010111101011001011000;
        end
        7903: begin
            cosine_reg0 <= 36'sb100000001100100100001011001111001100;
            sine_reg0   <= 36'sb11100010100001000000001101100010;
        end
        7904: begin
            cosine_reg0 <= 36'sb100000001100011110101000000010100110;
            sine_reg0   <= 36'sb11100001101111000010111000111101;
        end
        7905: begin
            cosine_reg0 <= 36'sb100000001100011001000110000100011101;
            sine_reg0   <= 36'sb11100000111101000101011011101011;
        end
        7906: begin
            cosine_reg0 <= 36'sb100000001100010011100101010100110100;
            sine_reg0   <= 36'sb11100000001011000111110101101101;
        end
        7907: begin
            cosine_reg0 <= 36'sb100000001100001110000101110011101001;
            sine_reg0   <= 36'sb11011111011001001010000111000111;
        end
        7908: begin
            cosine_reg0 <= 36'sb100000001100001000100111100000111110;
            sine_reg0   <= 36'sb11011110100111001100001111111001;
        end
        7909: begin
            cosine_reg0 <= 36'sb100000001100000011001010011100110010;
            sine_reg0   <= 36'sb11011101110101001110010000000111;
        end
        7910: begin
            cosine_reg0 <= 36'sb100000001011111101101110100111000101;
            sine_reg0   <= 36'sb11011101000011010000000111110000;
        end
        7911: begin
            cosine_reg0 <= 36'sb100000001011111000010011111111111000;
            sine_reg0   <= 36'sb11011100010001010001110110111001;
        end
        7912: begin
            cosine_reg0 <= 36'sb100000001011110010111010100111001011;
            sine_reg0   <= 36'sb11011011011111010011011101100010;
        end
        7913: begin
            cosine_reg0 <= 36'sb100000001011101101100010011100111110;
            sine_reg0   <= 36'sb11011010101101010100111011101101;
        end
        7914: begin
            cosine_reg0 <= 36'sb100000001011101000001011100001010001;
            sine_reg0   <= 36'sb11011001111011010110010001011101;
        end
        7915: begin
            cosine_reg0 <= 36'sb100000001011100010110101110100000101;
            sine_reg0   <= 36'sb11011001001001010111011110110011;
        end
        7916: begin
            cosine_reg0 <= 36'sb100000001011011101100001010101011010;
            sine_reg0   <= 36'sb11011000010111011000100011110001;
        end
        7917: begin
            cosine_reg0 <= 36'sb100000001011011000001110000101010000;
            sine_reg0   <= 36'sb11010111100101011001100000011001;
        end
        7918: begin
            cosine_reg0 <= 36'sb100000001011010010111100000011100111;
            sine_reg0   <= 36'sb11010110110011011010010100101110;
        end
        7919: begin
            cosine_reg0 <= 36'sb100000001011001101101011010000011111;
            sine_reg0   <= 36'sb11010110000001011011000000110000;
        end
        7920: begin
            cosine_reg0 <= 36'sb100000001011001000011011101011111000;
            sine_reg0   <= 36'sb11010101001111011011100100100010;
        end
        7921: begin
            cosine_reg0 <= 36'sb100000001011000011001101010101110100;
            sine_reg0   <= 36'sb11010100011101011100000000000110;
        end
        7922: begin
            cosine_reg0 <= 36'sb100000001010111110000000001110010010;
            sine_reg0   <= 36'sb11010011101011011100010011011110;
        end
        7923: begin
            cosine_reg0 <= 36'sb100000001010111000110100010101010001;
            sine_reg0   <= 36'sb11010010111001011100011110101100;
        end
        7924: begin
            cosine_reg0 <= 36'sb100000001010110011101001101010110011;
            sine_reg0   <= 36'sb11010010000111011100100001110001;
        end
        7925: begin
            cosine_reg0 <= 36'sb100000001010101110100000001110111000;
            sine_reg0   <= 36'sb11010001010101011100011100110000;
        end
        7926: begin
            cosine_reg0 <= 36'sb100000001010101001011000000001011111;
            sine_reg0   <= 36'sb11010000100011011100001111101010;
        end
        7927: begin
            cosine_reg0 <= 36'sb100000001010100100010001000010101010;
            sine_reg0   <= 36'sb11001111110001011011111010100010;
        end
        7928: begin
            cosine_reg0 <= 36'sb100000001010011111001011010010010111;
            sine_reg0   <= 36'sb11001110111111011011011101011001;
        end
        7929: begin
            cosine_reg0 <= 36'sb100000001010011010000110110000101000;
            sine_reg0   <= 36'sb11001110001101011010111000010001;
        end
        7930: begin
            cosine_reg0 <= 36'sb100000001010010101000011011101011100;
            sine_reg0   <= 36'sb11001101011011011010001011001101;
        end
        7931: begin
            cosine_reg0 <= 36'sb100000001010010000000001011000110101;
            sine_reg0   <= 36'sb11001100101001011001010110001110;
        end
        7932: begin
            cosine_reg0 <= 36'sb100000001010001011000000100010110001;
            sine_reg0   <= 36'sb11001011110111011000011001010101;
        end
        7933: begin
            cosine_reg0 <= 36'sb100000001010000110000000111011010001;
            sine_reg0   <= 36'sb11001011000101010111010100100110;
        end
        7934: begin
            cosine_reg0 <= 36'sb100000001010000001000010100010010110;
            sine_reg0   <= 36'sb11001010010011010110001000000010;
        end
        7935: begin
            cosine_reg0 <= 36'sb100000001001111100000101010111111111;
            sine_reg0   <= 36'sb11001001100001010100110011101010;
        end
        7936: begin
            cosine_reg0 <= 36'sb100000001001110111001001011100001101;
            sine_reg0   <= 36'sb11001000101111010011010111100001;
        end
        7937: begin
            cosine_reg0 <= 36'sb100000001001110010001110101110111111;
            sine_reg0   <= 36'sb11000111111101010001110011101001;
        end
        7938: begin
            cosine_reg0 <= 36'sb100000001001101101010101010000010111;
            sine_reg0   <= 36'sb11000111001011010000001000000100;
        end
        7939: begin
            cosine_reg0 <= 36'sb100000001001101000011101000000010100;
            sine_reg0   <= 36'sb11000110011001001110010100110011;
        end
        7940: begin
            cosine_reg0 <= 36'sb100000001001100011100101111110110111;
            sine_reg0   <= 36'sb11000101100111001100011001111000;
        end
        7941: begin
            cosine_reg0 <= 36'sb100000001001011110110000001011111111;
            sine_reg0   <= 36'sb11000100110101001010010111010110;
        end
        7942: begin
            cosine_reg0 <= 36'sb100000001001011001111011100111101101;
            sine_reg0   <= 36'sb11000100000011001000001101001111;
        end
        7943: begin
            cosine_reg0 <= 36'sb100000001001010101001000010010000010;
            sine_reg0   <= 36'sb11000011010001000101111011100011;
        end
        7944: begin
            cosine_reg0 <= 36'sb100000001001010000010110001010111100;
            sine_reg0   <= 36'sb11000010011111000011100010010110;
        end
        7945: begin
            cosine_reg0 <= 36'sb100000001001001011100101010010011101;
            sine_reg0   <= 36'sb11000001101101000001000001101001;
        end
        7946: begin
            cosine_reg0 <= 36'sb100000001001000110110101101000100100;
            sine_reg0   <= 36'sb11000000111010111110011001011110;
        end
        7947: begin
            cosine_reg0 <= 36'sb100000001001000010000111001101010010;
            sine_reg0   <= 36'sb11000000001000111011101001110111;
        end
        7948: begin
            cosine_reg0 <= 36'sb100000001000111101011010000000100111;
            sine_reg0   <= 36'sb10111111010110111000110010110110;
        end
        7949: begin
            cosine_reg0 <= 36'sb100000001000111000101110000010100011;
            sine_reg0   <= 36'sb10111110100100110101110100011100;
        end
        7950: begin
            cosine_reg0 <= 36'sb100000001000110100000011010011000111;
            sine_reg0   <= 36'sb10111101110010110010101110101101;
        end
        7951: begin
            cosine_reg0 <= 36'sb100000001000101111011001110010010010;
            sine_reg0   <= 36'sb10111101000000101111100001101001;
        end
        7952: begin
            cosine_reg0 <= 36'sb100000001000101010110001100000000101;
            sine_reg0   <= 36'sb10111100001110101100001101010011;
        end
        7953: begin
            cosine_reg0 <= 36'sb100000001000100110001010011100011111;
            sine_reg0   <= 36'sb10111011011100101000110001101100;
        end
        7954: begin
            cosine_reg0 <= 36'sb100000001000100001100100100111100010;
            sine_reg0   <= 36'sb10111010101010100101001110110111;
        end
        7955: begin
            cosine_reg0 <= 36'sb100000001000011101000000000001001100;
            sine_reg0   <= 36'sb10111001111000100001100100110101;
        end
        7956: begin
            cosine_reg0 <= 36'sb100000001000011000011100101001011111;
            sine_reg0   <= 36'sb10111001000110011101110011101001;
        end
        7957: begin
            cosine_reg0 <= 36'sb100000001000010011111010100000011011;
            sine_reg0   <= 36'sb10111000010100011001111011010100;
        end
        7958: begin
            cosine_reg0 <= 36'sb100000001000001111011001100101111111;
            sine_reg0   <= 36'sb10110111100010010101111011111000;
        end
        7959: begin
            cosine_reg0 <= 36'sb100000001000001010111001111010001101;
            sine_reg0   <= 36'sb10110110110000010001110101010111;
        end
        7960: begin
            cosine_reg0 <= 36'sb100000001000000110011011011101000011;
            sine_reg0   <= 36'sb10110101111110001101100111110100;
        end
        7961: begin
            cosine_reg0 <= 36'sb100000001000000001111110001110100011;
            sine_reg0   <= 36'sb10110101001100001001010011001111;
        end
        7962: begin
            cosine_reg0 <= 36'sb100000000111111101100010001110101100;
            sine_reg0   <= 36'sb10110100011010000100110111101011;
        end
        7963: begin
            cosine_reg0 <= 36'sb100000000111111001000111011101011111;
            sine_reg0   <= 36'sb10110011101000000000010101001011;
        end
        7964: begin
            cosine_reg0 <= 36'sb100000000111110100101101111010111011;
            sine_reg0   <= 36'sb10110010110101111011101011101110;
        end
        7965: begin
            cosine_reg0 <= 36'sb100000000111110000010101100111000001;
            sine_reg0   <= 36'sb10110010000011110110111011011001;
        end
        7966: begin
            cosine_reg0 <= 36'sb100000000111101011111110100001110010;
            sine_reg0   <= 36'sb10110001010001110010000100001100;
        end
        7967: begin
            cosine_reg0 <= 36'sb100000000111100111101000101011001100;
            sine_reg0   <= 36'sb10110000011111101101000110001010;
        end
        7968: begin
            cosine_reg0 <= 36'sb100000000111100011010100000011010010;
            sine_reg0   <= 36'sb10101111101101101000000001010101;
        end
        7969: begin
            cosine_reg0 <= 36'sb100000000111011111000000101010000001;
            sine_reg0   <= 36'sb10101110111011100010110101101110;
        end
        7970: begin
            cosine_reg0 <= 36'sb100000000111011010101110011111011100;
            sine_reg0   <= 36'sb10101110001001011101100011010111;
        end
        7971: begin
            cosine_reg0 <= 36'sb100000000111010110011101100011100001;
            sine_reg0   <= 36'sb10101101010111011000001010010010;
        end
        7972: begin
            cosine_reg0 <= 36'sb100000000111010010001101110110010010;
            sine_reg0   <= 36'sb10101100100101010010101010100010;
        end
        7973: begin
            cosine_reg0 <= 36'sb100000000111001101111111010111101110;
            sine_reg0   <= 36'sb10101011110011001101000100001000;
        end
        7974: begin
            cosine_reg0 <= 36'sb100000000111001001110010000111110101;
            sine_reg0   <= 36'sb10101011000001000111010111000110;
        end
        7975: begin
            cosine_reg0 <= 36'sb100000000111000101100110000110101000;
            sine_reg0   <= 36'sb10101010001111000001100011011110;
        end
        7976: begin
            cosine_reg0 <= 36'sb100000000111000001011011010100000111;
            sine_reg0   <= 36'sb10101001011100111011101001010010;
        end
        7977: begin
            cosine_reg0 <= 36'sb100000000110111101010001110000010001;
            sine_reg0   <= 36'sb10101000101010110101101000100100;
        end
        7978: begin
            cosine_reg0 <= 36'sb100000000110111001001001011011001000;
            sine_reg0   <= 36'sb10100111111000101111100001010110;
        end
        7979: begin
            cosine_reg0 <= 36'sb100000000110110101000010010100101010;
            sine_reg0   <= 36'sb10100111000110101001010011101010;
        end
        7980: begin
            cosine_reg0 <= 36'sb100000000110110000111100011100111010;
            sine_reg0   <= 36'sb10100110010100100010111111100001;
        end
        7981: begin
            cosine_reg0 <= 36'sb100000000110101100110111110011110101;
            sine_reg0   <= 36'sb10100101100010011100100100111110;
        end
        7982: begin
            cosine_reg0 <= 36'sb100000000110101000110100011001011110;
            sine_reg0   <= 36'sb10100100110000010110000100000010;
        end
        7983: begin
            cosine_reg0 <= 36'sb100000000110100100110010001101110011;
            sine_reg0   <= 36'sb10100011111110001111011100110000;
        end
        7984: begin
            cosine_reg0 <= 36'sb100000000110100000110001010000110101;
            sine_reg0   <= 36'sb10100011001100001000101111001001;
        end
        7985: begin
            cosine_reg0 <= 36'sb100000000110011100110001100010100101;
            sine_reg0   <= 36'sb10100010011010000001111011010000;
        end
        7986: begin
            cosine_reg0 <= 36'sb100000000110011000110011000011000010;
            sine_reg0   <= 36'sb10100001100111111011000001000110;
        end
        7987: begin
            cosine_reg0 <= 36'sb100000000110010100110101110010001100;
            sine_reg0   <= 36'sb10100000110101110100000000101101;
        end
        7988: begin
            cosine_reg0 <= 36'sb100000000110010000111001110000000100;
            sine_reg0   <= 36'sb10100000000011101100111010000111;
        end
        7989: begin
            cosine_reg0 <= 36'sb100000000110001100111110111100101010;
            sine_reg0   <= 36'sb10011111010001100101101101010110;
        end
        7990: begin
            cosine_reg0 <= 36'sb100000000110001001000101010111111101;
            sine_reg0   <= 36'sb10011110011111011110011010011101;
        end
        7991: begin
            cosine_reg0 <= 36'sb100000000110000101001101000001111111;
            sine_reg0   <= 36'sb10011101101101010111000001011100;
        end
        7992: begin
            cosine_reg0 <= 36'sb100000000110000001010101111010101111;
            sine_reg0   <= 36'sb10011100111011001111100010010110;
        end
        7993: begin
            cosine_reg0 <= 36'sb100000000101111101100000000010001101;
            sine_reg0   <= 36'sb10011100001001000111111101001101;
        end
        7994: begin
            cosine_reg0 <= 36'sb100000000101111001101011011000011010;
            sine_reg0   <= 36'sb10011011010111000000010010000011;
        end
        7995: begin
            cosine_reg0 <= 36'sb100000000101110101110111111101010110;
            sine_reg0   <= 36'sb10011010100100111000100000111001;
        end
        7996: begin
            cosine_reg0 <= 36'sb100000000101110010000101110001000000;
            sine_reg0   <= 36'sb10011001110010110000101001110010;
        end
        7997: begin
            cosine_reg0 <= 36'sb100000000101101110010100110011011001;
            sine_reg0   <= 36'sb10011001000000101000101100101111;
        end
        7998: begin
            cosine_reg0 <= 36'sb100000000101101010100101000100100010;
            sine_reg0   <= 36'sb10011000001110100000101001110011;
        end
        7999: begin
            cosine_reg0 <= 36'sb100000000101100110110110100100011010;
            sine_reg0   <= 36'sb10010111011100011000100001000000;
        end
        8000: begin
            cosine_reg0 <= 36'sb100000000101100011001001010011000001;
            sine_reg0   <= 36'sb10010110101010010000010010010110;
        end
        8001: begin
            cosine_reg0 <= 36'sb100000000101011111011101010000010111;
            sine_reg0   <= 36'sb10010101111000000111111101111001;
        end
        8002: begin
            cosine_reg0 <= 36'sb100000000101011011110010011100011110;
            sine_reg0   <= 36'sb10010101000101111111100011101010;
        end
        8003: begin
            cosine_reg0 <= 36'sb100000000101011000001000110111010100;
            sine_reg0   <= 36'sb10010100010011110111000011101100;
        end
        8004: begin
            cosine_reg0 <= 36'sb100000000101010100100000100000111010;
            sine_reg0   <= 36'sb10010011100001101110011101111111;
        end
        8005: begin
            cosine_reg0 <= 36'sb100000000101010000111001011001010000;
            sine_reg0   <= 36'sb10010010101111100101110010100110;
        end
        8006: begin
            cosine_reg0 <= 36'sb100000000101001101010011100000010111;
            sine_reg0   <= 36'sb10010001111101011101000001100011;
        end
        8007: begin
            cosine_reg0 <= 36'sb100000000101001001101110110110001110;
            sine_reg0   <= 36'sb10010001001011010100001010111000;
        end
        8008: begin
            cosine_reg0 <= 36'sb100000000101000110001011011010110101;
            sine_reg0   <= 36'sb10010000011001001011001110100111;
        end
        8009: begin
            cosine_reg0 <= 36'sb100000000101000010101001001110001101;
            sine_reg0   <= 36'sb10001111100111000010001100110010;
        end
        8010: begin
            cosine_reg0 <= 36'sb100000000100111111001000010000010110;
            sine_reg0   <= 36'sb10001110110100111001000101011010;
        end
        8011: begin
            cosine_reg0 <= 36'sb100000000100111011101000100001010000;
            sine_reg0   <= 36'sb10001110000010101111111000100010;
        end
        8012: begin
            cosine_reg0 <= 36'sb100000000100111000001010000000111011;
            sine_reg0   <= 36'sb10001101010000100110100110001011;
        end
        8013: begin
            cosine_reg0 <= 36'sb100000000100110100101100101111010111;
            sine_reg0   <= 36'sb10001100011110011101001110011000;
        end
        8014: begin
            cosine_reg0 <= 36'sb100000000100110001010000101100100100;
            sine_reg0   <= 36'sb10001011101100010011110001001010;
        end
        8015: begin
            cosine_reg0 <= 36'sb100000000100101101110101111000100011;
            sine_reg0   <= 36'sb10001010111010001010001110100100;
        end
        8016: begin
            cosine_reg0 <= 36'sb100000000100101010011100010011010011;
            sine_reg0   <= 36'sb10001010001000000000100110100111;
        end
        8017: begin
            cosine_reg0 <= 36'sb100000000100100111000011111100110110;
            sine_reg0   <= 36'sb10001001010101110110111001010101;
        end
        8018: begin
            cosine_reg0 <= 36'sb100000000100100011101100110101001010;
            sine_reg0   <= 36'sb10001000100011101101000110110000;
        end
        8019: begin
            cosine_reg0 <= 36'sb100000000100100000010110111100010000;
            sine_reg0   <= 36'sb10000111110001100011001110111010;
        end
        8020: begin
            cosine_reg0 <= 36'sb100000000100011101000010010010001000;
            sine_reg0   <= 36'sb10000110111111011001010001110101;
        end
        8021: begin
            cosine_reg0 <= 36'sb100000000100011001101110110110110010;
            sine_reg0   <= 36'sb10000110001101001111001111100011;
        end
        8022: begin
            cosine_reg0 <= 36'sb100000000100010110011100101010001111;
            sine_reg0   <= 36'sb10000101011011000101001000000110;
        end
        8023: begin
            cosine_reg0 <= 36'sb100000000100010011001011101100011110;
            sine_reg0   <= 36'sb10000100101000111010111011100000;
        end
        8024: begin
            cosine_reg0 <= 36'sb100000000100001111111011111101100000;
            sine_reg0   <= 36'sb10000011110110110000101001110010;
        end
        8025: begin
            cosine_reg0 <= 36'sb100000000100001100101101011101010101;
            sine_reg0   <= 36'sb10000011000100100110010010111111;
        end
        8026: begin
            cosine_reg0 <= 36'sb100000000100001001100000001011111101;
            sine_reg0   <= 36'sb10000010010010011011110111001001;
        end
        8027: begin
            cosine_reg0 <= 36'sb100000000100000110010100001001010111;
            sine_reg0   <= 36'sb10000001100000010001010110010001;
        end
        8028: begin
            cosine_reg0 <= 36'sb100000000100000011001001010101100101;
            sine_reg0   <= 36'sb10000000101110000110110000011010;
        end
        8029: begin
            cosine_reg0 <= 36'sb100000000011111111111111110000100110;
            sine_reg0   <= 36'sb1111111111011111100000101100101;
        end
        8030: begin
            cosine_reg0 <= 36'sb100000000011111100110111011010011010;
            sine_reg0   <= 36'sb1111111001001110001010101110100;
        end
        8031: begin
            cosine_reg0 <= 36'sb100000000011111001110000010011000010;
            sine_reg0   <= 36'sb1111110010111100110100001001010;
        end
        8032: begin
            cosine_reg0 <= 36'sb100000000011110110101010011010011101;
            sine_reg0   <= 36'sb1111101100101011011100111101000;
        end
        8033: begin
            cosine_reg0 <= 36'sb100000000011110011100101110000101101;
            sine_reg0   <= 36'sb1111100110011010000101001010000;
        end
        8034: begin
            cosine_reg0 <= 36'sb100000000011110000100010010101110000;
            sine_reg0   <= 36'sb1111100000001000101100110000100;
        end
        8035: begin
            cosine_reg0 <= 36'sb100000000011101101100000001001100110;
            sine_reg0   <= 36'sb1111011001110111010011110000110;
        end
        8036: begin
            cosine_reg0 <= 36'sb100000000011101010011111001100010001;
            sine_reg0   <= 36'sb1111010011100101111010001011000;
        end
        8037: begin
            cosine_reg0 <= 36'sb100000000011100111011111011101110001;
            sine_reg0   <= 36'sb1111001101010100011111111111100;
        end
        8038: begin
            cosine_reg0 <= 36'sb100000000011100100100000111110000100;
            sine_reg0   <= 36'sb1111000111000011000101001110011;
        end
        8039: begin
            cosine_reg0 <= 36'sb100000000011100001100011101101001100;
            sine_reg0   <= 36'sb1111000000110001101001111000001;
        end
        8040: begin
            cosine_reg0 <= 36'sb100000000011011110100111101011001001;
            sine_reg0   <= 36'sb1110111010100000001101111100110;
        end
        8041: begin
            cosine_reg0 <= 36'sb100000000011011011101100110111111010;
            sine_reg0   <= 36'sb1110110100001110110001011100101;
        end
        8042: begin
            cosine_reg0 <= 36'sb100000000011011000110011010011100000;
            sine_reg0   <= 36'sb1110101101111101010100010111111;
        end
        8043: begin
            cosine_reg0 <= 36'sb100000000011010101111010111101111011;
            sine_reg0   <= 36'sb1110100111101011110110101110111;
        end
        8044: begin
            cosine_reg0 <= 36'sb100000000011010011000011110111001010;
            sine_reg0   <= 36'sb1110100001011010011000100001110;
        end
        8045: begin
            cosine_reg0 <= 36'sb100000000011010000001101111111001111;
            sine_reg0   <= 36'sb1110011011001000111001110000110;
        end
        8046: begin
            cosine_reg0 <= 36'sb100000000011001101011001010110001001;
            sine_reg0   <= 36'sb1110010100110111011010011100010;
        end
        8047: begin
            cosine_reg0 <= 36'sb100000000011001010100101111011111001;
            sine_reg0   <= 36'sb1110001110100101111010100100011;
        end
        8048: begin
            cosine_reg0 <= 36'sb100000000011000111110011110000011110;
            sine_reg0   <= 36'sb1110001000010100011010001001011;
        end
        8049: begin
            cosine_reg0 <= 36'sb100000000011000101000010110011111000;
            sine_reg0   <= 36'sb1110000010000010111001001011100;
        end
        8050: begin
            cosine_reg0 <= 36'sb100000000011000010010011000110001000;
            sine_reg0   <= 36'sb1101111011110001010111101011000;
        end
        8051: begin
            cosine_reg0 <= 36'sb100000000010111111100100100111001110;
            sine_reg0   <= 36'sb1101110101011111110101101000010;
        end
        8052: begin
            cosine_reg0 <= 36'sb100000000010111100110111010111001001;
            sine_reg0   <= 36'sb1101101111001110010011000011010;
        end
        8053: begin
            cosine_reg0 <= 36'sb100000000010111010001011010101111011;
            sine_reg0   <= 36'sb1101101000111100101111111100010;
        end
        8054: begin
            cosine_reg0 <= 36'sb100000000010110111100000100011100011;
            sine_reg0   <= 36'sb1101100010101011001100010011110;
        end
        8055: begin
            cosine_reg0 <= 36'sb100000000010110100110111000000000000;
            sine_reg0   <= 36'sb1101011100011001101000001001110;
        end
        8056: begin
            cosine_reg0 <= 36'sb100000000010110010001110101011010101;
            sine_reg0   <= 36'sb1101010110001000000011011110101;
        end
        8057: begin
            cosine_reg0 <= 36'sb100000000010101111100111100101011111;
            sine_reg0   <= 36'sb1101001111110110011110010010101;
        end
        8058: begin
            cosine_reg0 <= 36'sb100000000010101101000001101110100000;
            sine_reg0   <= 36'sb1101001001100100111000100101111;
        end
        8059: begin
            cosine_reg0 <= 36'sb100000000010101010011101000110010111;
            sine_reg0   <= 36'sb1101000011010011010010011000101;
        end
        8060: begin
            cosine_reg0 <= 36'sb100000000010100111111001101101000101;
            sine_reg0   <= 36'sb1100111101000001101011101011010;
        end
        8061: begin
            cosine_reg0 <= 36'sb100000000010100101010111100010101010;
            sine_reg0   <= 36'sb1100110110110000000100011101111;
        end
        8062: begin
            cosine_reg0 <= 36'sb100000000010100010110110100111000110;
            sine_reg0   <= 36'sb1100110000011110011100110000111;
        end
        8063: begin
            cosine_reg0 <= 36'sb100000000010100000010110111010011001;
            sine_reg0   <= 36'sb1100101010001100110100100100010;
        end
        8064: begin
            cosine_reg0 <= 36'sb100000000010011101111000011100100011;
            sine_reg0   <= 36'sb1100100011111011001011111000100;
        end
        8065: begin
            cosine_reg0 <= 36'sb100000000010011011011011001101100100;
            sine_reg0   <= 36'sb1100011101101001100010101101110;
        end
        8066: begin
            cosine_reg0 <= 36'sb100000000010011000111111001101011100;
            sine_reg0   <= 36'sb1100010111010111111001000100010;
        end
        8067: begin
            cosine_reg0 <= 36'sb100000000010010110100100011100001011;
            sine_reg0   <= 36'sb1100010001000110001110111100001;
        end
        8068: begin
            cosine_reg0 <= 36'sb100000000010010100001010111001110010;
            sine_reg0   <= 36'sb1100001010110100100100010101111;
        end
        8069: begin
            cosine_reg0 <= 36'sb100000000010010001110010100110010001;
            sine_reg0   <= 36'sb1100000100100010111001010001100;
        end
        8070: begin
            cosine_reg0 <= 36'sb100000000010001111011011100001100111;
            sine_reg0   <= 36'sb1011111110010001001101101111011;
        end
        8071: begin
            cosine_reg0 <= 36'sb100000000010001101000101101011110101;
            sine_reg0   <= 36'sb1011110111111111100001101111110;
        end
        8072: begin
            cosine_reg0 <= 36'sb100000000010001010110001000100111010;
            sine_reg0   <= 36'sb1011110001101101110101010010110;
        end
        8073: begin
            cosine_reg0 <= 36'sb100000000010001000011101101100111000;
            sine_reg0   <= 36'sb1011101011011100001000011000110;
        end
        8074: begin
            cosine_reg0 <= 36'sb100000000010000110001011100011101101;
            sine_reg0   <= 36'sb1011100101001010011011000001111;
        end
        8075: begin
            cosine_reg0 <= 36'sb100000000010000011111010101001011011;
            sine_reg0   <= 36'sb1011011110111000101101001110100;
        end
        8076: begin
            cosine_reg0 <= 36'sb100000000010000001101010111110000000;
            sine_reg0   <= 36'sb1011011000100110111110111110110;
        end
        8077: begin
            cosine_reg0 <= 36'sb100000000001111111011100100001011110;
            sine_reg0   <= 36'sb1011010010010101010000010010111;
        end
        8078: begin
            cosine_reg0 <= 36'sb100000000001111101001111010011110100;
            sine_reg0   <= 36'sb1011001100000011100001001011010;
        end
        8079: begin
            cosine_reg0 <= 36'sb100000000001111011000011010101000011;
            sine_reg0   <= 36'sb1011000101110001110001100111111;
        end
        8080: begin
            cosine_reg0 <= 36'sb100000000001111000111000100101001010;
            sine_reg0   <= 36'sb1010111111100000000001101001010;
        end
        8081: begin
            cosine_reg0 <= 36'sb100000000001110110101111000100001010;
            sine_reg0   <= 36'sb1010111001001110010001001111100;
        end
        8082: begin
            cosine_reg0 <= 36'sb100000000001110100100110110010000010;
            sine_reg0   <= 36'sb1010110010111100100000011010111;
        end
        8083: begin
            cosine_reg0 <= 36'sb100000000001110010011111101110110011;
            sine_reg0   <= 36'sb1010101100101010101111001011100;
        end
        8084: begin
            cosine_reg0 <= 36'sb100000000001110000011001111010011101;
            sine_reg0   <= 36'sb1010100110011000111101100001111;
        end
        8085: begin
            cosine_reg0 <= 36'sb100000000001101110010101010101000000;
            sine_reg0   <= 36'sb1010100000000111001011011110000;
        end
        8086: begin
            cosine_reg0 <= 36'sb100000000001101100010001111110011100;
            sine_reg0   <= 36'sb1010011001110101011001000000010;
        end
        8087: begin
            cosine_reg0 <= 36'sb100000000001101010001111110110110001;
            sine_reg0   <= 36'sb1010010011100011100110001000111;
        end
        8088: begin
            cosine_reg0 <= 36'sb100000000001101000001110111101111111;
            sine_reg0   <= 36'sb1010001101010001110010111000000;
        end
        8089: begin
            cosine_reg0 <= 36'sb100000000001100110001111010100000110;
            sine_reg0   <= 36'sb1010000110111111111111001110000;
        end
        8090: begin
            cosine_reg0 <= 36'sb100000000001100100010000111001000111;
            sine_reg0   <= 36'sb1010000000101110001011001011000;
        end
        8091: begin
            cosine_reg0 <= 36'sb100000000001100010010011101101000001;
            sine_reg0   <= 36'sb1001111010011100010110101111010;
        end
        8092: begin
            cosine_reg0 <= 36'sb100000000001100000010111101111110100;
            sine_reg0   <= 36'sb1001110100001010100001111011001;
        end
        8093: begin
            cosine_reg0 <= 36'sb100000000001011110011101000001100001;
            sine_reg0   <= 36'sb1001101101111000101100101110110;
        end
        8094: begin
            cosine_reg0 <= 36'sb100000000001011100100011100010000111;
            sine_reg0   <= 36'sb1001100111100110110111001010011;
        end
        8095: begin
            cosine_reg0 <= 36'sb100000000001011010101011010001100111;
            sine_reg0   <= 36'sb1001100001010101000001001110011;
        end
        8096: begin
            cosine_reg0 <= 36'sb100000000001011000110100010000000001;
            sine_reg0   <= 36'sb1001011011000011001010111010110;
        end
        8097: begin
            cosine_reg0 <= 36'sb100000000001010110111110011101010101;
            sine_reg0   <= 36'sb1001010100110001010100010000000;
        end
        8098: begin
            cosine_reg0 <= 36'sb100000000001010101001001111001100011;
            sine_reg0   <= 36'sb1001001110011111011101001110001;
        end
        8099: begin
            cosine_reg0 <= 36'sb100000000001010011010110100100101010;
            sine_reg0   <= 36'sb1001001000001101100101110101101;
        end
        8100: begin
            cosine_reg0 <= 36'sb100000000001010001100100011110101100;
            sine_reg0   <= 36'sb1001000001111011101110000110100;
        end
        8101: begin
            cosine_reg0 <= 36'sb100000000001001111110011100111100111;
            sine_reg0   <= 36'sb1000111011101001110110000001001;
        end
        8102: begin
            cosine_reg0 <= 36'sb100000000001001110000011111111011101;
            sine_reg0   <= 36'sb1000110101010111111101100101101;
        end
        8103: begin
            cosine_reg0 <= 36'sb100000000001001100010101100110001101;
            sine_reg0   <= 36'sb1000101111000110000100110100011;
        end
        8104: begin
            cosine_reg0 <= 36'sb100000000001001010101000011011111000;
            sine_reg0   <= 36'sb1000101000110100001011101101101;
        end
        8105: begin
            cosine_reg0 <= 36'sb100000000001001000111100100000011100;
            sine_reg0   <= 36'sb1000100010100010010010010001100;
        end
        8106: begin
            cosine_reg0 <= 36'sb100000000001000111010001110011111011;
            sine_reg0   <= 36'sb1000011100010000011000100000011;
        end
        8107: begin
            cosine_reg0 <= 36'sb100000000001000101101000010110010101;
            sine_reg0   <= 36'sb1000010101111110011110011010011;
        end
        8108: begin
            cosine_reg0 <= 36'sb100000000001000100000000000111101001;
            sine_reg0   <= 36'sb1000001111101100100011111111110;
        end
        8109: begin
            cosine_reg0 <= 36'sb100000000001000010011001000111111000;
            sine_reg0   <= 36'sb1000001001011010101001010000111;
        end
        8110: begin
            cosine_reg0 <= 36'sb100000000001000000110011010111000001;
            sine_reg0   <= 36'sb1000000011001000101110001101111;
        end
        8111: begin
            cosine_reg0 <= 36'sb100000000000111111001110110101000110;
            sine_reg0   <= 36'sb111111100110110110010110111000;
        end
        8112: begin
            cosine_reg0 <= 36'sb100000000000111101101011100010000101;
            sine_reg0   <= 36'sb111110110100100110111001100100;
        end
        8113: begin
            cosine_reg0 <= 36'sb100000000000111100001001011101111110;
            sine_reg0   <= 36'sb111110000010010111011001110101;
        end
        8114: begin
            cosine_reg0 <= 36'sb100000000000111010101000101000110011;
            sine_reg0   <= 36'sb111101010000000111110111101100;
        end
        8115: begin
            cosine_reg0 <= 36'sb100000000000111001001001000010100011;
            sine_reg0   <= 36'sb111100011101111000010011001101;
        end
        8116: begin
            cosine_reg0 <= 36'sb100000000000110111101010101011001110;
            sine_reg0   <= 36'sb111011101011101000101100011001;
        end
        8117: begin
            cosine_reg0 <= 36'sb100000000000110110001101100010110100;
            sine_reg0   <= 36'sb111010111001011001000011010001;
        end
        8118: begin
            cosine_reg0 <= 36'sb100000000000110100110001101001010101;
            sine_reg0   <= 36'sb111010000111001001010111111000;
        end
        8119: begin
            cosine_reg0 <= 36'sb100000000000110011010110111110110001;
            sine_reg0   <= 36'sb111001010100111001101010010000;
        end
        8120: begin
            cosine_reg0 <= 36'sb100000000000110001111101100011001000;
            sine_reg0   <= 36'sb111000100010101001111010011010;
        end
        8121: begin
            cosine_reg0 <= 36'sb100000000000110000100101010110011011;
            sine_reg0   <= 36'sb110111110000011010001000011000;
        end
        8122: begin
            cosine_reg0 <= 36'sb100000000000101111001110011000101001;
            sine_reg0   <= 36'sb110110111110001010010100001101;
        end
        8123: begin
            cosine_reg0 <= 36'sb100000000000101101111000101001110011;
            sine_reg0   <= 36'sb110110001011111010011101111011;
        end
        8124: begin
            cosine_reg0 <= 36'sb100000000000101100100100001001111000;
            sine_reg0   <= 36'sb110101011001101010100101100011;
        end
        8125: begin
            cosine_reg0 <= 36'sb100000000000101011010000111000111000;
            sine_reg0   <= 36'sb110100100111011010101011000111;
        end
        8126: begin
            cosine_reg0 <= 36'sb100000000000101001111110110110110101;
            sine_reg0   <= 36'sb110011110101001010101110101001;
        end
        8127: begin
            cosine_reg0 <= 36'sb100000000000101000101110000011101100;
            sine_reg0   <= 36'sb110011000010111010110000001011;
        end
        8128: begin
            cosine_reg0 <= 36'sb100000000000100111011110011111100000;
            sine_reg0   <= 36'sb110010010000101010101111101111;
        end
        8129: begin
            cosine_reg0 <= 36'sb100000000000100110010000001010001111;
            sine_reg0   <= 36'sb110001011110011010101101011000;
        end
        8130: begin
            cosine_reg0 <= 36'sb100000000000100101000011000011111010;
            sine_reg0   <= 36'sb110000101100001010101001000110;
        end
        8131: begin
            cosine_reg0 <= 36'sb100000000000100011110111001100100001;
            sine_reg0   <= 36'sb101111111001111010100010111100;
        end
        8132: begin
            cosine_reg0 <= 36'sb100000000000100010101100100100000011;
            sine_reg0   <= 36'sb101111000111101010011010111100;
        end
        8133: begin
            cosine_reg0 <= 36'sb100000000000100001100011001010100010;
            sine_reg0   <= 36'sb101110010101011010010001000111;
        end
        8134: begin
            cosine_reg0 <= 36'sb100000000000100000011010111111111100;
            sine_reg0   <= 36'sb101101100011001010000101100001;
        end
        8135: begin
            cosine_reg0 <= 36'sb100000000000011111010100000100010010;
            sine_reg0   <= 36'sb101100110000111001111000001001;
        end
        8136: begin
            cosine_reg0 <= 36'sb100000000000011110001110010111100101;
            sine_reg0   <= 36'sb101011111110101001101001000100;
        end
        8137: begin
            cosine_reg0 <= 36'sb100000000000011101001001111001110011;
            sine_reg0   <= 36'sb101011001100011001011000010010;
        end
        8138: begin
            cosine_reg0 <= 36'sb100000000000011100000110101010111110;
            sine_reg0   <= 36'sb101010011010001001000101110101;
        end
        8139: begin
            cosine_reg0 <= 36'sb100000000000011011000100101011000101;
            sine_reg0   <= 36'sb101001100111111000110001110000;
        end
        8140: begin
            cosine_reg0 <= 36'sb100000000000011010000011111010001000;
            sine_reg0   <= 36'sb101000110101101000011100000100;
        end
        8141: begin
            cosine_reg0 <= 36'sb100000000000011001000100011000000111;
            sine_reg0   <= 36'sb101000000011011000000100110011;
        end
        8142: begin
            cosine_reg0 <= 36'sb100000000000011000000110000101000010;
            sine_reg0   <= 36'sb100111010001000111101100000000;
        end
        8143: begin
            cosine_reg0 <= 36'sb100000000000010111001001000000111010;
            sine_reg0   <= 36'sb100110011110110111010001101011;
        end
        8144: begin
            cosine_reg0 <= 36'sb100000000000010110001101001011101110;
            sine_reg0   <= 36'sb100101101100100110110101111000;
        end
        8145: begin
            cosine_reg0 <= 36'sb100000000000010101010010100101011111;
            sine_reg0   <= 36'sb100100111010010110011000100111;
        end
        8146: begin
            cosine_reg0 <= 36'sb100000000000010100011001001110001100;
            sine_reg0   <= 36'sb100100001000000101111001111100;
        end
        8147: begin
            cosine_reg0 <= 36'sb100000000000010011100001000101110101;
            sine_reg0   <= 36'sb100011010101110101011001110111;
        end
        8148: begin
            cosine_reg0 <= 36'sb100000000000010010101010001100011011;
            sine_reg0   <= 36'sb100010100011100100111000011011;
        end
        8149: begin
            cosine_reg0 <= 36'sb100000000000010001110100100001111101;
            sine_reg0   <= 36'sb100001110001010100010101101010;
        end
        8150: begin
            cosine_reg0 <= 36'sb100000000000010001000000000110011100;
            sine_reg0   <= 36'sb100000111111000011110001100110;
        end
        8151: begin
            cosine_reg0 <= 36'sb100000000000010000001100111001111000;
            sine_reg0   <= 36'sb100000001100110011001100010000;
        end
        8152: begin
            cosine_reg0 <= 36'sb100000000000001111011010111100010000;
            sine_reg0   <= 36'sb11111011010100010100101101011;
        end
        8153: begin
            cosine_reg0 <= 36'sb100000000000001110101010001101100100;
            sine_reg0   <= 36'sb11110101000010001111101111000;
        end
        8154: begin
            cosine_reg0 <= 36'sb100000000000001101111010101101110110;
            sine_reg0   <= 36'sb11101110110000001010100111010;
        end
        8155: begin
            cosine_reg0 <= 36'sb100000000000001101001100011101000100;
            sine_reg0   <= 36'sb11101000011110000101010110010;
        end
        8156: begin
            cosine_reg0 <= 36'sb100000000000001100011111011011001111;
            sine_reg0   <= 36'sb11100010001011111111111100010;
        end
        8157: begin
            cosine_reg0 <= 36'sb100000000000001011110011101000010110;
            sine_reg0   <= 36'sb11011011111001111010011001100;
        end
        8158: begin
            cosine_reg0 <= 36'sb100000000000001011001001000100011011;
            sine_reg0   <= 36'sb11010101100111110100101110011;
        end
        8159: begin
            cosine_reg0 <= 36'sb100000000000001010011111101111011100;
            sine_reg0   <= 36'sb11001111010101101110111011000;
        end
        8160: begin
            cosine_reg0 <= 36'sb100000000000001001110111101001011010;
            sine_reg0   <= 36'sb11001001000011101000111111101;
        end
        8161: begin
            cosine_reg0 <= 36'sb100000000000001001010000110010010101;
            sine_reg0   <= 36'sb11000010110001100010111100100;
        end
        8162: begin
            cosine_reg0 <= 36'sb100000000000001000101011001010001101;
            sine_reg0   <= 36'sb10111100011111011100110001111;
        end
        8163: begin
            cosine_reg0 <= 36'sb100000000000001000000110110001000001;
            sine_reg0   <= 36'sb10110110001101010110011111111;
        end
        8164: begin
            cosine_reg0 <= 36'sb100000000000000111100011100110110011;
            sine_reg0   <= 36'sb10101111111011010000000111000;
        end
        8165: begin
            cosine_reg0 <= 36'sb100000000000000111000001101011100010;
            sine_reg0   <= 36'sb10101001101001001001100111010;
        end
        8166: begin
            cosine_reg0 <= 36'sb100000000000000110100000111111001101;
            sine_reg0   <= 36'sb10100011010111000011000001000;
        end
        8167: begin
            cosine_reg0 <= 36'sb100000000000000110000001100001110110;
            sine_reg0   <= 36'sb10011101000100111100010100011;
        end
        8168: begin
            cosine_reg0 <= 36'sb100000000000000101100011010011011011;
            sine_reg0   <= 36'sb10010110110010110101100001110;
        end
        8169: begin
            cosine_reg0 <= 36'sb100000000000000101000110010011111110;
            sine_reg0   <= 36'sb10010000100000101110101001011;
        end
        8170: begin
            cosine_reg0 <= 36'sb100000000000000100101010100011011101;
            sine_reg0   <= 36'sb10001010001110100111101011011;
        end
        8171: begin
            cosine_reg0 <= 36'sb100000000000000100010000000001111010;
            sine_reg0   <= 36'sb10000011111100100000101000000;
        end
        8172: begin
            cosine_reg0 <= 36'sb100000000000000011110110101111010100;
            sine_reg0   <= 36'sb1111101101010011001011111101;
        end
        8173: begin
            cosine_reg0 <= 36'sb100000000000000011011110101011101010;
            sine_reg0   <= 36'sb1110111011000010010010010011;
        end
        8174: begin
            cosine_reg0 <= 36'sb100000000000000011000111110110111110;
            sine_reg0   <= 36'sb1110001000110001011000000100;
        end
        8175: begin
            cosine_reg0 <= 36'sb100000000000000010110010010001001111;
            sine_reg0   <= 36'sb1101010110100000011101010010;
        end
        8176: begin
            cosine_reg0 <= 36'sb100000000000000010011101111010011101;
            sine_reg0   <= 36'sb1100100100001111100001111111;
        end
        8177: begin
            cosine_reg0 <= 36'sb100000000000000010001010110010101001;
            sine_reg0   <= 36'sb1011110001111110100110001101;
        end
        8178: begin
            cosine_reg0 <= 36'sb100000000000000001111000111001110001;
            sine_reg0   <= 36'sb1010111111101101101001111111;
        end
        8179: begin
            cosine_reg0 <= 36'sb100000000000000001101000001111110111;
            sine_reg0   <= 36'sb1010001101011100101101010101;
        end
        8180: begin
            cosine_reg0 <= 36'sb100000000000000001011000110100111001;
            sine_reg0   <= 36'sb1001011011001011110000010001;
        end
        8181: begin
            cosine_reg0 <= 36'sb100000000000000001001010101000111001;
            sine_reg0   <= 36'sb1000101000111010110010110111;
        end
        8182: begin
            cosine_reg0 <= 36'sb100000000000000000111101101011110111;
            sine_reg0   <= 36'sb111110110101001110101000111;
        end
        8183: begin
            cosine_reg0 <= 36'sb100000000000000000110001111101110001;
            sine_reg0   <= 36'sb111000100011000110111000100;
        end
        8184: begin
            cosine_reg0 <= 36'sb100000000000000000100111011110101000;
            sine_reg0   <= 36'sb110010010000111111000110000;
        end
        8185: begin
            cosine_reg0 <= 36'sb100000000000000000011110001110011101;
            sine_reg0   <= 36'sb101011111110110111010001100;
        end
        8186: begin
            cosine_reg0 <= 36'sb100000000000000000010110001101001111;
            sine_reg0   <= 36'sb100101101100101111011011010;
        end
        8187: begin
            cosine_reg0 <= 36'sb100000000000000000001111011010111110;
            sine_reg0   <= 36'sb11111011010100111100011101;
        end
        8188: begin
            cosine_reg0 <= 36'sb100000000000000000001001110111101011;
            sine_reg0   <= 36'sb11001001000011111101010110;
        end
        8189: begin
            cosine_reg0 <= 36'sb100000000000000000000101100011010101;
            sine_reg0   <= 36'sb10010110110010111110000111;
        end
        8190: begin
            cosine_reg0 <= 36'sb100000000000000000000010011101111011;
            sine_reg0   <= 36'sb1100100100001111110110011;
        end
        8191: begin
            cosine_reg0 <= 36'sb100000000000000000000000100111100000;
            sine_reg0   <= 36'sb110010010000111111011010;
        end
        8192: begin
            cosine_reg0 <= 36'sb100000000000000000000000000000000001;
            sine_reg0   <= 36'sb0;
        end
        8193: begin
            cosine_reg0 <= 36'sb100000000000000000000000100111100000;
            sine_reg0   <= 36'sb111111111111001101101111000000100110;
        end
        8194: begin
            cosine_reg0 <= 36'sb100000000000000000000010011101111011;
            sine_reg0   <= 36'sb111111111110011011011110000001001101;
        end
        8195: begin
            cosine_reg0 <= 36'sb100000000000000000000101100011010101;
            sine_reg0   <= 36'sb111111111101101001001101000001111001;
        end
        8196: begin
            cosine_reg0 <= 36'sb100000000000000000001001110111101011;
            sine_reg0   <= 36'sb111111111100110110111100000010101010;
        end
        8197: begin
            cosine_reg0 <= 36'sb100000000000000000001111011010111110;
            sine_reg0   <= 36'sb111111111100000100101011000011100011;
        end
        8198: begin
            cosine_reg0 <= 36'sb100000000000000000010110001101001111;
            sine_reg0   <= 36'sb111111111011010010011010000100100110;
        end
        8199: begin
            cosine_reg0 <= 36'sb100000000000000000011110001110011101;
            sine_reg0   <= 36'sb111111111010100000001001000101110100;
        end
        8200: begin
            cosine_reg0 <= 36'sb100000000000000000100111011110101000;
            sine_reg0   <= 36'sb111111111001101101111000000111010000;
        end
        8201: begin
            cosine_reg0 <= 36'sb100000000000000000110001111101110001;
            sine_reg0   <= 36'sb111111111000111011100111001000111100;
        end
        8202: begin
            cosine_reg0 <= 36'sb100000000000000000111101101011110111;
            sine_reg0   <= 36'sb111111111000001001010110001010111001;
        end
        8203: begin
            cosine_reg0 <= 36'sb100000000000000001001010101000111001;
            sine_reg0   <= 36'sb111111110111010111000101001101001001;
        end
        8204: begin
            cosine_reg0 <= 36'sb100000000000000001011000110100111001;
            sine_reg0   <= 36'sb111111110110100100110100001111101111;
        end
        8205: begin
            cosine_reg0 <= 36'sb100000000000000001101000001111110111;
            sine_reg0   <= 36'sb111111110101110010100011010010101011;
        end
        8206: begin
            cosine_reg0 <= 36'sb100000000000000001111000111001110001;
            sine_reg0   <= 36'sb111111110101000000010010010110000001;
        end
        8207: begin
            cosine_reg0 <= 36'sb100000000000000010001010110010101001;
            sine_reg0   <= 36'sb111111110100001110000001011001110011;
        end
        8208: begin
            cosine_reg0 <= 36'sb100000000000000010011101111010011101;
            sine_reg0   <= 36'sb111111110011011011110000011110000001;
        end
        8209: begin
            cosine_reg0 <= 36'sb100000000000000010110010010001001111;
            sine_reg0   <= 36'sb111111110010101001011111100010101110;
        end
        8210: begin
            cosine_reg0 <= 36'sb100000000000000011000111110110111110;
            sine_reg0   <= 36'sb111111110001110111001110100111111100;
        end
        8211: begin
            cosine_reg0 <= 36'sb100000000000000011011110101011101010;
            sine_reg0   <= 36'sb111111110001000100111101101101101101;
        end
        8212: begin
            cosine_reg0 <= 36'sb100000000000000011110110101111010100;
            sine_reg0   <= 36'sb111111110000010010101100110100000011;
        end
        8213: begin
            cosine_reg0 <= 36'sb100000000000000100010000000001111010;
            sine_reg0   <= 36'sb111111101111100000011011111011000000;
        end
        8214: begin
            cosine_reg0 <= 36'sb100000000000000100101010100011011101;
            sine_reg0   <= 36'sb111111101110101110001011000010100101;
        end
        8215: begin
            cosine_reg0 <= 36'sb100000000000000101000110010011111110;
            sine_reg0   <= 36'sb111111101101111011111010001010110101;
        end
        8216: begin
            cosine_reg0 <= 36'sb100000000000000101100011010011011011;
            sine_reg0   <= 36'sb111111101101001001101001010011110010;
        end
        8217: begin
            cosine_reg0 <= 36'sb100000000000000110000001100001110110;
            sine_reg0   <= 36'sb111111101100010111011000011101011101;
        end
        8218: begin
            cosine_reg0 <= 36'sb100000000000000110100000111111001101;
            sine_reg0   <= 36'sb111111101011100101000111100111111000;
        end
        8219: begin
            cosine_reg0 <= 36'sb100000000000000111000001101011100010;
            sine_reg0   <= 36'sb111111101010110010110110110011000110;
        end
        8220: begin
            cosine_reg0 <= 36'sb100000000000000111100011100110110011;
            sine_reg0   <= 36'sb111111101010000000100101111111001000;
        end
        8221: begin
            cosine_reg0 <= 36'sb100000000000001000000110110001000001;
            sine_reg0   <= 36'sb111111101001001110010101001100000001;
        end
        8222: begin
            cosine_reg0 <= 36'sb100000000000001000101011001010001101;
            sine_reg0   <= 36'sb111111101000011100000100011001110001;
        end
        8223: begin
            cosine_reg0 <= 36'sb100000000000001001010000110010010101;
            sine_reg0   <= 36'sb111111100111101001110011101000011100;
        end
        8224: begin
            cosine_reg0 <= 36'sb100000000000001001110111101001011010;
            sine_reg0   <= 36'sb111111100110110111100010111000000011;
        end
        8225: begin
            cosine_reg0 <= 36'sb100000000000001010011111101111011100;
            sine_reg0   <= 36'sb111111100110000101010010001000101000;
        end
        8226: begin
            cosine_reg0 <= 36'sb100000000000001011001001000100011011;
            sine_reg0   <= 36'sb111111100101010011000001011010001101;
        end
        8227: begin
            cosine_reg0 <= 36'sb100000000000001011110011101000010110;
            sine_reg0   <= 36'sb111111100100100000110000101100110100;
        end
        8228: begin
            cosine_reg0 <= 36'sb100000000000001100011111011011001111;
            sine_reg0   <= 36'sb111111100011101110100000000000011110;
        end
        8229: begin
            cosine_reg0 <= 36'sb100000000000001101001100011101000100;
            sine_reg0   <= 36'sb111111100010111100001111010101001110;
        end
        8230: begin
            cosine_reg0 <= 36'sb100000000000001101111010101101110110;
            sine_reg0   <= 36'sb111111100010001001111110101011000110;
        end
        8231: begin
            cosine_reg0 <= 36'sb100000000000001110101010001101100100;
            sine_reg0   <= 36'sb111111100001010111101110000010001000;
        end
        8232: begin
            cosine_reg0 <= 36'sb100000000000001111011010111100010000;
            sine_reg0   <= 36'sb111111100000100101011101011010010101;
        end
        8233: begin
            cosine_reg0 <= 36'sb100000000000010000001100111001111000;
            sine_reg0   <= 36'sb111111011111110011001100110011110000;
        end
        8234: begin
            cosine_reg0 <= 36'sb100000000000010001000000000110011100;
            sine_reg0   <= 36'sb111111011111000000111100001110011010;
        end
        8235: begin
            cosine_reg0 <= 36'sb100000000000010001110100100001111101;
            sine_reg0   <= 36'sb111111011110001110101011101010010110;
        end
        8236: begin
            cosine_reg0 <= 36'sb100000000000010010101010001100011011;
            sine_reg0   <= 36'sb111111011101011100011011000111100101;
        end
        8237: begin
            cosine_reg0 <= 36'sb100000000000010011100001000101110101;
            sine_reg0   <= 36'sb111111011100101010001010100110001001;
        end
        8238: begin
            cosine_reg0 <= 36'sb100000000000010100011001001110001100;
            sine_reg0   <= 36'sb111111011011110111111010000110000100;
        end
        8239: begin
            cosine_reg0 <= 36'sb100000000000010101010010100101011111;
            sine_reg0   <= 36'sb111111011011000101101001100111011001;
        end
        8240: begin
            cosine_reg0 <= 36'sb100000000000010110001101001011101110;
            sine_reg0   <= 36'sb111111011010010011011001001010001000;
        end
        8241: begin
            cosine_reg0 <= 36'sb100000000000010111001001000000111010;
            sine_reg0   <= 36'sb111111011001100001001000101110010101;
        end
        8242: begin
            cosine_reg0 <= 36'sb100000000000011000000110000101000010;
            sine_reg0   <= 36'sb111111011000101110111000010100000000;
        end
        8243: begin
            cosine_reg0 <= 36'sb100000000000011001000100011000000111;
            sine_reg0   <= 36'sb111111010111111100100111111011001101;
        end
        8244: begin
            cosine_reg0 <= 36'sb100000000000011010000011111010001000;
            sine_reg0   <= 36'sb111111010111001010010111100011111100;
        end
        8245: begin
            cosine_reg0 <= 36'sb100000000000011011000100101011000101;
            sine_reg0   <= 36'sb111111010110011000000111001110010000;
        end
        8246: begin
            cosine_reg0 <= 36'sb100000000000011100000110101010111110;
            sine_reg0   <= 36'sb111111010101100101110110111010001011;
        end
        8247: begin
            cosine_reg0 <= 36'sb100000000000011101001001111001110011;
            sine_reg0   <= 36'sb111111010100110011100110100111101110;
        end
        8248: begin
            cosine_reg0 <= 36'sb100000000000011110001110010111100101;
            sine_reg0   <= 36'sb111111010100000001010110010110111100;
        end
        8249: begin
            cosine_reg0 <= 36'sb100000000000011111010100000100010010;
            sine_reg0   <= 36'sb111111010011001111000110000111110111;
        end
        8250: begin
            cosine_reg0 <= 36'sb100000000000100000011010111111111100;
            sine_reg0   <= 36'sb111111010010011100110101111010011111;
        end
        8251: begin
            cosine_reg0 <= 36'sb100000000000100001100011001010100010;
            sine_reg0   <= 36'sb111111010001101010100101101110111001;
        end
        8252: begin
            cosine_reg0 <= 36'sb100000000000100010101100100100000011;
            sine_reg0   <= 36'sb111111010000111000010101100101000100;
        end
        8253: begin
            cosine_reg0 <= 36'sb100000000000100011110111001100100001;
            sine_reg0   <= 36'sb111111010000000110000101011101000100;
        end
        8254: begin
            cosine_reg0 <= 36'sb100000000000100101000011000011111010;
            sine_reg0   <= 36'sb111111001111010011110101010110111010;
        end
        8255: begin
            cosine_reg0 <= 36'sb100000000000100110010000001010001111;
            sine_reg0   <= 36'sb111111001110100001100101010010101000;
        end
        8256: begin
            cosine_reg0 <= 36'sb100000000000100111011110011111100000;
            sine_reg0   <= 36'sb111111001101101111010101010000010001;
        end
        8257: begin
            cosine_reg0 <= 36'sb100000000000101000101110000011101100;
            sine_reg0   <= 36'sb111111001100111101000101001111110101;
        end
        8258: begin
            cosine_reg0 <= 36'sb100000000000101001111110110110110101;
            sine_reg0   <= 36'sb111111001100001010110101010001010111;
        end
        8259: begin
            cosine_reg0 <= 36'sb100000000000101011010000111000111000;
            sine_reg0   <= 36'sb111111001011011000100101010100111001;
        end
        8260: begin
            cosine_reg0 <= 36'sb100000000000101100100100001001111000;
            sine_reg0   <= 36'sb111111001010100110010101011010011101;
        end
        8261: begin
            cosine_reg0 <= 36'sb100000000000101101111000101001110011;
            sine_reg0   <= 36'sb111111001001110100000101100010000101;
        end
        8262: begin
            cosine_reg0 <= 36'sb100000000000101111001110011000101001;
            sine_reg0   <= 36'sb111111001001000001110101101011110011;
        end
        8263: begin
            cosine_reg0 <= 36'sb100000000000110000100101010110011011;
            sine_reg0   <= 36'sb111111001000001111100101110111101000;
        end
        8264: begin
            cosine_reg0 <= 36'sb100000000000110001111101100011001000;
            sine_reg0   <= 36'sb111111000111011101010110000101100110;
        end
        8265: begin
            cosine_reg0 <= 36'sb100000000000110011010110111110110001;
            sine_reg0   <= 36'sb111111000110101011000110010101110000;
        end
        8266: begin
            cosine_reg0 <= 36'sb100000000000110100110001101001010101;
            sine_reg0   <= 36'sb111111000101111000110110101000001000;
        end
        8267: begin
            cosine_reg0 <= 36'sb100000000000110110001101100010110100;
            sine_reg0   <= 36'sb111111000101000110100110111100101111;
        end
        8268: begin
            cosine_reg0 <= 36'sb100000000000110111101010101011001110;
            sine_reg0   <= 36'sb111111000100010100010111010011100111;
        end
        8269: begin
            cosine_reg0 <= 36'sb100000000000111001001001000010100011;
            sine_reg0   <= 36'sb111111000011100010000111101100110011;
        end
        8270: begin
            cosine_reg0 <= 36'sb100000000000111010101000101000110011;
            sine_reg0   <= 36'sb111111000010101111111000001000010100;
        end
        8271: begin
            cosine_reg0 <= 36'sb100000000000111100001001011101111110;
            sine_reg0   <= 36'sb111111000001111101101000100110001011;
        end
        8272: begin
            cosine_reg0 <= 36'sb100000000000111101101011100010000101;
            sine_reg0   <= 36'sb111111000001001011011001000110011100;
        end
        8273: begin
            cosine_reg0 <= 36'sb100000000000111111001110110101000110;
            sine_reg0   <= 36'sb111111000000011001001001101001001000;
        end
        8274: begin
            cosine_reg0 <= 36'sb100000000001000000110011010111000001;
            sine_reg0   <= 36'sb111110111111100110111010001110010001;
        end
        8275: begin
            cosine_reg0 <= 36'sb100000000001000010011001000111111000;
            sine_reg0   <= 36'sb111110111110110100101010110101111001;
        end
        8276: begin
            cosine_reg0 <= 36'sb100000000001000100000000000111101001;
            sine_reg0   <= 36'sb111110111110000010011011100000000010;
        end
        8277: begin
            cosine_reg0 <= 36'sb100000000001000101101000010110010101;
            sine_reg0   <= 36'sb111110111101010000001100001100101101;
        end
        8278: begin
            cosine_reg0 <= 36'sb100000000001000111010001110011111011;
            sine_reg0   <= 36'sb111110111100011101111100111011111101;
        end
        8279: begin
            cosine_reg0 <= 36'sb100000000001001000111100100000011100;
            sine_reg0   <= 36'sb111110111011101011101101101101110100;
        end
        8280: begin
            cosine_reg0 <= 36'sb100000000001001010101000011011111000;
            sine_reg0   <= 36'sb111110111010111001011110100010010011;
        end
        8281: begin
            cosine_reg0 <= 36'sb100000000001001100010101100110001101;
            sine_reg0   <= 36'sb111110111010000111001111011001011101;
        end
        8282: begin
            cosine_reg0 <= 36'sb100000000001001110000011111111011101;
            sine_reg0   <= 36'sb111110111001010101000000010011010011;
        end
        8283: begin
            cosine_reg0 <= 36'sb100000000001001111110011100111100111;
            sine_reg0   <= 36'sb111110111000100010110001001111110111;
        end
        8284: begin
            cosine_reg0 <= 36'sb100000000001010001100100011110101100;
            sine_reg0   <= 36'sb111110110111110000100010001111001100;
        end
        8285: begin
            cosine_reg0 <= 36'sb100000000001010011010110100100101010;
            sine_reg0   <= 36'sb111110110110111110010011010001010011;
        end
        8286: begin
            cosine_reg0 <= 36'sb100000000001010101001001111001100011;
            sine_reg0   <= 36'sb111110110110001100000100010110001111;
        end
        8287: begin
            cosine_reg0 <= 36'sb100000000001010110111110011101010101;
            sine_reg0   <= 36'sb111110110101011001110101011110000000;
        end
        8288: begin
            cosine_reg0 <= 36'sb100000000001011000110100010000000001;
            sine_reg0   <= 36'sb111110110100100111100110101000101010;
        end
        8289: begin
            cosine_reg0 <= 36'sb100000000001011010101011010001100111;
            sine_reg0   <= 36'sb111110110011110101010111110110001101;
        end
        8290: begin
            cosine_reg0 <= 36'sb100000000001011100100011100010000111;
            sine_reg0   <= 36'sb111110110011000011001001000110101101;
        end
        8291: begin
            cosine_reg0 <= 36'sb100000000001011110011101000001100001;
            sine_reg0   <= 36'sb111110110010010000111010011010001010;
        end
        8292: begin
            cosine_reg0 <= 36'sb100000000001100000010111101111110100;
            sine_reg0   <= 36'sb111110110001011110101011110000100111;
        end
        8293: begin
            cosine_reg0 <= 36'sb100000000001100010010011101101000001;
            sine_reg0   <= 36'sb111110110000101100011101001010000110;
        end
        8294: begin
            cosine_reg0 <= 36'sb100000000001100100010000111001000111;
            sine_reg0   <= 36'sb111110101111111010001110100110101000;
        end
        8295: begin
            cosine_reg0 <= 36'sb100000000001100110001111010100000110;
            sine_reg0   <= 36'sb111110101111001000000000000110010000;
        end
        8296: begin
            cosine_reg0 <= 36'sb100000000001101000001110111101111111;
            sine_reg0   <= 36'sb111110101110010101110001101001000000;
        end
        8297: begin
            cosine_reg0 <= 36'sb100000000001101010001111110110110001;
            sine_reg0   <= 36'sb111110101101100011100011001110111001;
        end
        8298: begin
            cosine_reg0 <= 36'sb100000000001101100010001111110011100;
            sine_reg0   <= 36'sb111110101100110001010100110111111110;
        end
        8299: begin
            cosine_reg0 <= 36'sb100000000001101110010101010101000000;
            sine_reg0   <= 36'sb111110101011111111000110100100010000;
        end
        8300: begin
            cosine_reg0 <= 36'sb100000000001110000011001111010011101;
            sine_reg0   <= 36'sb111110101011001100111000010011110001;
        end
        8301: begin
            cosine_reg0 <= 36'sb100000000001110010011111101110110011;
            sine_reg0   <= 36'sb111110101010011010101010000110100100;
        end
        8302: begin
            cosine_reg0 <= 36'sb100000000001110100100110110010000010;
            sine_reg0   <= 36'sb111110101001101000011011111100101001;
        end
        8303: begin
            cosine_reg0 <= 36'sb100000000001110110101111000100001010;
            sine_reg0   <= 36'sb111110101000110110001101110110000100;
        end
        8304: begin
            cosine_reg0 <= 36'sb100000000001111000111000100101001010;
            sine_reg0   <= 36'sb111110101000000011111111110010110110;
        end
        8305: begin
            cosine_reg0 <= 36'sb100000000001111011000011010101000011;
            sine_reg0   <= 36'sb111110100111010001110001110011000001;
        end
        8306: begin
            cosine_reg0 <= 36'sb100000000001111101001111010011110100;
            sine_reg0   <= 36'sb111110100110011111100011110110100110;
        end
        8307: begin
            cosine_reg0 <= 36'sb100000000001111111011100100001011110;
            sine_reg0   <= 36'sb111110100101101101010101111101101001;
        end
        8308: begin
            cosine_reg0 <= 36'sb100000000010000001101010111110000000;
            sine_reg0   <= 36'sb111110100100111011001000001000001010;
        end
        8309: begin
            cosine_reg0 <= 36'sb100000000010000011111010101001011011;
            sine_reg0   <= 36'sb111110100100001000111010010110001100;
        end
        8310: begin
            cosine_reg0 <= 36'sb100000000010000110001011100011101101;
            sine_reg0   <= 36'sb111110100011010110101100100111110001;
        end
        8311: begin
            cosine_reg0 <= 36'sb100000000010001000011101101100111000;
            sine_reg0   <= 36'sb111110100010100100011110111100111010;
        end
        8312: begin
            cosine_reg0 <= 36'sb100000000010001010110001000100111010;
            sine_reg0   <= 36'sb111110100001110010010001010101101010;
        end
        8313: begin
            cosine_reg0 <= 36'sb100000000010001101000101101011110101;
            sine_reg0   <= 36'sb111110100001000000000011110010000010;
        end
        8314: begin
            cosine_reg0 <= 36'sb100000000010001111011011100001100111;
            sine_reg0   <= 36'sb111110100000001101110110010010000101;
        end
        8315: begin
            cosine_reg0 <= 36'sb100000000010010001110010100110010001;
            sine_reg0   <= 36'sb111110011111011011101000110101110100;
        end
        8316: begin
            cosine_reg0 <= 36'sb100000000010010100001010111001110010;
            sine_reg0   <= 36'sb111110011110101001011011011101010001;
        end
        8317: begin
            cosine_reg0 <= 36'sb100000000010010110100100011100001011;
            sine_reg0   <= 36'sb111110011101110111001110001000011111;
        end
        8318: begin
            cosine_reg0 <= 36'sb100000000010011000111111001101011100;
            sine_reg0   <= 36'sb111110011101000101000000110111011110;
        end
        8319: begin
            cosine_reg0 <= 36'sb100000000010011011011011001101100100;
            sine_reg0   <= 36'sb111110011100010010110011101010010010;
        end
        8320: begin
            cosine_reg0 <= 36'sb100000000010011101111000011100100011;
            sine_reg0   <= 36'sb111110011011100000100110100000111100;
        end
        8321: begin
            cosine_reg0 <= 36'sb100000000010100000010110111010011001;
            sine_reg0   <= 36'sb111110011010101110011001011011011110;
        end
        8322: begin
            cosine_reg0 <= 36'sb100000000010100010110110100111000110;
            sine_reg0   <= 36'sb111110011001111100001100011001111001;
        end
        8323: begin
            cosine_reg0 <= 36'sb100000000010100101010111100010101010;
            sine_reg0   <= 36'sb111110011001001001111111011100010001;
        end
        8324: begin
            cosine_reg0 <= 36'sb100000000010100111111001101101000101;
            sine_reg0   <= 36'sb111110011000010111110010100010100110;
        end
        8325: begin
            cosine_reg0 <= 36'sb100000000010101010011101000110010111;
            sine_reg0   <= 36'sb111110010111100101100101101100111011;
        end
        8326: begin
            cosine_reg0 <= 36'sb100000000010101101000001101110100000;
            sine_reg0   <= 36'sb111110010110110011011000111011010001;
        end
        8327: begin
            cosine_reg0 <= 36'sb100000000010101111100111100101011111;
            sine_reg0   <= 36'sb111110010110000001001100001101101011;
        end
        8328: begin
            cosine_reg0 <= 36'sb100000000010110010001110101011010101;
            sine_reg0   <= 36'sb111110010101001110111111100100001011;
        end
        8329: begin
            cosine_reg0 <= 36'sb100000000010110100110111000000000000;
            sine_reg0   <= 36'sb111110010100011100110010111110110010;
        end
        8330: begin
            cosine_reg0 <= 36'sb100000000010110111100000100011100011;
            sine_reg0   <= 36'sb111110010011101010100110011101100010;
        end
        8331: begin
            cosine_reg0 <= 36'sb100000000010111010001011010101111011;
            sine_reg0   <= 36'sb111110010010111000011010000000011110;
        end
        8332: begin
            cosine_reg0 <= 36'sb100000000010111100110111010111001001;
            sine_reg0   <= 36'sb111110010010000110001101100111100110;
        end
        8333: begin
            cosine_reg0 <= 36'sb100000000010111111100100100111001110;
            sine_reg0   <= 36'sb111110010001010100000001010010111110;
        end
        8334: begin
            cosine_reg0 <= 36'sb100000000011000010010011000110001000;
            sine_reg0   <= 36'sb111110010000100001110101000010101000;
        end
        8335: begin
            cosine_reg0 <= 36'sb100000000011000101000010110011111000;
            sine_reg0   <= 36'sb111110001111101111101000110110100100;
        end
        8336: begin
            cosine_reg0 <= 36'sb100000000011000111110011110000011110;
            sine_reg0   <= 36'sb111110001110111101011100101110110101;
        end
        8337: begin
            cosine_reg0 <= 36'sb100000000011001010100101111011111001;
            sine_reg0   <= 36'sb111110001110001011010000101011011101;
        end
        8338: begin
            cosine_reg0 <= 36'sb100000000011001101011001010110001001;
            sine_reg0   <= 36'sb111110001101011001000100101100011110;
        end
        8339: begin
            cosine_reg0 <= 36'sb100000000011010000001101111111001111;
            sine_reg0   <= 36'sb111110001100100110111000110001111010;
        end
        8340: begin
            cosine_reg0 <= 36'sb100000000011010011000011110111001010;
            sine_reg0   <= 36'sb111110001011110100101100111011110010;
        end
        8341: begin
            cosine_reg0 <= 36'sb100000000011010101111010111101111011;
            sine_reg0   <= 36'sb111110001011000010100001001010001001;
        end
        8342: begin
            cosine_reg0 <= 36'sb100000000011011000110011010011100000;
            sine_reg0   <= 36'sb111110001010010000010101011101000001;
        end
        8343: begin
            cosine_reg0 <= 36'sb100000000011011011101100110111111010;
            sine_reg0   <= 36'sb111110001001011110001001110100011011;
        end
        8344: begin
            cosine_reg0 <= 36'sb100000000011011110100111101011001001;
            sine_reg0   <= 36'sb111110001000101011111110010000011010;
        end
        8345: begin
            cosine_reg0 <= 36'sb100000000011100001100011101101001100;
            sine_reg0   <= 36'sb111110000111111001110010110000111111;
        end
        8346: begin
            cosine_reg0 <= 36'sb100000000011100100100000111110000100;
            sine_reg0   <= 36'sb111110000111000111100111010110001101;
        end
        8347: begin
            cosine_reg0 <= 36'sb100000000011100111011111011101110001;
            sine_reg0   <= 36'sb111110000110010101011100000000000100;
        end
        8348: begin
            cosine_reg0 <= 36'sb100000000011101010011111001100010001;
            sine_reg0   <= 36'sb111110000101100011010000101110101000;
        end
        8349: begin
            cosine_reg0 <= 36'sb100000000011101101100000001001100110;
            sine_reg0   <= 36'sb111110000100110001000101100001111010;
        end
        8350: begin
            cosine_reg0 <= 36'sb100000000011110000100010010101110000;
            sine_reg0   <= 36'sb111110000011111110111010011001111100;
        end
        8351: begin
            cosine_reg0 <= 36'sb100000000011110011100101110000101101;
            sine_reg0   <= 36'sb111110000011001100101111010110110000;
        end
        8352: begin
            cosine_reg0 <= 36'sb100000000011110110101010011010011101;
            sine_reg0   <= 36'sb111110000010011010100100011000011000;
        end
        8353: begin
            cosine_reg0 <= 36'sb100000000011111001110000010011000010;
            sine_reg0   <= 36'sb111110000001101000011001011110110110;
        end
        8354: begin
            cosine_reg0 <= 36'sb100000000011111100110111011010011010;
            sine_reg0   <= 36'sb111110000000110110001110101010001100;
        end
        8355: begin
            cosine_reg0 <= 36'sb100000000011111111111111110000100110;
            sine_reg0   <= 36'sb111110000000000100000011111010011011;
        end
        8356: begin
            cosine_reg0 <= 36'sb100000000100000011001001010101100101;
            sine_reg0   <= 36'sb111101111111010001111001001111100110;
        end
        8357: begin
            cosine_reg0 <= 36'sb100000000100000110010100001001010111;
            sine_reg0   <= 36'sb111101111110011111101110101001101111;
        end
        8358: begin
            cosine_reg0 <= 36'sb100000000100001001100000001011111101;
            sine_reg0   <= 36'sb111101111101101101100100001000110111;
        end
        8359: begin
            cosine_reg0 <= 36'sb100000000100001100101101011101010101;
            sine_reg0   <= 36'sb111101111100111011011001101101000001;
        end
        8360: begin
            cosine_reg0 <= 36'sb100000000100001111111011111101100000;
            sine_reg0   <= 36'sb111101111100001001001111010110001110;
        end
        8361: begin
            cosine_reg0 <= 36'sb100000000100010011001011101100011110;
            sine_reg0   <= 36'sb111101111011010111000101000100100000;
        end
        8362: begin
            cosine_reg0 <= 36'sb100000000100010110011100101010001111;
            sine_reg0   <= 36'sb111101111010100100111010110111111010;
        end
        8363: begin
            cosine_reg0 <= 36'sb100000000100011001101110110110110010;
            sine_reg0   <= 36'sb111101111001110010110000110000011101;
        end
        8364: begin
            cosine_reg0 <= 36'sb100000000100011101000010010010001000;
            sine_reg0   <= 36'sb111101111001000000100110101110001011;
        end
        8365: begin
            cosine_reg0 <= 36'sb100000000100100000010110111100010000;
            sine_reg0   <= 36'sb111101111000001110011100110001000110;
        end
        8366: begin
            cosine_reg0 <= 36'sb100000000100100011101100110101001010;
            sine_reg0   <= 36'sb111101110111011100010010111001010000;
        end
        8367: begin
            cosine_reg0 <= 36'sb100000000100100111000011111100110110;
            sine_reg0   <= 36'sb111101110110101010001001000110101011;
        end
        8368: begin
            cosine_reg0 <= 36'sb100000000100101010011100010011010011;
            sine_reg0   <= 36'sb111101110101110111111111011001011001;
        end
        8369: begin
            cosine_reg0 <= 36'sb100000000100101101110101111000100011;
            sine_reg0   <= 36'sb111101110101000101110101110001011100;
        end
        8370: begin
            cosine_reg0 <= 36'sb100000000100110001010000101100100100;
            sine_reg0   <= 36'sb111101110100010011101100001110110110;
        end
        8371: begin
            cosine_reg0 <= 36'sb100000000100110100101100101111010111;
            sine_reg0   <= 36'sb111101110011100001100010110001101000;
        end
        8372: begin
            cosine_reg0 <= 36'sb100000000100111000001010000000111011;
            sine_reg0   <= 36'sb111101110010101111011001011001110101;
        end
        8373: begin
            cosine_reg0 <= 36'sb100000000100111011101000100001010000;
            sine_reg0   <= 36'sb111101110001111101010000000111011110;
        end
        8374: begin
            cosine_reg0 <= 36'sb100000000100111111001000010000010110;
            sine_reg0   <= 36'sb111101110001001011000110111010100110;
        end
        8375: begin
            cosine_reg0 <= 36'sb100000000101000010101001001110001101;
            sine_reg0   <= 36'sb111101110000011000111101110011001110;
        end
        8376: begin
            cosine_reg0 <= 36'sb100000000101000110001011011010110101;
            sine_reg0   <= 36'sb111101101111100110110100110001011001;
        end
        8377: begin
            cosine_reg0 <= 36'sb100000000101001001101110110110001110;
            sine_reg0   <= 36'sb111101101110110100101011110101001000;
        end
        8378: begin
            cosine_reg0 <= 36'sb100000000101001101010011100000010111;
            sine_reg0   <= 36'sb111101101110000010100010111110011101;
        end
        8379: begin
            cosine_reg0 <= 36'sb100000000101010000111001011001010000;
            sine_reg0   <= 36'sb111101101101010000011010001101011010;
        end
        8380: begin
            cosine_reg0 <= 36'sb100000000101010100100000100000111010;
            sine_reg0   <= 36'sb111101101100011110010001100010000001;
        end
        8381: begin
            cosine_reg0 <= 36'sb100000000101011000001000110111010100;
            sine_reg0   <= 36'sb111101101011101100001000111100010100;
        end
        8382: begin
            cosine_reg0 <= 36'sb100000000101011011110010011100011110;
            sine_reg0   <= 36'sb111101101010111010000000011100010110;
        end
        8383: begin
            cosine_reg0 <= 36'sb100000000101011111011101010000010111;
            sine_reg0   <= 36'sb111101101010000111111000000010000111;
        end
        8384: begin
            cosine_reg0 <= 36'sb100000000101100011001001010011000001;
            sine_reg0   <= 36'sb111101101001010101101111101101101010;
        end
        8385: begin
            cosine_reg0 <= 36'sb100000000101100110110110100100011010;
            sine_reg0   <= 36'sb111101101000100011100111011111000000;
        end
        8386: begin
            cosine_reg0 <= 36'sb100000000101101010100101000100100010;
            sine_reg0   <= 36'sb111101100111110001011111010110001101;
        end
        8387: begin
            cosine_reg0 <= 36'sb100000000101101110010100110011011001;
            sine_reg0   <= 36'sb111101100110111111010111010011010001;
        end
        8388: begin
            cosine_reg0 <= 36'sb100000000101110010000101110001000000;
            sine_reg0   <= 36'sb111101100110001101001111010110001110;
        end
        8389: begin
            cosine_reg0 <= 36'sb100000000101110101110111111101010110;
            sine_reg0   <= 36'sb111101100101011011000111011111000111;
        end
        8390: begin
            cosine_reg0 <= 36'sb100000000101111001101011011000011010;
            sine_reg0   <= 36'sb111101100100101000111111101101111101;
        end
        8391: begin
            cosine_reg0 <= 36'sb100000000101111101100000000010001101;
            sine_reg0   <= 36'sb111101100011110110111000000010110011;
        end
        8392: begin
            cosine_reg0 <= 36'sb100000000110000001010101111010101111;
            sine_reg0   <= 36'sb111101100011000100110000011101101010;
        end
        8393: begin
            cosine_reg0 <= 36'sb100000000110000101001101000001111111;
            sine_reg0   <= 36'sb111101100010010010101000111110100100;
        end
        8394: begin
            cosine_reg0 <= 36'sb100000000110001001000101010111111101;
            sine_reg0   <= 36'sb111101100001100000100001100101100011;
        end
        8395: begin
            cosine_reg0 <= 36'sb100000000110001100111110111100101010;
            sine_reg0   <= 36'sb111101100000101110011010010010101010;
        end
        8396: begin
            cosine_reg0 <= 36'sb100000000110010000111001110000000100;
            sine_reg0   <= 36'sb111101011111111100010011000101111001;
        end
        8397: begin
            cosine_reg0 <= 36'sb100000000110010100110101110010001100;
            sine_reg0   <= 36'sb111101011111001010001011111111010011;
        end
        8398: begin
            cosine_reg0 <= 36'sb100000000110011000110011000011000010;
            sine_reg0   <= 36'sb111101011110011000000100111110111010;
        end
        8399: begin
            cosine_reg0 <= 36'sb100000000110011100110001100010100101;
            sine_reg0   <= 36'sb111101011101100101111110000100110000;
        end
        8400: begin
            cosine_reg0 <= 36'sb100000000110100000110001010000110101;
            sine_reg0   <= 36'sb111101011100110011110111010000110111;
        end
        8401: begin
            cosine_reg0 <= 36'sb100000000110100100110010001101110011;
            sine_reg0   <= 36'sb111101011100000001110000100011010000;
        end
        8402: begin
            cosine_reg0 <= 36'sb100000000110101000110100011001011110;
            sine_reg0   <= 36'sb111101011011001111101001111011111110;
        end
        8403: begin
            cosine_reg0 <= 36'sb100000000110101100110111110011110101;
            sine_reg0   <= 36'sb111101011010011101100011011011000010;
        end
        8404: begin
            cosine_reg0 <= 36'sb100000000110110000111100011100111010;
            sine_reg0   <= 36'sb111101011001101011011101000000011111;
        end
        8405: begin
            cosine_reg0 <= 36'sb100000000110110101000010010100101010;
            sine_reg0   <= 36'sb111101011000111001010110101100010110;
        end
        8406: begin
            cosine_reg0 <= 36'sb100000000110111001001001011011001000;
            sine_reg0   <= 36'sb111101011000000111010000011110101010;
        end
        8407: begin
            cosine_reg0 <= 36'sb100000000110111101010001110000010001;
            sine_reg0   <= 36'sb111101010111010101001010010111011100;
        end
        8408: begin
            cosine_reg0 <= 36'sb100000000111000001011011010100000111;
            sine_reg0   <= 36'sb111101010110100011000100010110101110;
        end
        8409: begin
            cosine_reg0 <= 36'sb100000000111000101100110000110101000;
            sine_reg0   <= 36'sb111101010101110000111110011100100010;
        end
        8410: begin
            cosine_reg0 <= 36'sb100000000111001001110010000111110101;
            sine_reg0   <= 36'sb111101010100111110111000101000111010;
        end
        8411: begin
            cosine_reg0 <= 36'sb100000000111001101111111010111101110;
            sine_reg0   <= 36'sb111101010100001100110010111011111000;
        end
        8412: begin
            cosine_reg0 <= 36'sb100000000111010010001101110110010010;
            sine_reg0   <= 36'sb111101010011011010101101010101011110;
        end
        8413: begin
            cosine_reg0 <= 36'sb100000000111010110011101100011100001;
            sine_reg0   <= 36'sb111101010010101000100111110101101110;
        end
        8414: begin
            cosine_reg0 <= 36'sb100000000111011010101110011111011100;
            sine_reg0   <= 36'sb111101010001110110100010011100101001;
        end
        8415: begin
            cosine_reg0 <= 36'sb100000000111011111000000101010000001;
            sine_reg0   <= 36'sb111101010001000100011101001010010010;
        end
        8416: begin
            cosine_reg0 <= 36'sb100000000111100011010100000011010010;
            sine_reg0   <= 36'sb111101010000010010010111111110101011;
        end
        8417: begin
            cosine_reg0 <= 36'sb100000000111100111101000101011001100;
            sine_reg0   <= 36'sb111101001111100000010010111001110110;
        end
        8418: begin
            cosine_reg0 <= 36'sb100000000111101011111110100001110010;
            sine_reg0   <= 36'sb111101001110101110001101111011110100;
        end
        8419: begin
            cosine_reg0 <= 36'sb100000000111110000010101100111000001;
            sine_reg0   <= 36'sb111101001101111100001001000100100111;
        end
        8420: begin
            cosine_reg0 <= 36'sb100000000111110100101101111010111011;
            sine_reg0   <= 36'sb111101001101001010000100010100010010;
        end
        8421: begin
            cosine_reg0 <= 36'sb100000000111111001000111011101011111;
            sine_reg0   <= 36'sb111101001100010111111111101010110101;
        end
        8422: begin
            cosine_reg0 <= 36'sb100000000111111101100010001110101100;
            sine_reg0   <= 36'sb111101001011100101111011001000010101;
        end
        8423: begin
            cosine_reg0 <= 36'sb100000001000000001111110001110100011;
            sine_reg0   <= 36'sb111101001010110011110110101100110001;
        end
        8424: begin
            cosine_reg0 <= 36'sb100000001000000110011011011101000011;
            sine_reg0   <= 36'sb111101001010000001110010011000001100;
        end
        8425: begin
            cosine_reg0 <= 36'sb100000001000001010111001111010001101;
            sine_reg0   <= 36'sb111101001001001111101110001010101001;
        end
        8426: begin
            cosine_reg0 <= 36'sb100000001000001111011001100101111111;
            sine_reg0   <= 36'sb111101001000011101101010000100001000;
        end
        8427: begin
            cosine_reg0 <= 36'sb100000001000010011111010100000011011;
            sine_reg0   <= 36'sb111101000111101011100110000100101100;
        end
        8428: begin
            cosine_reg0 <= 36'sb100000001000011000011100101001011111;
            sine_reg0   <= 36'sb111101000110111001100010001100010111;
        end
        8429: begin
            cosine_reg0 <= 36'sb100000001000011101000000000001001100;
            sine_reg0   <= 36'sb111101000110000111011110011011001011;
        end
        8430: begin
            cosine_reg0 <= 36'sb100000001000100001100100100111100010;
            sine_reg0   <= 36'sb111101000101010101011010110001001001;
        end
        8431: begin
            cosine_reg0 <= 36'sb100000001000100110001010011100011111;
            sine_reg0   <= 36'sb111101000100100011010111001110010100;
        end
        8432: begin
            cosine_reg0 <= 36'sb100000001000101010110001100000000101;
            sine_reg0   <= 36'sb111101000011110001010011110010101101;
        end
        8433: begin
            cosine_reg0 <= 36'sb100000001000101111011001110010010010;
            sine_reg0   <= 36'sb111101000010111111010000011110010111;
        end
        8434: begin
            cosine_reg0 <= 36'sb100000001000110100000011010011000111;
            sine_reg0   <= 36'sb111101000010001101001101010001010011;
        end
        8435: begin
            cosine_reg0 <= 36'sb100000001000111000101110000010100011;
            sine_reg0   <= 36'sb111101000001011011001010001011100100;
        end
        8436: begin
            cosine_reg0 <= 36'sb100000001000111101011010000000100111;
            sine_reg0   <= 36'sb111101000000101001000111001101001010;
        end
        8437: begin
            cosine_reg0 <= 36'sb100000001001000010000111001101010010;
            sine_reg0   <= 36'sb111100111111110111000100010110001001;
        end
        8438: begin
            cosine_reg0 <= 36'sb100000001001000110110101101000100100;
            sine_reg0   <= 36'sb111100111111000101000001100110100010;
        end
        8439: begin
            cosine_reg0 <= 36'sb100000001001001011100101010010011101;
            sine_reg0   <= 36'sb111100111110010010111110111110010111;
        end
        8440: begin
            cosine_reg0 <= 36'sb100000001001010000010110001010111100;
            sine_reg0   <= 36'sb111100111101100000111100011101101010;
        end
        8441: begin
            cosine_reg0 <= 36'sb100000001001010101001000010010000010;
            sine_reg0   <= 36'sb111100111100101110111010000100011101;
        end
        8442: begin
            cosine_reg0 <= 36'sb100000001001011001111011100111101101;
            sine_reg0   <= 36'sb111100111011111100110111110010110001;
        end
        8443: begin
            cosine_reg0 <= 36'sb100000001001011110110000001011111111;
            sine_reg0   <= 36'sb111100111011001010110101101000101010;
        end
        8444: begin
            cosine_reg0 <= 36'sb100000001001100011100101111110110111;
            sine_reg0   <= 36'sb111100111010011000110011100110001000;
        end
        8445: begin
            cosine_reg0 <= 36'sb100000001001101000011101000000010100;
            sine_reg0   <= 36'sb111100111001100110110001101011001101;
        end
        8446: begin
            cosine_reg0 <= 36'sb100000001001101101010101010000010111;
            sine_reg0   <= 36'sb111100111000110100101111110111111100;
        end
        8447: begin
            cosine_reg0 <= 36'sb100000001001110010001110101110111111;
            sine_reg0   <= 36'sb111100111000000010101110001100010111;
        end
        8448: begin
            cosine_reg0 <= 36'sb100000001001110111001001011100001101;
            sine_reg0   <= 36'sb111100110111010000101100101000011111;
        end
        8449: begin
            cosine_reg0 <= 36'sb100000001001111100000101010111111111;
            sine_reg0   <= 36'sb111100110110011110101011001100010110;
        end
        8450: begin
            cosine_reg0 <= 36'sb100000001010000001000010100010010110;
            sine_reg0   <= 36'sb111100110101101100101001110111111110;
        end
        8451: begin
            cosine_reg0 <= 36'sb100000001010000110000000111011010001;
            sine_reg0   <= 36'sb111100110100111010101000101011011010;
        end
        8452: begin
            cosine_reg0 <= 36'sb100000001010001011000000100010110001;
            sine_reg0   <= 36'sb111100110100001000100111100110101011;
        end
        8453: begin
            cosine_reg0 <= 36'sb100000001010010000000001011000110101;
            sine_reg0   <= 36'sb111100110011010110100110101001110010;
        end
        8454: begin
            cosine_reg0 <= 36'sb100000001010010101000011011101011100;
            sine_reg0   <= 36'sb111100110010100100100101110100110011;
        end
        8455: begin
            cosine_reg0 <= 36'sb100000001010011010000110110000101000;
            sine_reg0   <= 36'sb111100110001110010100101000111101111;
        end
        8456: begin
            cosine_reg0 <= 36'sb100000001010011111001011010010010111;
            sine_reg0   <= 36'sb111100110001000000100100100010100111;
        end
        8457: begin
            cosine_reg0 <= 36'sb100000001010100100010001000010101010;
            sine_reg0   <= 36'sb111100110000001110100100000101011110;
        end
        8458: begin
            cosine_reg0 <= 36'sb100000001010101001011000000001011111;
            sine_reg0   <= 36'sb111100101111011100100011110000010110;
        end
        8459: begin
            cosine_reg0 <= 36'sb100000001010101110100000001110111000;
            sine_reg0   <= 36'sb111100101110101010100011100011010000;
        end
        8460: begin
            cosine_reg0 <= 36'sb100000001010110011101001101010110011;
            sine_reg0   <= 36'sb111100101101111000100011011110001111;
        end
        8461: begin
            cosine_reg0 <= 36'sb100000001010111000110100010101010001;
            sine_reg0   <= 36'sb111100101101000110100011100001010100;
        end
        8462: begin
            cosine_reg0 <= 36'sb100000001010111110000000001110010010;
            sine_reg0   <= 36'sb111100101100010100100011101100100010;
        end
        8463: begin
            cosine_reg0 <= 36'sb100000001011000011001101010101110100;
            sine_reg0   <= 36'sb111100101011100010100011111111111010;
        end
        8464: begin
            cosine_reg0 <= 36'sb100000001011001000011011101011111000;
            sine_reg0   <= 36'sb111100101010110000100100011011011110;
        end
        8465: begin
            cosine_reg0 <= 36'sb100000001011001101101011010000011111;
            sine_reg0   <= 36'sb111100101001111110100100111111010000;
        end
        8466: begin
            cosine_reg0 <= 36'sb100000001011010010111100000011100111;
            sine_reg0   <= 36'sb111100101001001100100101101011010010;
        end
        8467: begin
            cosine_reg0 <= 36'sb100000001011011000001110000101010000;
            sine_reg0   <= 36'sb111100101000011010100110011111100111;
        end
        8468: begin
            cosine_reg0 <= 36'sb100000001011011101100001010101011010;
            sine_reg0   <= 36'sb111100100111101000100111011100001111;
        end
        8469: begin
            cosine_reg0 <= 36'sb100000001011100010110101110100000101;
            sine_reg0   <= 36'sb111100100110110110101000100001001101;
        end
        8470: begin
            cosine_reg0 <= 36'sb100000001011101000001011100001010001;
            sine_reg0   <= 36'sb111100100110000100101001101110100011;
        end
        8471: begin
            cosine_reg0 <= 36'sb100000001011101101100010011100111110;
            sine_reg0   <= 36'sb111100100101010010101011000100010011;
        end
        8472: begin
            cosine_reg0 <= 36'sb100000001011110010111010100111001011;
            sine_reg0   <= 36'sb111100100100100000101100100010011110;
        end
        8473: begin
            cosine_reg0 <= 36'sb100000001011111000010011111111111000;
            sine_reg0   <= 36'sb111100100011101110101110001001000111;
        end
        8474: begin
            cosine_reg0 <= 36'sb100000001011111101101110100111000101;
            sine_reg0   <= 36'sb111100100010111100101111111000010000;
        end
        8475: begin
            cosine_reg0 <= 36'sb100000001100000011001010011100110010;
            sine_reg0   <= 36'sb111100100010001010110001101111111001;
        end
        8476: begin
            cosine_reg0 <= 36'sb100000001100001000100111100000111110;
            sine_reg0   <= 36'sb111100100001011000110011110000000111;
        end
        8477: begin
            cosine_reg0 <= 36'sb100000001100001110000101110011101001;
            sine_reg0   <= 36'sb111100100000100110110101111000111001;
        end
        8478: begin
            cosine_reg0 <= 36'sb100000001100010011100101010100110100;
            sine_reg0   <= 36'sb111100011111110100111000001010010011;
        end
        8479: begin
            cosine_reg0 <= 36'sb100000001100011001000110000100011101;
            sine_reg0   <= 36'sb111100011111000010111010100100010101;
        end
        8480: begin
            cosine_reg0 <= 36'sb100000001100011110101000000010100110;
            sine_reg0   <= 36'sb111100011110010000111101000111000011;
        end
        8481: begin
            cosine_reg0 <= 36'sb100000001100100100001011001111001100;
            sine_reg0   <= 36'sb111100011101011110111111110010011110;
        end
        8482: begin
            cosine_reg0 <= 36'sb100000001100101001101111101010010001;
            sine_reg0   <= 36'sb111100011100101101000010100110101000;
        end
        8483: begin
            cosine_reg0 <= 36'sb100000001100101111010101010011110100;
            sine_reg0   <= 36'sb111100011011111011000101100011100010;
        end
        8484: begin
            cosine_reg0 <= 36'sb100000001100110100111100001011110100;
            sine_reg0   <= 36'sb111100011011001001001000101001001111;
        end
        8485: begin
            cosine_reg0 <= 36'sb100000001100111010100100010010010011;
            sine_reg0   <= 36'sb111100011010010111001011110111110001;
        end
        8486: begin
            cosine_reg0 <= 36'sb100000001101000000001101100111001110;
            sine_reg0   <= 36'sb111100011001100101001111001111001010;
        end
        8487: begin
            cosine_reg0 <= 36'sb100000001101000101111000001010100111;
            sine_reg0   <= 36'sb111100011000110011010010101111011011;
        end
        8488: begin
            cosine_reg0 <= 36'sb100000001101001011100011111100011101;
            sine_reg0   <= 36'sb111100011000000001010110011000100111;
        end
        8489: begin
            cosine_reg0 <= 36'sb100000001101010001010000111100101111;
            sine_reg0   <= 36'sb111100010111001111011010001010101111;
        end
        8490: begin
            cosine_reg0 <= 36'sb100000001101010110111111001011011110;
            sine_reg0   <= 36'sb111100010110011101011110000101110101;
        end
        8491: begin
            cosine_reg0 <= 36'sb100000001101011100101110101000101001;
            sine_reg0   <= 36'sb111100010101101011100010001001111011;
        end
        8492: begin
            cosine_reg0 <= 36'sb100000001101100010011111010100010000;
            sine_reg0   <= 36'sb111100010100111001100110010111000100;
        end
        8493: begin
            cosine_reg0 <= 36'sb100000001101101000010001001110010011;
            sine_reg0   <= 36'sb111100010100000111101010101101010001;
        end
        8494: begin
            cosine_reg0 <= 36'sb100000001101101110000100010110110010;
            sine_reg0   <= 36'sb111100010011010101101111001100100011;
        end
        8495: begin
            cosine_reg0 <= 36'sb100000001101110011111000101101101100;
            sine_reg0   <= 36'sb111100010010100011110011110100111110;
        end
        8496: begin
            cosine_reg0 <= 36'sb100000001101111001101110010011000001;
            sine_reg0   <= 36'sb111100010001110001111000100110100011;
        end
        8497: begin
            cosine_reg0 <= 36'sb100000001101111111100101000110110001;
            sine_reg0   <= 36'sb111100010000111111111101100001010011;
        end
        8498: begin
            cosine_reg0 <= 36'sb100000001110000101011101001000111100;
            sine_reg0   <= 36'sb111100010000001110000010100101010001;
        end
        8499: begin
            cosine_reg0 <= 36'sb100000001110001011010110011001100010;
            sine_reg0   <= 36'sb111100001111011100000111110010011111;
        end
        8500: begin
            cosine_reg0 <= 36'sb100000001110010001010000111000100001;
            sine_reg0   <= 36'sb111100001110101010001101001000111110;
        end
        8501: begin
            cosine_reg0 <= 36'sb100000001110010111001100100101111011;
            sine_reg0   <= 36'sb111100001101111000010010101000110001;
        end
        8502: begin
            cosine_reg0 <= 36'sb100000001110011101001001100001101110;
            sine_reg0   <= 36'sb111100001101000110011000010001111001;
        end
        8503: begin
            cosine_reg0 <= 36'sb100000001110100011000111101011111011;
            sine_reg0   <= 36'sb111100001100010100011110000100011000;
        end
        8504: begin
            cosine_reg0 <= 36'sb100000001110101001000111000100100010;
            sine_reg0   <= 36'sb111100001011100010100100000000010001;
        end
        8505: begin
            cosine_reg0 <= 36'sb100000001110101111000111101011100001;
            sine_reg0   <= 36'sb111100001010110000101010000101100101;
        end
        8506: begin
            cosine_reg0 <= 36'sb100000001110110101001001100000111001;
            sine_reg0   <= 36'sb111100001001111110110000010100010110;
        end
        8507: begin
            cosine_reg0 <= 36'sb100000001110111011001100100100101010;
            sine_reg0   <= 36'sb111100001001001100110110101100100110;
        end
        8508: begin
            cosine_reg0 <= 36'sb100000001111000001010000110110110100;
            sine_reg0   <= 36'sb111100001000011010111101001110010111;
        end
        8509: begin
            cosine_reg0 <= 36'sb100000001111000111010110010111010101;
            sine_reg0   <= 36'sb111100000111101001000011111001101011;
        end
        8510: begin
            cosine_reg0 <= 36'sb100000001111001101011101000110001111;
            sine_reg0   <= 36'sb111100000110110111001010101110100011;
        end
        8511: begin
            cosine_reg0 <= 36'sb100000001111010011100101000011100000;
            sine_reg0   <= 36'sb111100000110000101010001101101000011;
        end
        8512: begin
            cosine_reg0 <= 36'sb100000001111011001101110001111001001;
            sine_reg0   <= 36'sb111100000101010011011000110101001011;
        end
        8513: begin
            cosine_reg0 <= 36'sb100000001111011111111000101001001000;
            sine_reg0   <= 36'sb111100000100100001100000000110111101;
        end
        8514: begin
            cosine_reg0 <= 36'sb100000001111100110000100010001011111;
            sine_reg0   <= 36'sb111100000011101111100111100010011101;
        end
        8515: begin
            cosine_reg0 <= 36'sb100000001111101100010001001000001101;
            sine_reg0   <= 36'sb111100000010111101101111000111101010;
        end
        8516: begin
            cosine_reg0 <= 36'sb100000001111110010011111001101010001;
            sine_reg0   <= 36'sb111100000010001011110110110110101000;
        end
        8517: begin
            cosine_reg0 <= 36'sb100000001111111000101110100000101100;
            sine_reg0   <= 36'sb111100000001011001111110101111011000;
        end
        8518: begin
            cosine_reg0 <= 36'sb100000001111111110111111000010011100;
            sine_reg0   <= 36'sb111100000000101000000110110001111100;
        end
        8519: begin
            cosine_reg0 <= 36'sb100000010000000101010000110010100010;
            sine_reg0   <= 36'sb111011111111110110001110111110010111;
        end
        8520: begin
            cosine_reg0 <= 36'sb100000010000001011100011110000111110;
            sine_reg0   <= 36'sb111011111111000100010111010100101001;
        end
        8521: begin
            cosine_reg0 <= 36'sb100000010000010001110111111101110000;
            sine_reg0   <= 36'sb111011111110010010011111110100110110;
        end
        8522: begin
            cosine_reg0 <= 36'sb100000010000011000001101011000110110;
            sine_reg0   <= 36'sb111011111101100000101000011110111110;
        end
        8523: begin
            cosine_reg0 <= 36'sb100000010000011110100100000010010001;
            sine_reg0   <= 36'sb111011111100101110110001010011000100;
        end
        8524: begin
            cosine_reg0 <= 36'sb100000010000100100111011111010000000;
            sine_reg0   <= 36'sb111011111011111100111010010001001010;
        end
        8525: begin
            cosine_reg0 <= 36'sb100000010000101011010101000000000100;
            sine_reg0   <= 36'sb111011111011001011000011011001010001;
        end
        8526: begin
            cosine_reg0 <= 36'sb100000010000110001101111010100011101;
            sine_reg0   <= 36'sb111011111010011001001100101011011100;
        end
        8527: begin
            cosine_reg0 <= 36'sb100000010000111000001010110111001000;
            sine_reg0   <= 36'sb111011111001100111010110000111101101;
        end
        8528: begin
            cosine_reg0 <= 36'sb100000010000111110100111101000001000;
            sine_reg0   <= 36'sb111011111000110101011111101110000100;
        end
        8529: begin
            cosine_reg0 <= 36'sb100000010001000101000101100111011011;
            sine_reg0   <= 36'sb111011111000000011101001011110100110;
        end
        8530: begin
            cosine_reg0 <= 36'sb100000010001001011100100110101000001;
            sine_reg0   <= 36'sb111011110111010001110011011001010010;
        end
        8531: begin
            cosine_reg0 <= 36'sb100000010001010010000101010000111010;
            sine_reg0   <= 36'sb111011110110011111111101011110001100;
        end
        8532: begin
            cosine_reg0 <= 36'sb100000010001011000100110111011000101;
            sine_reg0   <= 36'sb111011110101101110000111101101010101;
        end
        8533: begin
            cosine_reg0 <= 36'sb100000010001011111001001110011100011;
            sine_reg0   <= 36'sb111011110100111100010010000110101110;
        end
        8534: begin
            cosine_reg0 <= 36'sb100000010001100101101101111010010010;
            sine_reg0   <= 36'sb111011110100001010011100101010011011;
        end
        8535: begin
            cosine_reg0 <= 36'sb100000010001101100010011001111010100;
            sine_reg0   <= 36'sb111011110011011000100111011000011101;
        end
        8536: begin
            cosine_reg0 <= 36'sb100000010001110010111001110010100111;
            sine_reg0   <= 36'sb111011110010100110110010010000110101;
        end
        8537: begin
            cosine_reg0 <= 36'sb100000010001111001100001100100001100;
            sine_reg0   <= 36'sb111011110001110100111101010011100110;
        end
        8538: begin
            cosine_reg0 <= 36'sb100000010010000000001010100100000010;
            sine_reg0   <= 36'sb111011110001000011001000100000110010;
        end
        8539: begin
            cosine_reg0 <= 36'sb100000010010000110110100110010001000;
            sine_reg0   <= 36'sb111011110000010001010011111000011010;
        end
        8540: begin
            cosine_reg0 <= 36'sb100000010010001101100000001110011111;
            sine_reg0   <= 36'sb111011101111011111011111011010100001;
        end
        8541: begin
            cosine_reg0 <= 36'sb100000010010010100001100111001000110;
            sine_reg0   <= 36'sb111011101110101101101011000111001000;
        end
        8542: begin
            cosine_reg0 <= 36'sb100000010010011010111010110001111110;
            sine_reg0   <= 36'sb111011101101111011110110111110010001;
        end
        8543: begin
            cosine_reg0 <= 36'sb100000010010100001101001111001000101;
            sine_reg0   <= 36'sb111011101101001010000010111111111111;
        end
        8544: begin
            cosine_reg0 <= 36'sb100000010010101000011010001110011100;
            sine_reg0   <= 36'sb111011101100011000001111001100010010;
        end
        8545: begin
            cosine_reg0 <= 36'sb100000010010101111001011110010000001;
            sine_reg0   <= 36'sb111011101011100110011011100011001110;
        end
        8546: begin
            cosine_reg0 <= 36'sb100000010010110101111110100011110110;
            sine_reg0   <= 36'sb111011101010110100101000000100110100;
        end
        8547: begin
            cosine_reg0 <= 36'sb100000010010111100110010100011111010;
            sine_reg0   <= 36'sb111011101010000010110100110001000110;
        end
        8548: begin
            cosine_reg0 <= 36'sb100000010011000011100111110010001100;
            sine_reg0   <= 36'sb111011101001010001000001101000000101;
        end
        8549: begin
            cosine_reg0 <= 36'sb100000010011001010011110001110101101;
            sine_reg0   <= 36'sb111011101000011111001110101001110101;
        end
        8550: begin
            cosine_reg0 <= 36'sb100000010011010001010101111001011011;
            sine_reg0   <= 36'sb111011100111101101011011110110010110;
        end
        8551: begin
            cosine_reg0 <= 36'sb100000010011011000001110110010010111;
            sine_reg0   <= 36'sb111011100110111011101001001101101010;
        end
        8552: begin
            cosine_reg0 <= 36'sb100000010011011111001000111001100001;
            sine_reg0   <= 36'sb111011100110001001110110101111110100;
        end
        8553: begin
            cosine_reg0 <= 36'sb100000010011100110000100001110110111;
            sine_reg0   <= 36'sb111011100101011000000100011100110110;
        end
        8554: begin
            cosine_reg0 <= 36'sb100000010011101101000000110010011011;
            sine_reg0   <= 36'sb111011100100100110010010010100110001;
        end
        8555: begin
            cosine_reg0 <= 36'sb100000010011110011111110100100001011;
            sine_reg0   <= 36'sb111011100011110100100000010111100111;
        end
        8556: begin
            cosine_reg0 <= 36'sb100000010011111010111101100100000111;
            sine_reg0   <= 36'sb111011100011000010101110100101011010;
        end
        8557: begin
            cosine_reg0 <= 36'sb100000010100000001111101110010010000;
            sine_reg0   <= 36'sb111011100010010000111100111110001100;
        end
        8558: begin
            cosine_reg0 <= 36'sb100000010100001000111111001110100100;
            sine_reg0   <= 36'sb111011100001011111001011100010000000;
        end
        8559: begin
            cosine_reg0 <= 36'sb100000010100010000000001111001000100;
            sine_reg0   <= 36'sb111011100000101101011010010000110110;
        end
        8560: begin
            cosine_reg0 <= 36'sb100000010100010111000101110001101111;
            sine_reg0   <= 36'sb111011011111111011101001001010110001;
        end
        8561: begin
            cosine_reg0 <= 36'sb100000010100011110001010111000100101;
            sine_reg0   <= 36'sb111011011111001001111000001111110011;
        end
        8562: begin
            cosine_reg0 <= 36'sb100000010100100101010001001101100110;
            sine_reg0   <= 36'sb111011011110011000000111011111111110;
        end
        8563: begin
            cosine_reg0 <= 36'sb100000010100101100011000110000110010;
            sine_reg0   <= 36'sb111011011101100110010110111011010011;
        end
        8564: begin
            cosine_reg0 <= 36'sb100000010100110011100001100010000111;
            sine_reg0   <= 36'sb111011011100110100100110100001110101;
        end
        8565: begin
            cosine_reg0 <= 36'sb100000010100111010101011100001100111;
            sine_reg0   <= 36'sb111011011100000010110110010011100110;
        end
        8566: begin
            cosine_reg0 <= 36'sb100000010101000001110110101111010000;
            sine_reg0   <= 36'sb111011011011010001000110010000100110;
        end
        8567: begin
            cosine_reg0 <= 36'sb100000010101001001000011001011000010;
            sine_reg0   <= 36'sb111011011010011111010110011000111001;
        end
        8568: begin
            cosine_reg0 <= 36'sb100000010101010000010000110100111110;
            sine_reg0   <= 36'sb111011011001101101100110101100100000;
        end
        8569: begin
            cosine_reg0 <= 36'sb100000010101010111011111101101000010;
            sine_reg0   <= 36'sb111011011000111011110111001011011110;
        end
        8570: begin
            cosine_reg0 <= 36'sb100000010101011110101111110011001111;
            sine_reg0   <= 36'sb111011011000001010000111110101110011;
        end
        8571: begin
            cosine_reg0 <= 36'sb100000010101100110000001000111100100;
            sine_reg0   <= 36'sb111011010111011000011000101011100010;
        end
        8572: begin
            cosine_reg0 <= 36'sb100000010101101101010011101010000001;
            sine_reg0   <= 36'sb111011010110100110101001101100101101;
        end
        8573: begin
            cosine_reg0 <= 36'sb100000010101110100100111011010100110;
            sine_reg0   <= 36'sb111011010101110100111010111001010110;
        end
        8574: begin
            cosine_reg0 <= 36'sb100000010101111011111100011001010010;
            sine_reg0   <= 36'sb111011010101000011001100010001011111;
        end
        8575: begin
            cosine_reg0 <= 36'sb100000010110000011010010100110000101;
            sine_reg0   <= 36'sb111011010100010001011101110101001001;
        end
        8576: begin
            cosine_reg0 <= 36'sb100000010110001010101010000000111111;
            sine_reg0   <= 36'sb111011010011011111101111100100010111;
        end
        8577: begin
            cosine_reg0 <= 36'sb100000010110010010000010101001111111;
            sine_reg0   <= 36'sb111011010010101110000001011111001011;
        end
        8578: begin
            cosine_reg0 <= 36'sb100000010110011001011100100001000110;
            sine_reg0   <= 36'sb111011010001111100010011100101100101;
        end
        8579: begin
            cosine_reg0 <= 36'sb100000010110100000110111100110010011;
            sine_reg0   <= 36'sb111011010001001010100101110111101001;
        end
        8580: begin
            cosine_reg0 <= 36'sb100000010110101000010011111001100101;
            sine_reg0   <= 36'sb111011010000011000111000010101011000;
        end
        8581: begin
            cosine_reg0 <= 36'sb100000010110101111110001011010111101;
            sine_reg0   <= 36'sb111011001111100111001010111110110101;
        end
        8582: begin
            cosine_reg0 <= 36'sb100000010110110111010000001010011010;
            sine_reg0   <= 36'sb111011001110110101011101110100000000;
        end
        8583: begin
            cosine_reg0 <= 36'sb100000010110111110110000000111111100;
            sine_reg0   <= 36'sb111011001110000011110000110100111101;
        end
        8584: begin
            cosine_reg0 <= 36'sb100000010111000110010001010011100010;
            sine_reg0   <= 36'sb111011001101010010000100000001101100;
        end
        8585: begin
            cosine_reg0 <= 36'sb100000010111001101110011101101001101;
            sine_reg0   <= 36'sb111011001100100000010111011010010000;
        end
        8586: begin
            cosine_reg0 <= 36'sb100000010111010101010111010100111100;
            sine_reg0   <= 36'sb111011001011101110101010111110101011;
        end
        8587: begin
            cosine_reg0 <= 36'sb100000010111011100111100001010101110;
            sine_reg0   <= 36'sb111011001010111100111110101110111110;
        end
        8588: begin
            cosine_reg0 <= 36'sb100000010111100100100010001110100011;
            sine_reg0   <= 36'sb111011001010001011010010101011001100;
        end
        8589: begin
            cosine_reg0 <= 36'sb100000010111101100001001100000011100;
            sine_reg0   <= 36'sb111011001001011001100110110011010110;
        end
        8590: begin
            cosine_reg0 <= 36'sb100000010111110011110010000000010111;
            sine_reg0   <= 36'sb111011001000100111111011000111011111;
        end
        8591: begin
            cosine_reg0 <= 36'sb100000010111111011011011101110010101;
            sine_reg0   <= 36'sb111011000111110110001111100111101000;
        end
        8592: begin
            cosine_reg0 <= 36'sb100000011000000011000110101010010110;
            sine_reg0   <= 36'sb111011000111000100100100010011110011;
        end
        8593: begin
            cosine_reg0 <= 36'sb100000011000001010110010110100011000;
            sine_reg0   <= 36'sb111011000110010010111001001100000011;
        end
        8594: begin
            cosine_reg0 <= 36'sb100000011000010010100000001100011011;
            sine_reg0   <= 36'sb111011000101100001001110010000011000;
        end
        8595: begin
            cosine_reg0 <= 36'sb100000011000011010001110110010100000;
            sine_reg0   <= 36'sb111011000100101111100011100000110101;
        end
        8596: begin
            cosine_reg0 <= 36'sb100000011000100001111110100110100110;
            sine_reg0   <= 36'sb111011000011111101111000111101011101;
        end
        8597: begin
            cosine_reg0 <= 36'sb100000011000101001101111101000101101;
            sine_reg0   <= 36'sb111011000011001100001110100110010000;
        end
        8598: begin
            cosine_reg0 <= 36'sb100000011000110001100001111000110100;
            sine_reg0   <= 36'sb111011000010011010100100011011010000;
        end
        8599: begin
            cosine_reg0 <= 36'sb100000011000111001010101010110111011;
            sine_reg0   <= 36'sb111011000001101000111010011100100001;
        end
        8600: begin
            cosine_reg0 <= 36'sb100000011001000001001010000011000010;
            sine_reg0   <= 36'sb111011000000110111010000101010000010;
        end
        8601: begin
            cosine_reg0 <= 36'sb100000011001001000111111111101001001;
            sine_reg0   <= 36'sb111011000000000101100111000011111000;
        end
        8602: begin
            cosine_reg0 <= 36'sb100000011001010000110111000101001110;
            sine_reg0   <= 36'sb111010111111010011111101101010000010;
        end
        8603: begin
            cosine_reg0 <= 36'sb100000011001011000101111011011010011;
            sine_reg0   <= 36'sb111010111110100010010100011100100100;
        end
        8604: begin
            cosine_reg0 <= 36'sb100000011001100000101000111111010110;
            sine_reg0   <= 36'sb111010111101110000101011011011011111;
        end
        8605: begin
            cosine_reg0 <= 36'sb100000011001101000100011110001011000;
            sine_reg0   <= 36'sb111010111100111111000010100110110101;
        end
        8606: begin
            cosine_reg0 <= 36'sb100000011001110000011111110001010111;
            sine_reg0   <= 36'sb111010111100001101011001111110101001;
        end
        8607: begin
            cosine_reg0 <= 36'sb100000011001111000011100111111010100;
            sine_reg0   <= 36'sb111010111011011011110001100010111011;
        end
        8608: begin
            cosine_reg0 <= 36'sb100000011010000000011011011011001111;
            sine_reg0   <= 36'sb111010111010101010001001010011101110;
        end
        8609: begin
            cosine_reg0 <= 36'sb100000011010001000011011000101000110;
            sine_reg0   <= 36'sb111010111001111000100001010001000011;
        end
        8610: begin
            cosine_reg0 <= 36'sb100000011010010000011011111100111011;
            sine_reg0   <= 36'sb111010111001000110111001011010111110;
        end
        8611: begin
            cosine_reg0 <= 36'sb100000011010011000011110000010101100;
            sine_reg0   <= 36'sb111010111000010101010001110001011110;
        end
        8612: begin
            cosine_reg0 <= 36'sb100000011010100000100001010110011001;
            sine_reg0   <= 36'sb111010110111100011101010010100101000;
        end
        8613: begin
            cosine_reg0 <= 36'sb100000011010101000100101111000000001;
            sine_reg0   <= 36'sb111010110110110010000011000100011100;
        end
        8614: begin
            cosine_reg0 <= 36'sb100000011010110000101011100111100110;
            sine_reg0   <= 36'sb111010110110000000011100000000111100;
        end
        8615: begin
            cosine_reg0 <= 36'sb100000011010111000110010100101000101;
            sine_reg0   <= 36'sb111010110101001110110101001010001010;
        end
        8616: begin
            cosine_reg0 <= 36'sb100000011011000000111010110000100000;
            sine_reg0   <= 36'sb111010110100011101001110100000001001;
        end
        8617: begin
            cosine_reg0 <= 36'sb100000011011001001000100001001110101;
            sine_reg0   <= 36'sb111010110011101011101000000010111001;
        end
        8618: begin
            cosine_reg0 <= 36'sb100000011011010001001110110001000100;
            sine_reg0   <= 36'sb111010110010111010000001110010011110;
        end
        8619: begin
            cosine_reg0 <= 36'sb100000011011011001011010100110001101;
            sine_reg0   <= 36'sb111010110010001000011011101110111000;
        end
        8620: begin
            cosine_reg0 <= 36'sb100000011011100001100111101001010000;
            sine_reg0   <= 36'sb111010110001010110110101111000001010;
        end
        8621: begin
            cosine_reg0 <= 36'sb100000011011101001110101111010001100;
            sine_reg0   <= 36'sb111010110000100101010000001110010110;
        end
        8622: begin
            cosine_reg0 <= 36'sb100000011011110010000101011001000001;
            sine_reg0   <= 36'sb111010101111110011101010110001011101;
        end
        8623: begin
            cosine_reg0 <= 36'sb100000011011111010010110000101101111;
            sine_reg0   <= 36'sb111010101111000010000101100001100010;
        end
        8624: begin
            cosine_reg0 <= 36'sb100000011100000010101000000000010101;
            sine_reg0   <= 36'sb111010101110010000100000011110100111;
        end
        8625: begin
            cosine_reg0 <= 36'sb100000011100001010111011001000110100;
            sine_reg0   <= 36'sb111010101101011110111011101000101100;
        end
        8626: begin
            cosine_reg0 <= 36'sb100000011100010011001111011111001010;
            sine_reg0   <= 36'sb111010101100101101010110111111110101;
        end
        8627: begin
            cosine_reg0 <= 36'sb100000011100011011100101000011010111;
            sine_reg0   <= 36'sb111010101011111011110010100100000100;
        end
        8628: begin
            cosine_reg0 <= 36'sb100000011100100011111011110101011100;
            sine_reg0   <= 36'sb111010101011001010001110010101011001;
        end
        8629: begin
            cosine_reg0 <= 36'sb100000011100101100010011110101010111;
            sine_reg0   <= 36'sb111010101010011000101010010011110111;
        end
        8630: begin
            cosine_reg0 <= 36'sb100000011100110100101101000011001001;
            sine_reg0   <= 36'sb111010101001100111000110011111100000;
        end
        8631: begin
            cosine_reg0 <= 36'sb100000011100111101000111011110110001;
            sine_reg0   <= 36'sb111010101000110101100010111000010110;
        end
        8632: begin
            cosine_reg0 <= 36'sb100000011101000101100011001000001110;
            sine_reg0   <= 36'sb111010101000000011111111011110011011;
        end
        8633: begin
            cosine_reg0 <= 36'sb100000011101001101111111111111100001;
            sine_reg0   <= 36'sb111010100111010010011100010001110000;
        end
        8634: begin
            cosine_reg0 <= 36'sb100000011101010110011110000100101010;
            sine_reg0   <= 36'sb111010100110100000111001010010011000;
        end
        8635: begin
            cosine_reg0 <= 36'sb100000011101011110111101010111100111;
            sine_reg0   <= 36'sb111010100101101111010110100000010100;
        end
        8636: begin
            cosine_reg0 <= 36'sb100000011101100111011101111000011000;
            sine_reg0   <= 36'sb111010100100111101110011111011100111;
        end
        8637: begin
            cosine_reg0 <= 36'sb100000011101101111111111100110111110;
            sine_reg0   <= 36'sb111010100100001100010001100100010010;
        end
        8638: begin
            cosine_reg0 <= 36'sb100000011101111000100010100011010111;
            sine_reg0   <= 36'sb111010100011011010101111011010010111;
        end
        8639: begin
            cosine_reg0 <= 36'sb100000011110000001000110101101100100;
            sine_reg0   <= 36'sb111010100010101001001101011101111000;
        end
        8640: begin
            cosine_reg0 <= 36'sb100000011110001001101100000101100101;
            sine_reg0   <= 36'sb111010100001110111101011101110110111;
        end
        8641: begin
            cosine_reg0 <= 36'sb100000011110010010010010101011011000;
            sine_reg0   <= 36'sb111010100001000110001010001101010111;
        end
        8642: begin
            cosine_reg0 <= 36'sb100000011110011010111010011110111101;
            sine_reg0   <= 36'sb111010100000010100101000111001011000;
        end
        8643: begin
            cosine_reg0 <= 36'sb100000011110100011100011100000010101;
            sine_reg0   <= 36'sb111010011111100011000111110010111100;
        end
        8644: begin
            cosine_reg0 <= 36'sb100000011110101100001101101111011111;
            sine_reg0   <= 36'sb111010011110110001100110111010000111;
        end
        8645: begin
            cosine_reg0 <= 36'sb100000011110110100111001001100011010;
            sine_reg0   <= 36'sb111010011110000000000110001110111000;
        end
        8646: begin
            cosine_reg0 <= 36'sb100000011110111101100101110111000110;
            sine_reg0   <= 36'sb111010011101001110100101110001010100;
        end
        8647: begin
            cosine_reg0 <= 36'sb100000011111000110010011101111100011;
            sine_reg0   <= 36'sb111010011100011101000101100001011010;
        end
        8648: begin
            cosine_reg0 <= 36'sb100000011111001111000010110101110001;
            sine_reg0   <= 36'sb111010011011101011100101011111001110;
        end
        8649: begin
            cosine_reg0 <= 36'sb100000011111010111110011001001101111;
            sine_reg0   <= 36'sb111010011010111010000101101010110001;
        end
        8650: begin
            cosine_reg0 <= 36'sb100000011111100000100100101011011100;
            sine_reg0   <= 36'sb111010011010001000100110000100000110;
        end
        8651: begin
            cosine_reg0 <= 36'sb100000011111101001010111011010111001;
            sine_reg0   <= 36'sb111010011001010111000110101011001101;
        end
        8652: begin
            cosine_reg0 <= 36'sb100000011111110010001011011000000110;
            sine_reg0   <= 36'sb111010011000100101100111100000001001;
        end
        8653: begin
            cosine_reg0 <= 36'sb100000011111111011000000100011000001;
            sine_reg0   <= 36'sb111010010111110100001000100010111100;
        end
        8654: begin
            cosine_reg0 <= 36'sb100000100000000011110110111011101010;
            sine_reg0   <= 36'sb111010010111000010101001110011101000;
        end
        8655: begin
            cosine_reg0 <= 36'sb100000100000001100101110100010000010;
            sine_reg0   <= 36'sb111010010110010001001011010010001110;
        end
        8656: begin
            cosine_reg0 <= 36'sb100000100000010101100111010110000111;
            sine_reg0   <= 36'sb111010010101011111101100111110110001;
        end
        8657: begin
            cosine_reg0 <= 36'sb100000100000011110100001010111111010;
            sine_reg0   <= 36'sb111010010100101110001110111001010010;
        end
        8658: begin
            cosine_reg0 <= 36'sb100000100000100111011100100111011010;
            sine_reg0   <= 36'sb111010010011111100110001000001110100;
        end
        8659: begin
            cosine_reg0 <= 36'sb100000100000110000011001000100100111;
            sine_reg0   <= 36'sb111010010011001011010011011000011000;
        end
        8660: begin
            cosine_reg0 <= 36'sb100000100000111001010110101111100000;
            sine_reg0   <= 36'sb111010010010011001110101111101000000;
        end
        8661: begin
            cosine_reg0 <= 36'sb100000100001000010010101101000000110;
            sine_reg0   <= 36'sb111010010001101000011000101111101110;
        end
        8662: begin
            cosine_reg0 <= 36'sb100000100001001011010101101110010111;
            sine_reg0   <= 36'sb111010010000110110111011110000100100;
        end
        8663: begin
            cosine_reg0 <= 36'sb100000100001010100010111000010010011;
            sine_reg0   <= 36'sb111010010000000101011110111111100100;
        end
        8664: begin
            cosine_reg0 <= 36'sb100000100001011101011001100011111010;
            sine_reg0   <= 36'sb111010001111010100000010011100110000;
        end
        8665: begin
            cosine_reg0 <= 36'sb100000100001100110011101010011001101;
            sine_reg0   <= 36'sb111010001110100010100110001000001001;
        end
        8666: begin
            cosine_reg0 <= 36'sb100000100001101111100010010000001001;
            sine_reg0   <= 36'sb111010001101110001001010000001110010;
        end
        8667: begin
            cosine_reg0 <= 36'sb100000100001111000101000011010101111;
            sine_reg0   <= 36'sb111010001100111111101110001001101101;
        end
        8668: begin
            cosine_reg0 <= 36'sb100000100010000001101111110010111111;
            sine_reg0   <= 36'sb111010001100001110010010011111111011;
        end
        8669: begin
            cosine_reg0 <= 36'sb100000100010001010111000011000111001;
            sine_reg0   <= 36'sb111010001011011100110111000100011110;
        end
        8670: begin
            cosine_reg0 <= 36'sb100000100010010100000010001100011011;
            sine_reg0   <= 36'sb111010001010101011011011110111011001;
        end
        8671: begin
            cosine_reg0 <= 36'sb100000100010011101001101001101100110;
            sine_reg0   <= 36'sb111010001001111010000000111000101100;
        end
        8672: begin
            cosine_reg0 <= 36'sb100000100010100110011001011100011001;
            sine_reg0   <= 36'sb111010001001001000100110001000011011;
        end
        8673: begin
            cosine_reg0 <= 36'sb100000100010101111100110111000110100;
            sine_reg0   <= 36'sb111010001000010111001011100110100111;
        end
        8674: begin
            cosine_reg0 <= 36'sb100000100010111000110101100010110110;
            sine_reg0   <= 36'sb111010000111100101110001010011010001;
        end
        8675: begin
            cosine_reg0 <= 36'sb100000100011000010000101011010100000;
            sine_reg0   <= 36'sb111010000110110100010111001110011101;
        end
        8676: begin
            cosine_reg0 <= 36'sb100000100011001011010110011111110000;
            sine_reg0   <= 36'sb111010000110000010111101011000001011;
        end
        8677: begin
            cosine_reg0 <= 36'sb100000100011010100101000110010100111;
            sine_reg0   <= 36'sb111010000101010001100011110000011101;
        end
        8678: begin
            cosine_reg0 <= 36'sb100000100011011101111100010011000100;
            sine_reg0   <= 36'sb111010000100100000001010010111010110;
        end
        8679: begin
            cosine_reg0 <= 36'sb100000100011100111010001000001000110;
            sine_reg0   <= 36'sb111010000011101110110001001100110111;
        end
        8680: begin
            cosine_reg0 <= 36'sb100000100011110000100110111100101110;
            sine_reg0   <= 36'sb111010000010111101011000010001000011;
        end
        8681: begin
            cosine_reg0 <= 36'sb100000100011111001111110000101111011;
            sine_reg0   <= 36'sb111010000010001011111111100011111011;
        end
        8682: begin
            cosine_reg0 <= 36'sb100000100100000011010110011100101101;
            sine_reg0   <= 36'sb111010000001011010100111000101100001;
        end
        8683: begin
            cosine_reg0 <= 36'sb100000100100001100110000000001000011;
            sine_reg0   <= 36'sb111010000000101001001110110101110111;
        end
        8684: begin
            cosine_reg0 <= 36'sb100000100100010110001010110010111100;
            sine_reg0   <= 36'sb111001111111110111110110110100111110;
        end
        8685: begin
            cosine_reg0 <= 36'sb100000100100011111100110110010011010;
            sine_reg0   <= 36'sb111001111111000110011111000010111010;
        end
        8686: begin
            cosine_reg0 <= 36'sb100000100100101001000011111111011010;
            sine_reg0   <= 36'sb111001111110010101000111011111101011;
        end
        8687: begin
            cosine_reg0 <= 36'sb100000100100110010100010011001111110;
            sine_reg0   <= 36'sb111001111101100011110000001011010100;
        end
        8688: begin
            cosine_reg0 <= 36'sb100000100100111100000010000010000100;
            sine_reg0   <= 36'sb111001111100110010011001000101110110;
        end
        8689: begin
            cosine_reg0 <= 36'sb100000100101000101100010110111101011;
            sine_reg0   <= 36'sb111001111100000001000010001111010100;
        end
        8690: begin
            cosine_reg0 <= 36'sb100000100101001111000100111010110101;
            sine_reg0   <= 36'sb111001111011001111101011100111101111;
        end
        8691: begin
            cosine_reg0 <= 36'sb100000100101011000101000001011100000;
            sine_reg0   <= 36'sb111001111010011110010101001111001010;
        end
        8692: begin
            cosine_reg0 <= 36'sb100000100101100010001100101001101100;
            sine_reg0   <= 36'sb111001111001101100111111000101100101;
        end
        8693: begin
            cosine_reg0 <= 36'sb100000100101101011110010010101011001;
            sine_reg0   <= 36'sb111001111000111011101001001011000011;
        end
        8694: begin
            cosine_reg0 <= 36'sb100000100101110101011001001110100110;
            sine_reg0   <= 36'sb111001111000001010010011011111100111;
        end
        8695: begin
            cosine_reg0 <= 36'sb100000100101111111000001010101010011;
            sine_reg0   <= 36'sb111001110111011000111110000011010001;
        end
        8696: begin
            cosine_reg0 <= 36'sb100000100110001000101010101001011111;
            sine_reg0   <= 36'sb111001110110100111101000110110000100;
        end
        8697: begin
            cosine_reg0 <= 36'sb100000100110010010010101001011001010;
            sine_reg0   <= 36'sb111001110101110110010011111000000001;
        end
        8698: begin
            cosine_reg0 <= 36'sb100000100110011100000000111010010101;
            sine_reg0   <= 36'sb111001110101000100111111001001001100;
        end
        8699: begin
            cosine_reg0 <= 36'sb100000100110100101101101110110111101;
            sine_reg0   <= 36'sb111001110100010011101010101001100100;
        end
        8700: begin
            cosine_reg0 <= 36'sb100000100110101111011100000001000100;
            sine_reg0   <= 36'sb111001110011100010010110011001001101;
        end
        8701: begin
            cosine_reg0 <= 36'sb100000100110111001001011011000101000;
            sine_reg0   <= 36'sb111001110010110001000010011000001000;
        end
        8702: begin
            cosine_reg0 <= 36'sb100000100111000010111011111101101010;
            sine_reg0   <= 36'sb111001110001111111101110100110010111;
        end
        8703: begin
            cosine_reg0 <= 36'sb100000100111001100101101110000001000;
            sine_reg0   <= 36'sb111001110001001110011011000011111100;
        end
        8704: begin
            cosine_reg0 <= 36'sb100000100111010110100000110000000011;
            sine_reg0   <= 36'sb111001110000011101000111110000111010;
        end
        8705: begin
            cosine_reg0 <= 36'sb100000100111100000010100111101011010;
            sine_reg0   <= 36'sb111001101111101011110100101101010001;
        end
        8706: begin
            cosine_reg0 <= 36'sb100000100111101010001010011000001101;
            sine_reg0   <= 36'sb111001101110111010100001111001000011;
        end
        8707: begin
            cosine_reg0 <= 36'sb100000100111110100000001000000011011;
            sine_reg0   <= 36'sb111001101110001001001111010100010100;
        end
        8708: begin
            cosine_reg0 <= 36'sb100000100111111101111000110110000101;
            sine_reg0   <= 36'sb111001101101010111111100111111000100;
        end
        8709: begin
            cosine_reg0 <= 36'sb100000101000000111110001111001001001;
            sine_reg0   <= 36'sb111001101100100110101010111001010101;
        end
        8710: begin
            cosine_reg0 <= 36'sb100000101000010001101100001001100111;
            sine_reg0   <= 36'sb111001101011110101011001000011001010;
        end
        8711: begin
            cosine_reg0 <= 36'sb100000101000011011100111100111011111;
            sine_reg0   <= 36'sb111001101011000100000111011100100100;
        end
        8712: begin
            cosine_reg0 <= 36'sb100000101000100101100100010010110000;
            sine_reg0   <= 36'sb111001101010010010110110000101100101;
        end
        8713: begin
            cosine_reg0 <= 36'sb100000101000101111100010001011011011;
            sine_reg0   <= 36'sb111001101001100001100100111110001111;
        end
        8714: begin
            cosine_reg0 <= 36'sb100000101000111001100001010001011110;
            sine_reg0   <= 36'sb111001101000110000010100000110100100;
        end
        8715: begin
            cosine_reg0 <= 36'sb100000101001000011100001100100111010;
            sine_reg0   <= 36'sb111001100111111111000011011110100110;
        end
        8716: begin
            cosine_reg0 <= 36'sb100000101001001101100011000101101101;
            sine_reg0   <= 36'sb111001100111001101110011000110010111;
        end
        8717: begin
            cosine_reg0 <= 36'sb100000101001010111100101110011111000;
            sine_reg0   <= 36'sb111001100110011100100010111101111000;
        end
        8718: begin
            cosine_reg0 <= 36'sb100000101001100001101001101111011010;
            sine_reg0   <= 36'sb111001100101101011010011000101001100;
        end
        8719: begin
            cosine_reg0 <= 36'sb100000101001101011101110111000010011;
            sine_reg0   <= 36'sb111001100100111010000011011100010100;
        end
        8720: begin
            cosine_reg0 <= 36'sb100000101001110101110101001110100011;
            sine_reg0   <= 36'sb111001100100001000110100000011010010;
        end
        8721: begin
            cosine_reg0 <= 36'sb100000101001111111111100110010001000;
            sine_reg0   <= 36'sb111001100011010111100100111010001001;
        end
        8722: begin
            cosine_reg0 <= 36'sb100000101010001010000101100011000011;
            sine_reg0   <= 36'sb111001100010100110010110000000111010;
        end
        8723: begin
            cosine_reg0 <= 36'sb100000101010010100001111100001010011;
            sine_reg0   <= 36'sb111001100001110101000111010111100111;
        end
        8724: begin
            cosine_reg0 <= 36'sb100000101010011110011010101100111001;
            sine_reg0   <= 36'sb111001100001000011111000111110010010;
        end
        8725: begin
            cosine_reg0 <= 36'sb100000101010101000100111000101110010;
            sine_reg0   <= 36'sb111001100000010010101010110100111101;
        end
        8726: begin
            cosine_reg0 <= 36'sb100000101010110010110100101100000000;
            sine_reg0   <= 36'sb111001011111100001011100111011101001;
        end
        8727: begin
            cosine_reg0 <= 36'sb100000101010111101000011011111100001;
            sine_reg0   <= 36'sb111001011110110000001111010010011001;
        end
        8728: begin
            cosine_reg0 <= 36'sb100000101011000111010011100000010101;
            sine_reg0   <= 36'sb111001011101111111000001111001001111;
        end
        8729: begin
            cosine_reg0 <= 36'sb100000101011010001100100101110011100;
            sine_reg0   <= 36'sb111001011101001101110100110000001100;
        end
        8730: begin
            cosine_reg0 <= 36'sb100000101011011011110111001001110110;
            sine_reg0   <= 36'sb111001011100011100100111110111010010;
        end
        8731: begin
            cosine_reg0 <= 36'sb100000101011100110001010110010100010;
            sine_reg0   <= 36'sb111001011011101011011011001110100011;
        end
        8732: begin
            cosine_reg0 <= 36'sb100000101011110000011111101000100000;
            sine_reg0   <= 36'sb111001011010111010001110110110000010;
        end
        8733: begin
            cosine_reg0 <= 36'sb100000101011111010110101101011101110;
            sine_reg0   <= 36'sb111001011010001001000010101101110000;
        end
        8734: begin
            cosine_reg0 <= 36'sb100000101100000101001100111100001110;
            sine_reg0   <= 36'sb111001011001010111110110110101101110;
        end
        8735: begin
            cosine_reg0 <= 36'sb100000101100001111100101011001111110;
            sine_reg0   <= 36'sb111001011000100110101011001101111111;
        end
        8736: begin
            cosine_reg0 <= 36'sb100000101100011001111111000100111110;
            sine_reg0   <= 36'sb111001010111110101011111110110100101;
        end
        8737: begin
            cosine_reg0 <= 36'sb100000101100100100011001111101001110;
            sine_reg0   <= 36'sb111001010111000100010100101111100010;
        end
        8738: begin
            cosine_reg0 <= 36'sb100000101100101110110110000010101101;
            sine_reg0   <= 36'sb111001010110010011001001111000110111;
        end
        8739: begin
            cosine_reg0 <= 36'sb100000101100111001010011010101011011;
            sine_reg0   <= 36'sb111001010101100001111111010010100110;
        end
        8740: begin
            cosine_reg0 <= 36'sb100000101101000011110001110101011000;
            sine_reg0   <= 36'sb111001010100110000110100111100110010;
        end
        8741: begin
            cosine_reg0 <= 36'sb100000101101001110010001100010100010;
            sine_reg0   <= 36'sb111001010011111111101010110111011100;
        end
        8742: begin
            cosine_reg0 <= 36'sb100000101101011000110010011100111010;
            sine_reg0   <= 36'sb111001010011001110100001000010100101;
        end
        8743: begin
            cosine_reg0 <= 36'sb100000101101100011010100100100100000;
            sine_reg0   <= 36'sb111001010010011101010111011110010001;
        end
        8744: begin
            cosine_reg0 <= 36'sb100000101101101101110111111001010010;
            sine_reg0   <= 36'sb111001010001101100001110001010100001;
        end
        8745: begin
            cosine_reg0 <= 36'sb100000101101111000011100011011010000;
            sine_reg0   <= 36'sb111001010000111011000101000111010110;
        end
        8746: begin
            cosine_reg0 <= 36'sb100000101110000011000010001010011011;
            sine_reg0   <= 36'sb111001010000001001111100010100110011;
        end
        8747: begin
            cosine_reg0 <= 36'sb100000101110001101101001000110110010;
            sine_reg0   <= 36'sb111001001111011000110011110010111010;
        end
        8748: begin
            cosine_reg0 <= 36'sb100000101110011000010001010000010011;
            sine_reg0   <= 36'sb111001001110100111101011100001101100;
        end
        8749: begin
            cosine_reg0 <= 36'sb100000101110100010111010100110111111;
            sine_reg0   <= 36'sb111001001101110110100011100001001011;
        end
        8750: begin
            cosine_reg0 <= 36'sb100000101110101101100101001010110110;
            sine_reg0   <= 36'sb111001001101000101011011110001011010;
        end
        8751: begin
            cosine_reg0 <= 36'sb100000101110111000010000111011110111;
            sine_reg0   <= 36'sb111001001100010100010100010010011010;
        end
        8752: begin
            cosine_reg0 <= 36'sb100000101111000010111101111010000001;
            sine_reg0   <= 36'sb111001001011100011001101000100001100;
        end
        8753: begin
            cosine_reg0 <= 36'sb100000101111001101101100000101010101;
            sine_reg0   <= 36'sb111001001010110010000110000110110100;
        end
        8754: begin
            cosine_reg0 <= 36'sb100000101111011000011011011101110001;
            sine_reg0   <= 36'sb111001001010000000111111011010010010;
        end
        8755: begin
            cosine_reg0 <= 36'sb100000101111100011001100000011010101;
            sine_reg0   <= 36'sb111001001001001111111000111110101001;
        end
        8756: begin
            cosine_reg0 <= 36'sb100000101111101101111101110110000010;
            sine_reg0   <= 36'sb111001001000011110110010110011111011;
        end
        8757: begin
            cosine_reg0 <= 36'sb100000101111111000110000110101110101;
            sine_reg0   <= 36'sb111001000111101101101100111010001001;
        end
        8758: begin
            cosine_reg0 <= 36'sb100000110000000011100101000010110000;
            sine_reg0   <= 36'sb111001000110111100100111010001010110;
        end
        8759: begin
            cosine_reg0 <= 36'sb100000110000001110011010011100110010;
            sine_reg0   <= 36'sb111001000110001011100001111001100010;
        end
        8760: begin
            cosine_reg0 <= 36'sb100000110000011001010001000011111010;
            sine_reg0   <= 36'sb111001000101011010011100110010110001;
        end
        8761: begin
            cosine_reg0 <= 36'sb100000110000100100001000111000001000;
            sine_reg0   <= 36'sb111001000100101001010111111101000100;
        end
        8762: begin
            cosine_reg0 <= 36'sb100000110000101111000001111001011011;
            sine_reg0   <= 36'sb111001000011111000010011011000011101;
        end
        8763: begin
            cosine_reg0 <= 36'sb100000110000111001111100000111110011;
            sine_reg0   <= 36'sb111001000011000111001111000100111110;
        end
        8764: begin
            cosine_reg0 <= 36'sb100000110001000100110111100011010000;
            sine_reg0   <= 36'sb111001000010010110001011000010101000;
        end
        8765: begin
            cosine_reg0 <= 36'sb100000110001001111110100001011110001;
            sine_reg0   <= 36'sb111001000001100101000111010001011110;
        end
        8766: begin
            cosine_reg0 <= 36'sb100000110001011010110010000001010101;
            sine_reg0   <= 36'sb111001000000110100000011110001100001;
        end
        8767: begin
            cosine_reg0 <= 36'sb100000110001100101110001000011111101;
            sine_reg0   <= 36'sb111001000000000011000000100010110100;
        end
        8768: begin
            cosine_reg0 <= 36'sb100000110001110000110001010011101000;
            sine_reg0   <= 36'sb111000111111010001111101100101011000;
        end
        8769: begin
            cosine_reg0 <= 36'sb100000110001111011110010110000010101;
            sine_reg0   <= 36'sb111000111110100000111010111001010000;
        end
        8770: begin
            cosine_reg0 <= 36'sb100000110010000110110101011010000100;
            sine_reg0   <= 36'sb111000111101101111111000011110011100;
        end
        8771: begin
            cosine_reg0 <= 36'sb100000110010010001111001010000110101;
            sine_reg0   <= 36'sb111000111100111110110110010100111111;
        end
        8772: begin
            cosine_reg0 <= 36'sb100000110010011100111110010100100111;
            sine_reg0   <= 36'sb111000111100001101110100011100111011;
        end
        8773: begin
            cosine_reg0 <= 36'sb100000110010101000000100100101011010;
            sine_reg0   <= 36'sb111000111011011100110010110110010010;
        end
        8774: begin
            cosine_reg0 <= 36'sb100000110010110011001100000011001101;
            sine_reg0   <= 36'sb111000111010101011110001100001000110;
        end
        8775: begin
            cosine_reg0 <= 36'sb100000110010111110010100101110000000;
            sine_reg0   <= 36'sb111000111001111010110000011101011000;
        end
        8776: begin
            cosine_reg0 <= 36'sb100000110011001001011110100101110010;
            sine_reg0   <= 36'sb111000111001001001101111101011001010;
        end
        8777: begin
            cosine_reg0 <= 36'sb100000110011010100101001101010100100;
            sine_reg0   <= 36'sb111000111000011000101111001010011111;
        end
        8778: begin
            cosine_reg0 <= 36'sb100000110011011111110101111100010100;
            sine_reg0   <= 36'sb111000110111100111101110111011011000;
        end
        8779: begin
            cosine_reg0 <= 36'sb100000110011101011000011011011000010;
            sine_reg0   <= 36'sb111000110110110110101110111101110111;
        end
        8780: begin
            cosine_reg0 <= 36'sb100000110011110110010010000110101110;
            sine_reg0   <= 36'sb111000110110000101101111010001111110;
        end
        8781: begin
            cosine_reg0 <= 36'sb100000110100000001100001111111010111;
            sine_reg0   <= 36'sb111000110101010100101111110111101111;
        end
        8782: begin
            cosine_reg0 <= 36'sb100000110100001100110011000100111110;
            sine_reg0   <= 36'sb111000110100100011110000101111001011;
        end
        8783: begin
            cosine_reg0 <= 36'sb100000110100011000000101010111100000;
            sine_reg0   <= 36'sb111000110011110010110001111000010101;
        end
        8784: begin
            cosine_reg0 <= 36'sb100000110100100011011000110110111111;
            sine_reg0   <= 36'sb111000110011000001110011010011001111;
        end
        8785: begin
            cosine_reg0 <= 36'sb100000110100101110101101100011011001;
            sine_reg0   <= 36'sb111000110010010000110100111111111010;
        end
        8786: begin
            cosine_reg0 <= 36'sb100000110100111010000011011100101110;
            sine_reg0   <= 36'sb111000110001011111110110111110011000;
        end
        8787: begin
            cosine_reg0 <= 36'sb100000110101000101011010100010111110;
            sine_reg0   <= 36'sb111000110000101110111001001110101100;
        end
        8788: begin
            cosine_reg0 <= 36'sb100000110101010000110010110110001001;
            sine_reg0   <= 36'sb111000101111111101111011110000110111;
        end
        8789: begin
            cosine_reg0 <= 36'sb100000110101011100001100010110001101;
            sine_reg0   <= 36'sb111000101111001100111110100100111010;
        end
        8790: begin
            cosine_reg0 <= 36'sb100000110101100111100111000011001010;
            sine_reg0   <= 36'sb111000101110011100000001101010111001;
        end
        8791: begin
            cosine_reg0 <= 36'sb100000110101110011000010111101000001;
            sine_reg0   <= 36'sb111000101101101011000101000010110100;
        end
        8792: begin
            cosine_reg0 <= 36'sb100000110101111110100000000011101111;
            sine_reg0   <= 36'sb111000101100111010001000101100101101;
        end
        8793: begin
            cosine_reg0 <= 36'sb100000110110001001111110010111010110;
            sine_reg0   <= 36'sb111000101100001001001100101000101000;
        end
        8794: begin
            cosine_reg0 <= 36'sb100000110110010101011101110111110101;
            sine_reg0   <= 36'sb111000101011011000010000110110100100;
        end
        8795: begin
            cosine_reg0 <= 36'sb100000110110100000111110100101001011;
            sine_reg0   <= 36'sb111000101010100111010101010110100101;
        end
        8796: begin
            cosine_reg0 <= 36'sb100000110110101100100000011111010111;
            sine_reg0   <= 36'sb111000101001110110011010001000101100;
        end
        8797: begin
            cosine_reg0 <= 36'sb100000110110111000000011100110011010;
            sine_reg0   <= 36'sb111000101001000101011111001100111011;
        end
        8798: begin
            cosine_reg0 <= 36'sb100000110111000011100111111010010011;
            sine_reg0   <= 36'sb111000101000010100100100100011010100;
        end
        8799: begin
            cosine_reg0 <= 36'sb100000110111001111001101011011000000;
            sine_reg0   <= 36'sb111000100111100011101010001011111001;
        end
        8800: begin
            cosine_reg0 <= 36'sb100000110111011010110100001000100011;
            sine_reg0   <= 36'sb111000100110110010110000000110101100;
        end
        8801: begin
            cosine_reg0 <= 36'sb100000110111100110011100000010111011;
            sine_reg0   <= 36'sb111000100110000001110110010011101110;
        end
        8802: begin
            cosine_reg0 <= 36'sb100000110111110010000101001010000110;
            sine_reg0   <= 36'sb111000100101010000111100110011000010;
        end
        8803: begin
            cosine_reg0 <= 36'sb100000110111111101101111011110000101;
            sine_reg0   <= 36'sb111000100100100000000011100100101001;
        end
        8804: begin
            cosine_reg0 <= 36'sb100000111000001001011010111110111000;
            sine_reg0   <= 36'sb111000100011101111001010101000100101;
        end
        8805: begin
            cosine_reg0 <= 36'sb100000111000010101000111101100011100;
            sine_reg0   <= 36'sb111000100010111110010001111110111000;
        end
        8806: begin
            cosine_reg0 <= 36'sb100000111000100000110101100110110100;
            sine_reg0   <= 36'sb111000100010001101011001100111100101;
        end
        8807: begin
            cosine_reg0 <= 36'sb100000111000101100100100101101111101;
            sine_reg0   <= 36'sb111000100001011100100001100010101100;
        end
        8808: begin
            cosine_reg0 <= 36'sb100000111000111000010101000001110111;
            sine_reg0   <= 36'sb111000100000101011101001110000010000;
        end
        8809: begin
            cosine_reg0 <= 36'sb100000111001000100000110100010100010;
            sine_reg0   <= 36'sb111000011111111010110010010000010011;
        end
        8810: begin
            cosine_reg0 <= 36'sb100000111001001111111001001111111110;
            sine_reg0   <= 36'sb111000011111001001111011000010110110;
        end
        8811: begin
            cosine_reg0 <= 36'sb100000111001011011101101001010001001;
            sine_reg0   <= 36'sb111000011110011001000100000111111100;
        end
        8812: begin
            cosine_reg0 <= 36'sb100000111001100111100010010001000100;
            sine_reg0   <= 36'sb111000011101101000001101011111100110;
        end
        8813: begin
            cosine_reg0 <= 36'sb100000111001110011011000100100101111;
            sine_reg0   <= 36'sb111000011100110111010111001001110110;
        end
        8814: begin
            cosine_reg0 <= 36'sb100000111001111111010000000101001000;
            sine_reg0   <= 36'sb111000011100000110100001000110101111;
        end
        8815: begin
            cosine_reg0 <= 36'sb100000111010001011001000110010001111;
            sine_reg0   <= 36'sb111000011011010101101011010110010001;
        end
        8816: begin
            cosine_reg0 <= 36'sb100000111010010111000010101100000011;
            sine_reg0   <= 36'sb111000011010100100110101111000011111;
        end
        8817: begin
            cosine_reg0 <= 36'sb100000111010100010111101110010100101;
            sine_reg0   <= 36'sb111000011001110100000000101101011011;
        end
        8818: begin
            cosine_reg0 <= 36'sb100000111010101110111010000101110100;
            sine_reg0   <= 36'sb111000011001000011001011110101000111;
        end
        8819: begin
            cosine_reg0 <= 36'sb100000111010111010110111100101101111;
            sine_reg0   <= 36'sb111000011000010010010111001111100100;
        end
        8820: begin
            cosine_reg0 <= 36'sb100000111011000110110110010010010110;
            sine_reg0   <= 36'sb111000010111100001100010111100110100;
        end
        8821: begin
            cosine_reg0 <= 36'sb100000111011010010110110001011101000;
            sine_reg0   <= 36'sb111000010110110000101110111100111010;
        end
        8822: begin
            cosine_reg0 <= 36'sb100000111011011110110111010001100101;
            sine_reg0   <= 36'sb111000010101111111111011001111110111;
        end
        8823: begin
            cosine_reg0 <= 36'sb100000111011101010111001100100001101;
            sine_reg0   <= 36'sb111000010101001111000111110101101101;
        end
        8824: begin
            cosine_reg0 <= 36'sb100000111011110110111101000011011111;
            sine_reg0   <= 36'sb111000010100011110010100101110011101;
        end
        8825: begin
            cosine_reg0 <= 36'sb100000111100000011000001101111011010;
            sine_reg0   <= 36'sb111000010011101101100001111010001011;
        end
        8826: begin
            cosine_reg0 <= 36'sb100000111100001111000111100111111110;
            sine_reg0   <= 36'sb111000010010111100101111011000110111;
        end
        8827: begin
            cosine_reg0 <= 36'sb100000111100011011001110101101001011;
            sine_reg0   <= 36'sb111000010010001011111101001010100100;
        end
        8828: begin
            cosine_reg0 <= 36'sb100000111100100111010110111111000000;
            sine_reg0   <= 36'sb111000010001011011001011001111010011;
        end
        8829: begin
            cosine_reg0 <= 36'sb100000111100110011100000011101011101;
            sine_reg0   <= 36'sb111000010000101010011001100111000111;
        end
        8830: begin
            cosine_reg0 <= 36'sb100000111100111111101011001000100001;
            sine_reg0   <= 36'sb111000001111111001101000010010000001;
        end
        8831: begin
            cosine_reg0 <= 36'sb100000111101001011110111000000001011;
            sine_reg0   <= 36'sb111000001111001000110111010000000010;
        end
        8832: begin
            cosine_reg0 <= 36'sb100000111101011000000100000100011100;
            sine_reg0   <= 36'sb111000001110011000000110100001001110;
        end
        8833: begin
            cosine_reg0 <= 36'sb100000111101100100010010010101010011;
            sine_reg0   <= 36'sb111000001101100111010110000101100110;
        end
        8834: begin
            cosine_reg0 <= 36'sb100000111101110000100001110010101111;
            sine_reg0   <= 36'sb111000001100110110100101111101001011;
        end
        8835: begin
            cosine_reg0 <= 36'sb100000111101111100110010011100110000;
            sine_reg0   <= 36'sb111000001100000101110110001000000000;
        end
        8836: begin
            cosine_reg0 <= 36'sb100000111110001001000100010011010101;
            sine_reg0   <= 36'sb111000001011010101000110100110000110;
        end
        8837: begin
            cosine_reg0 <= 36'sb100000111110010101010111010110011111;
            sine_reg0   <= 36'sb111000001010100100010111010111100000;
        end
        8838: begin
            cosine_reg0 <= 36'sb100000111110100001101011100110001011;
            sine_reg0   <= 36'sb111000001001110011101000011100001111;
        end
        8839: begin
            cosine_reg0 <= 36'sb100000111110101110000001000010011011;
            sine_reg0   <= 36'sb111000001001000010111001110100010101;
        end
        8840: begin
            cosine_reg0 <= 36'sb100000111110111010010111101011001101;
            sine_reg0   <= 36'sb111000001000010010001011011111110100;
        end
        8841: begin
            cosine_reg0 <= 36'sb100000111111000110101111100000100001;
            sine_reg0   <= 36'sb111000000111100001011101011110101110;
        end
        8842: begin
            cosine_reg0 <= 36'sb100000111111010011001000100010010111;
            sine_reg0   <= 36'sb111000000110110000101111110001000101;
        end
        8843: begin
            cosine_reg0 <= 36'sb100000111111011111100010110000101110;
            sine_reg0   <= 36'sb111000000110000000000010010110111010;
        end
        8844: begin
            cosine_reg0 <= 36'sb100000111111101011111110001011100101;
            sine_reg0   <= 36'sb111000000101001111010101010000010000;
        end
        8845: begin
            cosine_reg0 <= 36'sb100000111111111000011010110010111100;
            sine_reg0   <= 36'sb111000000100011110101000011101001001;
        end
        8846: begin
            cosine_reg0 <= 36'sb100001000000000100111000100110110011;
            sine_reg0   <= 36'sb111000000011101101111011111101100101;
        end
        8847: begin
            cosine_reg0 <= 36'sb100001000000010001010111100111001001;
            sine_reg0   <= 36'sb111000000010111101001111110001101000;
        end
        8848: begin
            cosine_reg0 <= 36'sb100001000000011101110111110011111110;
            sine_reg0   <= 36'sb111000000010001100100011111001010010;
        end
        8849: begin
            cosine_reg0 <= 36'sb100001000000101010011001001101010001;
            sine_reg0   <= 36'sb111000000001011011111000010100100111;
        end
        8850: begin
            cosine_reg0 <= 36'sb100001000000110110111011110011000010;
            sine_reg0   <= 36'sb111000000000101011001101000011100111;
        end
        8851: begin
            cosine_reg0 <= 36'sb100001000001000011011111100101001111;
            sine_reg0   <= 36'sb110111111111111010100010000110010101;
        end
        8852: begin
            cosine_reg0 <= 36'sb100001000001010000000100100011111010;
            sine_reg0   <= 36'sb110111111111001001110111011100110010;
        end
        8853: begin
            cosine_reg0 <= 36'sb100001000001011100101010101111000001;
            sine_reg0   <= 36'sb110111111110011001001101000111000001;
        end
        8854: begin
            cosine_reg0 <= 36'sb100001000001101001010010000110100011;
            sine_reg0   <= 36'sb110111111101101000100011000101000011;
        end
        8855: begin
            cosine_reg0 <= 36'sb100001000001110101111010101010100001;
            sine_reg0   <= 36'sb110111111100110111111001010110111011;
        end
        8856: begin
            cosine_reg0 <= 36'sb100001000010000010100100011010111010;
            sine_reg0   <= 36'sb110111111100000111001111111100101001;
        end
        8857: begin
            cosine_reg0 <= 36'sb100001000010001111001111010111101101;
            sine_reg0   <= 36'sb110111111011010110100110110110010000;
        end
        8858: begin
            cosine_reg0 <= 36'sb100001000010011011111011100000111001;
            sine_reg0   <= 36'sb110111111010100101111110000011110010;
        end
        8859: begin
            cosine_reg0 <= 36'sb100001000010101000101000110110011111;
            sine_reg0   <= 36'sb110111111001110101010101100101010001;
        end
        8860: begin
            cosine_reg0 <= 36'sb100001000010110101010111011000011110;
            sine_reg0   <= 36'sb110111111001000100101101011010101110;
        end
        8861: begin
            cosine_reg0 <= 36'sb100001000011000010000111000110110101;
            sine_reg0   <= 36'sb110111111000010100000101100100001011;
        end
        8862: begin
            cosine_reg0 <= 36'sb100001000011001110111000000001100100;
            sine_reg0   <= 36'sb110111110111100011011110000001101011;
        end
        8863: begin
            cosine_reg0 <= 36'sb100001000011011011101010001000101011;
            sine_reg0   <= 36'sb110111110110110010110110110011001111;
        end
        8864: begin
            cosine_reg0 <= 36'sb100001000011101000011101011100001000;
            sine_reg0   <= 36'sb110111110110000010001111111000111001;
        end
        8865: begin
            cosine_reg0 <= 36'sb100001000011110101010001111011111011;
            sine_reg0   <= 36'sb110111110101010001101001010010101011;
        end
        8866: begin
            cosine_reg0 <= 36'sb100001000100000010000111101000000101;
            sine_reg0   <= 36'sb110111110100100001000011000000100111;
        end
        8867: begin
            cosine_reg0 <= 36'sb100001000100001110111110100000100100;
            sine_reg0   <= 36'sb110111110011110000011101000010101110;
        end
        8868: begin
            cosine_reg0 <= 36'sb100001000100011011110110100101010111;
            sine_reg0   <= 36'sb110111110010111111110111011001000011;
        end
        8869: begin
            cosine_reg0 <= 36'sb100001000100101000101111110110011111;
            sine_reg0   <= 36'sb110111110010001111010010000011100111;
        end
        8870: begin
            cosine_reg0 <= 36'sb100001000100110101101010010011111011;
            sine_reg0   <= 36'sb110111110001011110101101000010011101;
        end
        8871: begin
            cosine_reg0 <= 36'sb100001000101000010100101111101101011;
            sine_reg0   <= 36'sb110111110000101110001000010101100101;
        end
        8872: begin
            cosine_reg0 <= 36'sb100001000101001111100010110011101101;
            sine_reg0   <= 36'sb110111101111111101100011111101000011;
        end
        8873: begin
            cosine_reg0 <= 36'sb100001000101011100100000110110000001;
            sine_reg0   <= 36'sb110111101111001100111111111000110111;
        end
        8874: begin
            cosine_reg0 <= 36'sb100001000101101001100000000100101000;
            sine_reg0   <= 36'sb110111101110011100011100001001000101;
        end
        8875: begin
            cosine_reg0 <= 36'sb100001000101110110100000011111100000;
            sine_reg0   <= 36'sb110111101101101011111000101101101100;
        end
        8876: begin
            cosine_reg0 <= 36'sb100001000110000011100010000110101001;
            sine_reg0   <= 36'sb110111101100111011010101100110110001;
        end
        8877: begin
            cosine_reg0 <= 36'sb100001000110010000100100111010000010;
            sine_reg0   <= 36'sb110111101100001010110010110100010100;
        end
        8878: begin
            cosine_reg0 <= 36'sb100001000110011101101000111001101011;
            sine_reg0   <= 36'sb110111101011011010010000010110010111;
        end
        8879: begin
            cosine_reg0 <= 36'sb100001000110101010101110000101100011;
            sine_reg0   <= 36'sb110111101010101001101110001100111100;
        end
        8880: begin
            cosine_reg0 <= 36'sb100001000110110111110100011101101010;
            sine_reg0   <= 36'sb110111101001111001001100011000000101;
        end
        8881: begin
            cosine_reg0 <= 36'sb100001000111000100111100000010000000;
            sine_reg0   <= 36'sb110111101001001000101010110111110100;
        end
        8882: begin
            cosine_reg0 <= 36'sb100001000111010010000100110010100011;
            sine_reg0   <= 36'sb110111101000011000001001101100001010;
        end
        8883: begin
            cosine_reg0 <= 36'sb100001000111011111001110101111010100;
            sine_reg0   <= 36'sb110111100111100111101000110101001011;
        end
        8884: begin
            cosine_reg0 <= 36'sb100001000111101100011001111000010010;
            sine_reg0   <= 36'sb110111100110110111001000010010110110;
        end
        8885: begin
            cosine_reg0 <= 36'sb100001000111111001100110001101011100;
            sine_reg0   <= 36'sb110111100110000110101000000101001111;
        end
        8886: begin
            cosine_reg0 <= 36'sb100001001000000110110011101110110010;
            sine_reg0   <= 36'sb110111100101010110001000001100011000;
        end
        8887: begin
            cosine_reg0 <= 36'sb100001001000010100000010011100010011;
            sine_reg0   <= 36'sb110111100100100101101000101000010001;
        end
        8888: begin
            cosine_reg0 <= 36'sb100001001000100001010010010101111111;
            sine_reg0   <= 36'sb110111100011110101001001011000111101;
        end
        8889: begin
            cosine_reg0 <= 36'sb100001001000101110100011011011110101;
            sine_reg0   <= 36'sb110111100011000100101010011110011110;
        end
        8890: begin
            cosine_reg0 <= 36'sb100001001000111011110101101101110101;
            sine_reg0   <= 36'sb110111100010010100001011111000110110;
        end
        8891: begin
            cosine_reg0 <= 36'sb100001001001001001001001001011111111;
            sine_reg0   <= 36'sb110111100001100011101101101000000111;
        end
        8892: begin
            cosine_reg0 <= 36'sb100001001001010110011101110110010001;
            sine_reg0   <= 36'sb110111100000110011001111101100010001;
        end
        8893: begin
            cosine_reg0 <= 36'sb100001001001100011110011101100101011;
            sine_reg0   <= 36'sb110111100000000010110010000101011000;
        end
        8894: begin
            cosine_reg0 <= 36'sb100001001001110001001010101111001101;
            sine_reg0   <= 36'sb110111011111010010010100110011011110;
        end
        8895: begin
            cosine_reg0 <= 36'sb100001001001111110100010111101110111;
            sine_reg0   <= 36'sb110111011110100001110111110110100011;
        end
        8896: begin
            cosine_reg0 <= 36'sb100001001010001011111100011000100111;
            sine_reg0   <= 36'sb110111011101110001011011001110101010;
        end
        8897: begin
            cosine_reg0 <= 36'sb100001001010011001010110111111011101;
            sine_reg0   <= 36'sb110111011101000000111110111011110101;
        end
        8898: begin
            cosine_reg0 <= 36'sb100001001010100110110010110010011001;
            sine_reg0   <= 36'sb110111011100010000100010111110000101;
        end
        8899: begin
            cosine_reg0 <= 36'sb100001001010110100001111110001011010;
            sine_reg0   <= 36'sb110111011011100000000111010101011101;
        end
        8900: begin
            cosine_reg0 <= 36'sb100001001011000001101101111100100000;
            sine_reg0   <= 36'sb110111011010101111101100000001111111;
        end
        8901: begin
            cosine_reg0 <= 36'sb100001001011001111001101010011101010;
            sine_reg0   <= 36'sb110111011001111111010001000011101100;
        end
        8902: begin
            cosine_reg0 <= 36'sb100001001011011100101101110110110111;
            sine_reg0   <= 36'sb110111011001001110110110011010100101;
        end
        8903: begin
            cosine_reg0 <= 36'sb100001001011101010001111100110001000;
            sine_reg0   <= 36'sb110111011000011110011100000110101110;
        end
        8904: begin
            cosine_reg0 <= 36'sb100001001011110111110010100001011011;
            sine_reg0   <= 36'sb110111010111101110000010001000000111;
        end
        8905: begin
            cosine_reg0 <= 36'sb100001001100000101010110101000110000;
            sine_reg0   <= 36'sb110111010110111101101000011110110100;
        end
        8906: begin
            cosine_reg0 <= 36'sb100001001100010010111011111100000110;
            sine_reg0   <= 36'sb110111010110001101001111001010110100;
        end
        8907: begin
            cosine_reg0 <= 36'sb100001001100100000100010011011011110;
            sine_reg0   <= 36'sb110111010101011100110110001100001100;
        end
        8908: begin
            cosine_reg0 <= 36'sb100001001100101110001010000110110110;
            sine_reg0   <= 36'sb110111010100101100011101100010111011;
        end
        8909: begin
            cosine_reg0 <= 36'sb100001001100111011110010111110001110;
            sine_reg0   <= 36'sb110111010011111100000101001111000101;
        end
        8910: begin
            cosine_reg0 <= 36'sb100001001101001001011101000001100101;
            sine_reg0   <= 36'sb110111010011001011101101010000101011;
        end
        8911: begin
            cosine_reg0 <= 36'sb100001001101010111001000010000111011;
            sine_reg0   <= 36'sb110111010010011011010101100111101110;
        end
        8912: begin
            cosine_reg0 <= 36'sb100001001101100100110100101100010000;
            sine_reg0   <= 36'sb110111010001101010111110010100010001;
        end
        8913: begin
            cosine_reg0 <= 36'sb100001001101110010100010010011100010;
            sine_reg0   <= 36'sb110111010000111010100111010110010110;
        end
        8914: begin
            cosine_reg0 <= 36'sb100001001110000000010001000110110010;
            sine_reg0   <= 36'sb110111010000001010010000101101111111;
        end
        8915: begin
            cosine_reg0 <= 36'sb100001001110001110000001000101111111;
            sine_reg0   <= 36'sb110111001111011001111010011011001101;
        end
        8916: begin
            cosine_reg0 <= 36'sb100001001110011011110010010001000111;
            sine_reg0   <= 36'sb110111001110101001100100011110000010;
        end
        8917: begin
            cosine_reg0 <= 36'sb100001001110101001100100101000001100;
            sine_reg0   <= 36'sb110111001101111001001110110110100000;
        end
        8918: begin
            cosine_reg0 <= 36'sb100001001110110111011000001011001100;
            sine_reg0   <= 36'sb110111001101001000111001100100101001;
        end
        8919: begin
            cosine_reg0 <= 36'sb100001001111000101001100111010000110;
            sine_reg0   <= 36'sb110111001100011000100100101000011111;
        end
        8920: begin
            cosine_reg0 <= 36'sb100001001111010011000010110100111010;
            sine_reg0   <= 36'sb110111001011101000010000000010000011;
        end
        8921: begin
            cosine_reg0 <= 36'sb100001001111100000111001111011101000;
            sine_reg0   <= 36'sb110111001010110111111011110001011000;
        end
        8922: begin
            cosine_reg0 <= 36'sb100001001111101110110010001110001111;
            sine_reg0   <= 36'sb110111001010000111100111110110100000;
        end
        8923: begin
            cosine_reg0 <= 36'sb100001001111111100101011101100101111;
            sine_reg0   <= 36'sb110111001001010111010100010001011011;
        end
        8924: begin
            cosine_reg0 <= 36'sb100001010000001010100110010111000110;
            sine_reg0   <= 36'sb110111001000100111000001000010001101;
        end
        8925: begin
            cosine_reg0 <= 36'sb100001010000011000100010001101010101;
            sine_reg0   <= 36'sb110111000111110110101110001000110111;
        end
        8926: begin
            cosine_reg0 <= 36'sb100001010000100110011111001111011011;
            sine_reg0   <= 36'sb110111000111000110011011100101011010;
        end
        8927: begin
            cosine_reg0 <= 36'sb100001010000110100011101011101010111;
            sine_reg0   <= 36'sb110111000110010110001001010111111010;
        end
        8928: begin
            cosine_reg0 <= 36'sb100001010001000010011100110111001001;
            sine_reg0   <= 36'sb110111000101100101110111100000010111;
        end
        8929: begin
            cosine_reg0 <= 36'sb100001010001010000011101011100110000;
            sine_reg0   <= 36'sb110111000100110101100101111110110011;
        end
        8930: begin
            cosine_reg0 <= 36'sb100001010001011110011111001110001101;
            sine_reg0   <= 36'sb110111000100000101010100110011010001;
        end
        8931: begin
            cosine_reg0 <= 36'sb100001010001101100100010001011011101;
            sine_reg0   <= 36'sb110111000011010101000011111101110001;
        end
        8932: begin
            cosine_reg0 <= 36'sb100001010001111010100110010100100001;
            sine_reg0   <= 36'sb110111000010100100110011011110010111;
        end
        8933: begin
            cosine_reg0 <= 36'sb100001010010001000101011101001011000;
            sine_reg0   <= 36'sb110111000001110100100011010101000100;
        end
        8934: begin
            cosine_reg0 <= 36'sb100001010010010110110010001010000001;
            sine_reg0   <= 36'sb110111000001000100010011100001111001;
        end
        8935: begin
            cosine_reg0 <= 36'sb100001010010100100111001110110011101;
            sine_reg0   <= 36'sb110111000000010100000100000100111001;
        end
        8936: begin
            cosine_reg0 <= 36'sb100001010010110011000010101110101010;
            sine_reg0   <= 36'sb110110111111100011110100111110000101;
        end
        8937: begin
            cosine_reg0 <= 36'sb100001010011000001001100110010101000;
            sine_reg0   <= 36'sb110110111110110011100110001101100000;
        end
        8938: begin
            cosine_reg0 <= 36'sb100001010011001111011000000010010111;
            sine_reg0   <= 36'sb110110111110000011010111110011001011;
        end
        8939: begin
            cosine_reg0 <= 36'sb100001010011011101100100011101110101;
            sine_reg0   <= 36'sb110110111101010011001001101111001000;
        end
        8940: begin
            cosine_reg0 <= 36'sb100001010011101011110010000101000011;
            sine_reg0   <= 36'sb110110111100100010111100000001011001;
        end
        8941: begin
            cosine_reg0 <= 36'sb100001010011111010000000110111111111;
            sine_reg0   <= 36'sb110110111011110010101110101001111111;
        end
        8942: begin
            cosine_reg0 <= 36'sb100001010100001000010000110110101001;
            sine_reg0   <= 36'sb110110111011000010100001101000111101;
        end
        8943: begin
            cosine_reg0 <= 36'sb100001010100010110100010000001000010;
            sine_reg0   <= 36'sb110110111010010010010100111110010101;
        end
        8944: begin
            cosine_reg0 <= 36'sb100001010100100100110100010111000111;
            sine_reg0   <= 36'sb110110111001100010001000101010001000;
        end
        8945: begin
            cosine_reg0 <= 36'sb100001010100110011000111111000111001;
            sine_reg0   <= 36'sb110110111000110001111100101100011000;
        end
        8946: begin
            cosine_reg0 <= 36'sb100001010101000001011100100110010111;
            sine_reg0   <= 36'sb110110111000000001110001000101000111;
        end
        8947: begin
            cosine_reg0 <= 36'sb100001010101001111110010011111100000;
            sine_reg0   <= 36'sb110110110111010001100101110100010111;
        end
        8948: begin
            cosine_reg0 <= 36'sb100001010101011110001001100100010100;
            sine_reg0   <= 36'sb110110110110100001011010111010001010;
        end
        8949: begin
            cosine_reg0 <= 36'sb100001010101101100100001110100110011;
            sine_reg0   <= 36'sb110110110101110001010000010110100001;
        end
        8950: begin
            cosine_reg0 <= 36'sb100001010101111010111011010000111011;
            sine_reg0   <= 36'sb110110110101000001000110001001011111;
        end
        8951: begin
            cosine_reg0 <= 36'sb100001010110001001010101111000101101;
            sine_reg0   <= 36'sb110110110100010000111100010011000101;
        end
        8952: begin
            cosine_reg0 <= 36'sb100001010110010111110001101100000111;
            sine_reg0   <= 36'sb110110110011100000110010110011010110;
        end
        8953: begin
            cosine_reg0 <= 36'sb100001010110100110001110101011001010;
            sine_reg0   <= 36'sb110110110010110000101001101010010010;
        end
        8954: begin
            cosine_reg0 <= 36'sb100001010110110100101100110101110100;
            sine_reg0   <= 36'sb110110110010000000100000110111111100;
        end
        8955: begin
            cosine_reg0 <= 36'sb100001010111000011001100001100000101;
            sine_reg0   <= 36'sb110110110001010000011000011100010110;
        end
        8956: begin
            cosine_reg0 <= 36'sb100001010111010001101100101101111100;
            sine_reg0   <= 36'sb110110110000100000010000010111100010;
        end
        8957: begin
            cosine_reg0 <= 36'sb100001010111100000001110011011011010;
            sine_reg0   <= 36'sb110110101111110000001000101001100001;
        end
        8958: begin
            cosine_reg0 <= 36'sb100001010111101110110001010100011100;
            sine_reg0   <= 36'sb110110101111000000000001010010010101;
        end
        8959: begin
            cosine_reg0 <= 36'sb100001010111111101010101011001000100;
            sine_reg0   <= 36'sb110110101110001111111010010010000001;
        end
        8960: begin
            cosine_reg0 <= 36'sb100001011000001011111010101001001111;
            sine_reg0   <= 36'sb110110101101011111110011101000100110;
        end
        8961: begin
            cosine_reg0 <= 36'sb100001011000011010100001000100111111;
            sine_reg0   <= 36'sb110110101100101111101101010110000101;
        end
        8962: begin
            cosine_reg0 <= 36'sb100001011000101001001000101100010001;
            sine_reg0   <= 36'sb110110101011111111100111011010100001;
        end
        8963: begin
            cosine_reg0 <= 36'sb100001011000110111110001011111000110;
            sine_reg0   <= 36'sb110110101011001111100001110101111100;
        end
        8964: begin
            cosine_reg0 <= 36'sb100001011001000110011011011101011101;
            sine_reg0   <= 36'sb110110101010011111011100101000010111;
        end
        8965: begin
            cosine_reg0 <= 36'sb100001011001010101000110100111010101;
            sine_reg0   <= 36'sb110110101001101111010111110001110101;
        end
        8966: begin
            cosine_reg0 <= 36'sb100001011001100011110010111100101110;
            sine_reg0   <= 36'sb110110101000111111010011010010010110;
        end
        8967: begin
            cosine_reg0 <= 36'sb100001011001110010100000011101101000;
            sine_reg0   <= 36'sb110110101000001111001111001001111110;
        end
        8968: begin
            cosine_reg0 <= 36'sb100001011010000001001111001010000001;
            sine_reg0   <= 36'sb110110100111011111001011011000101110;
        end
        8969: begin
            cosine_reg0 <= 36'sb100001011010001111111111000001111001;
            sine_reg0   <= 36'sb110110100110101111000111111110100111;
        end
        8970: begin
            cosine_reg0 <= 36'sb100001011010011110110000000101001111;
            sine_reg0   <= 36'sb110110100101111111000100111011101100;
        end
        8971: begin
            cosine_reg0 <= 36'sb100001011010101101100010010100000100;
            sine_reg0   <= 36'sb110110100101001111000010001111111110;
        end
        8972: begin
            cosine_reg0 <= 36'sb100001011010111100010101101110010110;
            sine_reg0   <= 36'sb110110100100011110111111111011011111;
        end
        8973: begin
            cosine_reg0 <= 36'sb100001011011001011001010010100000101;
            sine_reg0   <= 36'sb110110100011101110111101111110010010;
        end
        8974: begin
            cosine_reg0 <= 36'sb100001011011011010000000000101010000;
            sine_reg0   <= 36'sb110110100010111110111100011000010111;
        end
        8975: begin
            cosine_reg0 <= 36'sb100001011011101000110111000001110111;
            sine_reg0   <= 36'sb110110100010001110111011001001110010;
        end
        8976: begin
            cosine_reg0 <= 36'sb100001011011110111101111001001111001;
            sine_reg0   <= 36'sb110110100001011110111010010010100011;
        end
        8977: begin
            cosine_reg0 <= 36'sb100001011100000110101000011101010110;
            sine_reg0   <= 36'sb110110100000101110111001110010101100;
        end
        8978: begin
            cosine_reg0 <= 36'sb100001011100010101100010111100001101;
            sine_reg0   <= 36'sb110110011111111110111001101010010000;
        end
        8979: begin
            cosine_reg0 <= 36'sb100001011100100100011110100110011101;
            sine_reg0   <= 36'sb110110011111001110111001111001010000;
        end
        8980: begin
            cosine_reg0 <= 36'sb100001011100110011011011011100000110;
            sine_reg0   <= 36'sb110110011110011110111010011111101111;
        end
        8981: begin
            cosine_reg0 <= 36'sb100001011101000010011001011101000111;
            sine_reg0   <= 36'sb110110011101101110111011011101101101;
        end
        8982: begin
            cosine_reg0 <= 36'sb100001011101010001011000101001011111;
            sine_reg0   <= 36'sb110110011100111110111100110011001101;
        end
        8983: begin
            cosine_reg0 <= 36'sb100001011101100000011001000001001111;
            sine_reg0   <= 36'sb110110011100001110111110100000010000;
        end
        8984: begin
            cosine_reg0 <= 36'sb100001011101101111011010100100010110;
            sine_reg0   <= 36'sb110110011011011111000000100100111001;
        end
        8985: begin
            cosine_reg0 <= 36'sb100001011101111110011101010010110010;
            sine_reg0   <= 36'sb110110011010101111000011000001001010;
        end
        8986: begin
            cosine_reg0 <= 36'sb100001011110001101100001001100100100;
            sine_reg0   <= 36'sb110110011001111111000101110101000011;
        end
        8987: begin
            cosine_reg0 <= 36'sb100001011110011100100110010001101010;
            sine_reg0   <= 36'sb110110011001001111001001000000101000;
        end
        8988: begin
            cosine_reg0 <= 36'sb100001011110101011101100100010000101;
            sine_reg0   <= 36'sb110110011000011111001100100011111001;
        end
        8989: begin
            cosine_reg0 <= 36'sb100001011110111010110011111101110011;
            sine_reg0   <= 36'sb110110010111101111010000011110111001;
        end
        8990: begin
            cosine_reg0 <= 36'sb100001011111001001111100100100110100;
            sine_reg0   <= 36'sb110110010110111111010100110001101010;
        end
        8991: begin
            cosine_reg0 <= 36'sb100001011111011001000110010111001000;
            sine_reg0   <= 36'sb110110010110001111011001011100001101;
        end
        8992: begin
            cosine_reg0 <= 36'sb100001011111101000010001010100101110;
            sine_reg0   <= 36'sb110110010101011111011110011110100100;
        end
        8993: begin
            cosine_reg0 <= 36'sb100001011111110111011101011101100101;
            sine_reg0   <= 36'sb110110010100101111100011111000110010;
        end
        8994: begin
            cosine_reg0 <= 36'sb100001100000000110101010110001101100;
            sine_reg0   <= 36'sb110110010011111111101001101010110111;
        end
        8995: begin
            cosine_reg0 <= 36'sb100001100000010101111001010001000100;
            sine_reg0   <= 36'sb110110010011001111101111110100110110;
        end
        8996: begin
            cosine_reg0 <= 36'sb100001100000100101001000111011101011;
            sine_reg0   <= 36'sb110110010010011111110110010110110001;
        end
        8997: begin
            cosine_reg0 <= 36'sb100001100000110100011001110001100001;
            sine_reg0   <= 36'sb110110010001101111111101010000101001;
        end
        8998: begin
            cosine_reg0 <= 36'sb100001100001000011101011110010100110;
            sine_reg0   <= 36'sb110110010001000000000100100010100001;
        end
        8999: begin
            cosine_reg0 <= 36'sb100001100001010010111110111110111000;
            sine_reg0   <= 36'sb110110010000010000001100001100011010;
        end
        9000: begin
            cosine_reg0 <= 36'sb100001100001100010010011010110011000;
            sine_reg0   <= 36'sb110110001111100000010100001110010110;
        end
        9001: begin
            cosine_reg0 <= 36'sb100001100001110001101000111001000100;
            sine_reg0   <= 36'sb110110001110110000011100101000010111;
        end
        9002: begin
            cosine_reg0 <= 36'sb100001100010000000111111100110111100;
            sine_reg0   <= 36'sb110110001110000000100101011010011110;
        end
        9003: begin
            cosine_reg0 <= 36'sb100001100010010000010111011111111111;
            sine_reg0   <= 36'sb110110001101010000101110100100101110;
        end
        9004: begin
            cosine_reg0 <= 36'sb100001100010011111110000100100001101;
            sine_reg0   <= 36'sb110110001100100000111000000111001001;
        end
        9005: begin
            cosine_reg0 <= 36'sb100001100010101111001010110011100110;
            sine_reg0   <= 36'sb110110001011110001000010000001110000;
        end
        9006: begin
            cosine_reg0 <= 36'sb100001100010111110100110001110001000;
            sine_reg0   <= 36'sb110110001011000001001100010100100100;
        end
        9007: begin
            cosine_reg0 <= 36'sb100001100011001110000010110011110011;
            sine_reg0   <= 36'sb110110001010010001010110111111101001;
        end
        9008: begin
            cosine_reg0 <= 36'sb100001100011011101100000100100100110;
            sine_reg0   <= 36'sb110110001001100001100010000011000000;
        end
        9009: begin
            cosine_reg0 <= 36'sb100001100011101100111111100000100010;
            sine_reg0   <= 36'sb110110001000110001101101011110101010;
        end
        9010: begin
            cosine_reg0 <= 36'sb100001100011111100011111100111100100;
            sine_reg0   <= 36'sb110110001000000001111001010010101010;
        end
        9011: begin
            cosine_reg0 <= 36'sb100001100100001100000000111001101101;
            sine_reg0   <= 36'sb110110000111010010000101011111000001;
        end
        9012: begin
            cosine_reg0 <= 36'sb100001100100011011100011010110111100;
            sine_reg0   <= 36'sb110110000110100010010010000011110001;
        end
        9013: begin
            cosine_reg0 <= 36'sb100001100100101011000110111111010001;
            sine_reg0   <= 36'sb110110000101110010011111000000111100;
        end
        9014: begin
            cosine_reg0 <= 36'sb100001100100111010101011110010101011;
            sine_reg0   <= 36'sb110110000101000010101100010110100100;
        end
        9015: begin
            cosine_reg0 <= 36'sb100001100101001010010001110001001000;
            sine_reg0   <= 36'sb110110000100010010111010000100101011;
        end
        9016: begin
            cosine_reg0 <= 36'sb100001100101011001111000111010101010;
            sine_reg0   <= 36'sb110110000011100011001000001011010010;
        end
        9017: begin
            cosine_reg0 <= 36'sb100001100101101001100001001111001110;
            sine_reg0   <= 36'sb110110000010110011010110101010011100;
        end
        9018: begin
            cosine_reg0 <= 36'sb100001100101111001001010101110110101;
            sine_reg0   <= 36'sb110110000010000011100101100010001010;
        end
        9019: begin
            cosine_reg0 <= 36'sb100001100110001000110101011001011101;
            sine_reg0   <= 36'sb110110000001010011110100110010011110;
        end
        9020: begin
            cosine_reg0 <= 36'sb100001100110011000100001001111000111;
            sine_reg0   <= 36'sb110110000000100100000100011011011010;
        end
        9021: begin
            cosine_reg0 <= 36'sb100001100110101000001110001111110010;
            sine_reg0   <= 36'sb110101111111110100010100011101000000;
        end
        9022: begin
            cosine_reg0 <= 36'sb100001100110110111111100011011011100;
            sine_reg0   <= 36'sb110101111111000100100100110111010001;
        end
        9023: begin
            cosine_reg0 <= 36'sb100001100111000111101011110010000110;
            sine_reg0   <= 36'sb110101111110010100110101101010001111;
        end
        9024: begin
            cosine_reg0 <= 36'sb100001100111010111011100010011101111;
            sine_reg0   <= 36'sb110101111101100101000110110101111101;
        end
        9025: begin
            cosine_reg0 <= 36'sb100001100111100111001110000000010110;
            sine_reg0   <= 36'sb110101111100110101011000011010011100;
        end
        9026: begin
            cosine_reg0 <= 36'sb100001100111110111000000110111111010;
            sine_reg0   <= 36'sb110101111100000101101010010111101110;
        end
        9027: begin
            cosine_reg0 <= 36'sb100001101000000110110100111010011011;
            sine_reg0   <= 36'sb110101111011010101111100101101110101;
        end
        9028: begin
            cosine_reg0 <= 36'sb100001101000010110101010000111111001;
            sine_reg0   <= 36'sb110101111010100110001111011100110011;
        end
        9029: begin
            cosine_reg0 <= 36'sb100001101000100110100000100000010011;
            sine_reg0   <= 36'sb110101111001110110100010100100101000;
        end
        9030: begin
            cosine_reg0 <= 36'sb100001101000110110011000000011100111;
            sine_reg0   <= 36'sb110101111001000110110110000101011001;
        end
        9031: begin
            cosine_reg0 <= 36'sb100001101001000110010000110001110111;
            sine_reg0   <= 36'sb110101111000010111001001111111000101;
        end
        9032: begin
            cosine_reg0 <= 36'sb100001101001010110001010101011000000;
            sine_reg0   <= 36'sb110101110111100111011110010001101111;
        end
        9033: begin
            cosine_reg0 <= 36'sb100001101001100110000101101111000010;
            sine_reg0   <= 36'sb110101110110110111110010111101011001;
        end
        9034: begin
            cosine_reg0 <= 36'sb100001101001110110000001111101111101;
            sine_reg0   <= 36'sb110101110110001000001000000010000101;
        end
        9035: begin
            cosine_reg0 <= 36'sb100001101010000101111111010111110001;
            sine_reg0   <= 36'sb110101110101011000011101011111110100;
        end
        9036: begin
            cosine_reg0 <= 36'sb100001101010010101111101111100011011;
            sine_reg0   <= 36'sb110101110100101000110011010110101001;
        end
        9037: begin
            cosine_reg0 <= 36'sb100001101010100101111101101011111101;
            sine_reg0   <= 36'sb110101110011111001001001100110100101;
        end
        9038: begin
            cosine_reg0 <= 36'sb100001101010110101111110100110010101;
            sine_reg0   <= 36'sb110101110011001001100000001111101001;
        end
        9039: begin
            cosine_reg0 <= 36'sb100001101011000110000000101011100010;
            sine_reg0   <= 36'sb110101110010011001110111010001111001;
        end
        9040: begin
            cosine_reg0 <= 36'sb100001101011010110000011111011100100;
            sine_reg0   <= 36'sb110101110001101010001110101101010101;
        end
        9041: begin
            cosine_reg0 <= 36'sb100001101011100110001000010110011011;
            sine_reg0   <= 36'sb110101110000111010100110100010000000;
        end
        9042: begin
            cosine_reg0 <= 36'sb100001101011110110001101111100000110;
            sine_reg0   <= 36'sb110101110000001010111110101111111011;
        end
        9043: begin
            cosine_reg0 <= 36'sb100001101100000110010100101100100011;
            sine_reg0   <= 36'sb110101101111011011010111010111001001;
        end
        9044: begin
            cosine_reg0 <= 36'sb100001101100010110011100100111110011;
            sine_reg0   <= 36'sb110101101110101011110000010111101010;
        end
        9045: begin
            cosine_reg0 <= 36'sb100001101100100110100101101101110101;
            sine_reg0   <= 36'sb110101101101111100001001110001100010;
        end
        9046: begin
            cosine_reg0 <= 36'sb100001101100110110101111111110101001;
            sine_reg0   <= 36'sb110101101101001100100011100100110001;
        end
        9047: begin
            cosine_reg0 <= 36'sb100001101101000110111011011010001101;
            sine_reg0   <= 36'sb110101101100011100111101110001011001;
        end
        9048: begin
            cosine_reg0 <= 36'sb100001101101010111001000000000100000;
            sine_reg0   <= 36'sb110101101011101101011000010111011101;
        end
        9049: begin
            cosine_reg0 <= 36'sb100001101101100111010101110001100100;
            sine_reg0   <= 36'sb110101101010111101110011010110111110;
        end
        9050: begin
            cosine_reg0 <= 36'sb100001101101110111100100101101010110;
            sine_reg0   <= 36'sb110101101010001110001110101111111110;
        end
        9051: begin
            cosine_reg0 <= 36'sb100001101110000111110100110011110110;
            sine_reg0   <= 36'sb110101101001011110101010100010011111;
        end
        9052: begin
            cosine_reg0 <= 36'sb100001101110011000000110000101000100;
            sine_reg0   <= 36'sb110101101000101111000110101110100011;
        end
        9053: begin
            cosine_reg0 <= 36'sb100001101110101000011000100000111111;
            sine_reg0   <= 36'sb110101100111111111100011010100001011;
        end
        9054: begin
            cosine_reg0 <= 36'sb100001101110111000101100000111100110;
            sine_reg0   <= 36'sb110101100111010000000000010011011010;
        end
        9055: begin
            cosine_reg0 <= 36'sb100001101111001001000000111000111000;
            sine_reg0   <= 36'sb110101100110100000011101101100010000;
        end
        9056: begin
            cosine_reg0 <= 36'sb100001101111011001010110110100110110;
            sine_reg0   <= 36'sb110101100101110000111011011110110001;
        end
        9057: begin
            cosine_reg0 <= 36'sb100001101111101001101101111011011110;
            sine_reg0   <= 36'sb110101100101000001011001101010111110;
        end
        9058: begin
            cosine_reg0 <= 36'sb100001101111111010000110001100110000;
            sine_reg0   <= 36'sb110101100100010001111000010000111000;
        end
        9059: begin
            cosine_reg0 <= 36'sb100001110000001010011111101000101011;
            sine_reg0   <= 36'sb110101100011100010010111010000100010;
        end
        9060: begin
            cosine_reg0 <= 36'sb100001110000011010111010001111001110;
            sine_reg0   <= 36'sb110101100010110010110110101001111110;
        end
        9061: begin
            cosine_reg0 <= 36'sb100001110000101011010110000000011001;
            sine_reg0   <= 36'sb110101100010000011010110011101001100;
        end
        9062: begin
            cosine_reg0 <= 36'sb100001110000111011110010111100001100;
            sine_reg0   <= 36'sb110101100001010011110110101010010000;
        end
        9063: begin
            cosine_reg0 <= 36'sb100001110001001100010001000010100101;
            sine_reg0   <= 36'sb110101100000100100010111010001001010;
        end
        9064: begin
            cosine_reg0 <= 36'sb100001110001011100110000010011100011;
            sine_reg0   <= 36'sb110101011111110100111000010001111101;
        end
        9065: begin
            cosine_reg0 <= 36'sb100001110001101101010000101111001000;
            sine_reg0   <= 36'sb110101011111000101011001101100101011;
        end
        9066: begin
            cosine_reg0 <= 36'sb100001110001111101110010010101010001;
            sine_reg0   <= 36'sb110101011110010101111011100001010101;
        end
        9067: begin
            cosine_reg0 <= 36'sb100001110010001110010101000101111110;
            sine_reg0   <= 36'sb110101011101100110011101101111111101;
        end
        9068: begin
            cosine_reg0 <= 36'sb100001110010011110111001000001001110;
            sine_reg0   <= 36'sb110101011100110111000000011000100101;
        end
        9069: begin
            cosine_reg0 <= 36'sb100001110010101111011110000111000001;
            sine_reg0   <= 36'sb110101011100000111100011011011001111;
        end
        9070: begin
            cosine_reg0 <= 36'sb100001110011000000000100010111010110;
            sine_reg0   <= 36'sb110101011011011000000110110111111101;
        end
        9071: begin
            cosine_reg0 <= 36'sb100001110011010000101011110010001101;
            sine_reg0   <= 36'sb110101011010101000101010101110110000;
        end
        9072: begin
            cosine_reg0 <= 36'sb100001110011100001010100010111100101;
            sine_reg0   <= 36'sb110101011001111001001110111111101010;
        end
        9073: begin
            cosine_reg0 <= 36'sb100001110011110001111110000111011101;
            sine_reg0   <= 36'sb110101011001001001110011101010101110;
        end
        9074: begin
            cosine_reg0 <= 36'sb100001110100000010101001000001110100;
            sine_reg0   <= 36'sb110101011000011010011000101111111101;
        end
        9075: begin
            cosine_reg0 <= 36'sb100001110100010011010101000110101010;
            sine_reg0   <= 36'sb110101010111101010111110001111011000;
        end
        9076: begin
            cosine_reg0 <= 36'sb100001110100100100000010010101111111;
            sine_reg0   <= 36'sb110101010110111011100100001001000010;
        end
        9077: begin
            cosine_reg0 <= 36'sb100001110100110100110000101111110001;
            sine_reg0   <= 36'sb110101010110001100001010011100111101;
        end
        9078: begin
            cosine_reg0 <= 36'sb100001110101000101100000010100000000;
            sine_reg0   <= 36'sb110101010101011100110001001011001010;
        end
        9079: begin
            cosine_reg0 <= 36'sb100001110101010110010001000010101011;
            sine_reg0   <= 36'sb110101010100101101011000010011101011;
        end
        9080: begin
            cosine_reg0 <= 36'sb100001110101100111000010111011110011;
            sine_reg0   <= 36'sb110101010011111101111111110110100010;
        end
        9081: begin
            cosine_reg0 <= 36'sb100001110101110111110101111111010101;
            sine_reg0   <= 36'sb110101010011001110100111110011110001;
        end
        9082: begin
            cosine_reg0 <= 36'sb100001110110001000101010001101010010;
            sine_reg0   <= 36'sb110101010010011111010000001011011001;
        end
        9083: begin
            cosine_reg0 <= 36'sb100001110110011001011111100101101000;
            sine_reg0   <= 36'sb110101010001101111111000111101011101;
        end
        9084: begin
            cosine_reg0 <= 36'sb100001110110101010010110001000010111;
            sine_reg0   <= 36'sb110101010001000000100010001001111110;
        end
        9085: begin
            cosine_reg0 <= 36'sb100001110110111011001101110101011111;
            sine_reg0   <= 36'sb110101010000010001001011110000111110;
        end
        9086: begin
            cosine_reg0 <= 36'sb100001110111001100000110101100111111;
            sine_reg0   <= 36'sb110101001111100001110101110010011111;
        end
        9087: begin
            cosine_reg0 <= 36'sb100001110111011101000000101110110110;
            sine_reg0   <= 36'sb110101001110110010100000001110100011;
        end
        9088: begin
            cosine_reg0 <= 36'sb100001110111101101111011111011000011;
            sine_reg0   <= 36'sb110101001110000011001011000101001011;
        end
        9089: begin
            cosine_reg0 <= 36'sb100001110111111110111000010001100111;
            sine_reg0   <= 36'sb110101001101010011110110010110011010;
        end
        9090: begin
            cosine_reg0 <= 36'sb100001111000001111110101110010011111;
            sine_reg0   <= 36'sb110101001100100100100010000010010001;
        end
        9091: begin
            cosine_reg0 <= 36'sb100001111000100000110100011101101100;
            sine_reg0   <= 36'sb110101001011110101001110001000110010;
        end
        9092: begin
            cosine_reg0 <= 36'sb100001111000110001110100010011001101;
            sine_reg0   <= 36'sb110101001011000101111010101001111110;
        end
        9093: begin
            cosine_reg0 <= 36'sb100001111001000010110101010011000001;
            sine_reg0   <= 36'sb110101001010010110100111100101111001;
        end
        9094: begin
            cosine_reg0 <= 36'sb100001111001010011110111011101000111;
            sine_reg0   <= 36'sb110101001001100111010100111100100011;
        end
        9095: begin
            cosine_reg0 <= 36'sb100001111001100100111010110001100000;
            sine_reg0   <= 36'sb110101001000111000000010101101111110;
        end
        9096: begin
            cosine_reg0 <= 36'sb100001111001110101111111010000001010;
            sine_reg0   <= 36'sb110101001000001000110000111010001101;
        end
        9097: begin
            cosine_reg0 <= 36'sb100001111010000111000100111001000100;
            sine_reg0   <= 36'sb110101000111011001011111100001010000;
        end
        9098: begin
            cosine_reg0 <= 36'sb100001111010011000001011101100001111;
            sine_reg0   <= 36'sb110101000110101010001110100011001010;
        end
        9099: begin
            cosine_reg0 <= 36'sb100001111010101001010011101001101000;
            sine_reg0   <= 36'sb110101000101111010111101111111111101;
        end
        9100: begin
            cosine_reg0 <= 36'sb100001111010111010011100110001010001;
            sine_reg0   <= 36'sb110101000101001011101101110111101010;
        end
        9101: begin
            cosine_reg0 <= 36'sb100001111011001011100111000011000111;
            sine_reg0   <= 36'sb110101000100011100011110001010010100;
        end
        9102: begin
            cosine_reg0 <= 36'sb100001111011011100110010011111001010;
            sine_reg0   <= 36'sb110101000011101101001110110111111100;
        end
        9103: begin
            cosine_reg0 <= 36'sb100001111011101101111111000101011010;
            sine_reg0   <= 36'sb110101000010111110000000000000100011;
        end
        9104: begin
            cosine_reg0 <= 36'sb100001111011111111001100110101110111;
            sine_reg0   <= 36'sb110101000010001110110001100100001101;
        end
        9105: begin
            cosine_reg0 <= 36'sb100001111100010000011011110000011110;
            sine_reg0   <= 36'sb110101000001011111100011100010111001;
        end
        9106: begin
            cosine_reg0 <= 36'sb100001111100100001101011110101010000;
            sine_reg0   <= 36'sb110101000000110000010101111100101100;
        end
        9107: begin
            cosine_reg0 <= 36'sb100001111100110010111101000100001100;
            sine_reg0   <= 36'sb110101000000000001001000110001100101;
        end
        9108: begin
            cosine_reg0 <= 36'sb100001111101000100001111011101010010;
            sine_reg0   <= 36'sb110100111111010001111100000001100111;
        end
        9109: begin
            cosine_reg0 <= 36'sb100001111101010101100011000000100000;
            sine_reg0   <= 36'sb110100111110100010101111101100110100;
        end
        9110: begin
            cosine_reg0 <= 36'sb100001111101100110110111101101110110;
            sine_reg0   <= 36'sb110100111101110011100011110011001110;
        end
        9111: begin
            cosine_reg0 <= 36'sb100001111101111000001101100101010011;
            sine_reg0   <= 36'sb110100111101000100011000010100110111;
        end
        9112: begin
            cosine_reg0 <= 36'sb100001111110001001100100100110110111;
            sine_reg0   <= 36'sb110100111100010101001101010001101111;
        end
        9113: begin
            cosine_reg0 <= 36'sb100001111110011010111100110010100001;
            sine_reg0   <= 36'sb110100111011100110000010101001111010;
        end
        9114: begin
            cosine_reg0 <= 36'sb100001111110101100010110001000010000;
            sine_reg0   <= 36'sb110100111010110110111000011101011001;
        end
        9115: begin
            cosine_reg0 <= 36'sb100001111110111101110000101000000100;
            sine_reg0   <= 36'sb110100111010000111101110101100001101;
        end
        9116: begin
            cosine_reg0 <= 36'sb100001111111001111001100010001111100;
            sine_reg0   <= 36'sb110100111001011000100101010110011001;
        end
        9117: begin
            cosine_reg0 <= 36'sb100001111111100000101001000101110111;
            sine_reg0   <= 36'sb110100111000101001011100011011111110;
        end
        9118: begin
            cosine_reg0 <= 36'sb100001111111110010000111000011110101;
            sine_reg0   <= 36'sb110100110111111010010011111100111111;
        end
        9119: begin
            cosine_reg0 <= 36'sb100010000000000011100110001011110101;
            sine_reg0   <= 36'sb110100110111001011001011111001011100;
        end
        9120: begin
            cosine_reg0 <= 36'sb100010000000010101000110011101110110;
            sine_reg0   <= 36'sb110100110110011100000100010001011000;
        end
        9121: begin
            cosine_reg0 <= 36'sb100010000000100110100111111001110111;
            sine_reg0   <= 36'sb110100110101101100111101000100110101;
        end
        9122: begin
            cosine_reg0 <= 36'sb100010000000111000001010011111111001;
            sine_reg0   <= 36'sb110100110100111101110110010011110101;
        end
        9123: begin
            cosine_reg0 <= 36'sb100010000001001001101110001111111001;
            sine_reg0   <= 36'sb110100110100001110101111111110011001;
        end
        9124: begin
            cosine_reg0 <= 36'sb100010000001011011010011001001111001;
            sine_reg0   <= 36'sb110100110011011111101010000100100010;
        end
        9125: begin
            cosine_reg0 <= 36'sb100010000001101100111001001101110110;
            sine_reg0   <= 36'sb110100110010110000100100100110010100;
        end
        9126: begin
            cosine_reg0 <= 36'sb100010000001111110100000011011110000;
            sine_reg0   <= 36'sb110100110010000001011111100011101111;
        end
        9127: begin
            cosine_reg0 <= 36'sb100010000010010000001000110011100111;
            sine_reg0   <= 36'sb110100110001010010011010111100110110;
        end
        9128: begin
            cosine_reg0 <= 36'sb100010000010100001110010010101011010;
            sine_reg0   <= 36'sb110100110000100011010110110001101011;
        end
        9129: begin
            cosine_reg0 <= 36'sb100010000010110011011101000001001000;
            sine_reg0   <= 36'sb110100101111110100010011000010001110;
        end
        9130: begin
            cosine_reg0 <= 36'sb100010000011000101001000110110110000;
            sine_reg0   <= 36'sb110100101111000101001111101110100011;
        end
        9131: begin
            cosine_reg0 <= 36'sb100010000011010110110101110110010011;
            sine_reg0   <= 36'sb110100101110010110001100110110101010;
        end
        9132: begin
            cosine_reg0 <= 36'sb100010000011101000100011111111101110;
            sine_reg0   <= 36'sb110100101101100111001010011010100110;
        end
        9133: begin
            cosine_reg0 <= 36'sb100010000011111010010011010011000010;
            sine_reg0   <= 36'sb110100101100111000001000011010011000;
        end
        9134: begin
            cosine_reg0 <= 36'sb100010000100001100000011110000001110;
            sine_reg0   <= 36'sb110100101100001001000110110110000010;
        end
        9135: begin
            cosine_reg0 <= 36'sb100010000100011101110101010111010000;
            sine_reg0   <= 36'sb110100101011011010000101101101100111;
        end
        9136: begin
            cosine_reg0 <= 36'sb100010000100101111101000001000001001;
            sine_reg0   <= 36'sb110100101010101011000101000001000111;
        end
        9137: begin
            cosine_reg0 <= 36'sb100010000101000001011100000010111000;
            sine_reg0   <= 36'sb110100101001111100000100110000100110;
        end
        9138: begin
            cosine_reg0 <= 36'sb100010000101010011010001000111011100;
            sine_reg0   <= 36'sb110100101001001101000100111100000011;
        end
        9139: begin
            cosine_reg0 <= 36'sb100010000101100101000111010101110100;
            sine_reg0   <= 36'sb110100101000011110000101100011100010;
        end
        9140: begin
            cosine_reg0 <= 36'sb100010000101110110111110101110000000;
            sine_reg0   <= 36'sb110100100111101111000110100111000100;
        end
        9141: begin
            cosine_reg0 <= 36'sb100010000110001000110111001111111111;
            sine_reg0   <= 36'sb110100100111000000001000000110101011;
        end
        9142: begin
            cosine_reg0 <= 36'sb100010000110011010110000111011110000;
            sine_reg0   <= 36'sb110100100110010001001010000010011000;
        end
        9143: begin
            cosine_reg0 <= 36'sb100010000110101100101011110001010010;
            sine_reg0   <= 36'sb110100100101100010001100011010001111;
        end
        9144: begin
            cosine_reg0 <= 36'sb100010000110111110100111110000100110;
            sine_reg0   <= 36'sb110100100100110011001111001110001111;
        end
        9145: begin
            cosine_reg0 <= 36'sb100010000111010000100100111001101001;
            sine_reg0   <= 36'sb110100100100000100010010011110011100;
        end
        9146: begin
            cosine_reg0 <= 36'sb100010000111100010100011001100011100;
            sine_reg0   <= 36'sb110100100011010101010110001010110110;
        end
        9147: begin
            cosine_reg0 <= 36'sb100010000111110100100010101000111110;
            sine_reg0   <= 36'sb110100100010100110011010010011100001;
        end
        9148: begin
            cosine_reg0 <= 36'sb100010001000000110100011001111001110;
            sine_reg0   <= 36'sb110100100001110111011110111000011101;
        end
        9149: begin
            cosine_reg0 <= 36'sb100010001000011000100100111111001100;
            sine_reg0   <= 36'sb110100100001001000100011111001101100;
        end
        9150: begin
            cosine_reg0 <= 36'sb100010001000101010100111111000110110;
            sine_reg0   <= 36'sb110100100000011001101001010111010001;
        end
        9151: begin
            cosine_reg0 <= 36'sb100010001000111100101011111100001100;
            sine_reg0   <= 36'sb110100011111101010101111010001001101;
        end
        9152: begin
            cosine_reg0 <= 36'sb100010001001001110110001001001001110;
            sine_reg0   <= 36'sb110100011110111011110101100111100001;
        end
        9153: begin
            cosine_reg0 <= 36'sb100010001001100000110111011111111010;
            sine_reg0   <= 36'sb110100011110001100111100011010010000;
        end
        9154: begin
            cosine_reg0 <= 36'sb100010001001110010111111000000010000;
            sine_reg0   <= 36'sb110100011101011110000011101001011100;
        end
        9155: begin
            cosine_reg0 <= 36'sb100010001010000101000111101010001111;
            sine_reg0   <= 36'sb110100011100101111001011010101000110;
        end
        9156: begin
            cosine_reg0 <= 36'sb100010001010010111010001011101110111;
            sine_reg0   <= 36'sb110100011100000000010011011101001111;
        end
        9157: begin
            cosine_reg0 <= 36'sb100010001010101001011100011011000111;
            sine_reg0   <= 36'sb110100011011010001011100000001111011;
        end
        9158: begin
            cosine_reg0 <= 36'sb100010001010111011101000100001111110;
            sine_reg0   <= 36'sb110100011010100010100101000011001011;
        end
        9159: begin
            cosine_reg0 <= 36'sb100010001011001101110101110010011011;
            sine_reg0   <= 36'sb110100011001110011101110100000111111;
        end
        9160: begin
            cosine_reg0 <= 36'sb100010001011100000000100001100011110;
            sine_reg0   <= 36'sb110100011001000100111000011011011100;
        end
        9161: begin
            cosine_reg0 <= 36'sb100010001011110010010011110000000110;
            sine_reg0   <= 36'sb110100011000010110000010110010100001;
        end
        9162: begin
            cosine_reg0 <= 36'sb100010001100000100100100011101010011;
            sine_reg0   <= 36'sb110100010111100111001101100110010001;
        end
        9163: begin
            cosine_reg0 <= 36'sb100010001100010110110110010100000011;
            sine_reg0   <= 36'sb110100010110111000011000110110101110;
        end
        9164: begin
            cosine_reg0 <= 36'sb100010001100101001001001010100010110;
            sine_reg0   <= 36'sb110100010110001001100100100011111001;
        end
        9165: begin
            cosine_reg0 <= 36'sb100010001100111011011101011110001011;
            sine_reg0   <= 36'sb110100010101011010110000101101110101;
        end
        9166: begin
            cosine_reg0 <= 36'sb100010001101001101110010110001100010;
            sine_reg0   <= 36'sb110100010100101011111101010100100011;
        end
        9167: begin
            cosine_reg0 <= 36'sb100010001101100000001001001110011001;
            sine_reg0   <= 36'sb110100010011111101001010011000000100;
        end
        9168: begin
            cosine_reg0 <= 36'sb100010001101110010100000110100110001;
            sine_reg0   <= 36'sb110100010011001110010111111000011100;
        end
        9169: begin
            cosine_reg0 <= 36'sb100010001110000100111001100100101000;
            sine_reg0   <= 36'sb110100010010011111100101110101101011;
        end
        9170: begin
            cosine_reg0 <= 36'sb100010001110010111010011011101111101;
            sine_reg0   <= 36'sb110100010001110000110100001111110011;
        end
        9171: begin
            cosine_reg0 <= 36'sb100010001110101001101110100000110001;
            sine_reg0   <= 36'sb110100010001000010000011000110110111;
        end
        9172: begin
            cosine_reg0 <= 36'sb100010001110111100001010101101000010;
            sine_reg0   <= 36'sb110100010000010011010010011010110111;
        end
        9173: begin
            cosine_reg0 <= 36'sb100010001111001110101000000010101111;
            sine_reg0   <= 36'sb110100001111100100100010001011110110;
        end
        9174: begin
            cosine_reg0 <= 36'sb100010001111100001000110100001111000;
            sine_reg0   <= 36'sb110100001110110101110010011001110110;
        end
        9175: begin
            cosine_reg0 <= 36'sb100010001111110011100110001010011101;
            sine_reg0   <= 36'sb110100001110000111000011000100111000;
        end
        9176: begin
            cosine_reg0 <= 36'sb100010010000000110000110111100011100;
            sine_reg0   <= 36'sb110100001101011000010100001100111110;
        end
        9177: begin
            cosine_reg0 <= 36'sb100010010000011000101000110111110100;
            sine_reg0   <= 36'sb110100001100101001100101110010001010;
        end
        9178: begin
            cosine_reg0 <= 36'sb100010010000101011001011111100100101;
            sine_reg0   <= 36'sb110100001011111010110111110100011110;
        end
        9179: begin
            cosine_reg0 <= 36'sb100010010000111101110000001010101111;
            sine_reg0   <= 36'sb110100001011001100001010010011111011;
        end
        9180: begin
            cosine_reg0 <= 36'sb100010010001010000010101100010010000;
            sine_reg0   <= 36'sb110100001010011101011101010000100100;
        end
        9181: begin
            cosine_reg0 <= 36'sb100010010001100010111100000011001001;
            sine_reg0   <= 36'sb110100001001101110110000101010011010;
        end
        9182: begin
            cosine_reg0 <= 36'sb100010010001110101100011101101010111;
            sine_reg0   <= 36'sb110100001001000000000100100001011111;
        end
        9183: begin
            cosine_reg0 <= 36'sb100010010010001000001100100000111010;
            sine_reg0   <= 36'sb110100001000010001011000110101110100;
        end
        9184: begin
            cosine_reg0 <= 36'sb100010010010011010110110011101110011;
            sine_reg0   <= 36'sb110100000111100010101101100111011101;
        end
        9185: begin
            cosine_reg0 <= 36'sb100010010010101101100001100011111111;
            sine_reg0   <= 36'sb110100000110110100000010110110011001;
        end
        9186: begin
            cosine_reg0 <= 36'sb100010010011000000001101110011011111;
            sine_reg0   <= 36'sb110100000110000101011000100010101100;
        end
        9187: begin
            cosine_reg0 <= 36'sb100010010011010010111011001100010001;
            sine_reg0   <= 36'sb110100000101010110101110101100010111;
        end
        9188: begin
            cosine_reg0 <= 36'sb100010010011100101101001101110010100;
            sine_reg0   <= 36'sb110100000100101000000101010011011011;
        end
        9189: begin
            cosine_reg0 <= 36'sb100010010011111000011001011001101001;
            sine_reg0   <= 36'sb110100000011111001011100010111111011;
        end
        9190: begin
            cosine_reg0 <= 36'sb100010010100001011001010001110001111;
            sine_reg0   <= 36'sb110100000011001010110011111001111000;
        end
        9191: begin
            cosine_reg0 <= 36'sb100010010100011101111100001100000011;
            sine_reg0   <= 36'sb110100000010011100001011111001010101;
        end
        9192: begin
            cosine_reg0 <= 36'sb100010010100110000101111010011000111;
            sine_reg0   <= 36'sb110100000001101101100100010110010010;
        end
        9193: begin
            cosine_reg0 <= 36'sb100010010101000011100011100011011001;
            sine_reg0   <= 36'sb110100000000111110111101010000110010;
        end
        9194: begin
            cosine_reg0 <= 36'sb100010010101010110011000111100111001;
            sine_reg0   <= 36'sb110100000000010000010110101000110111;
        end
        9195: begin
            cosine_reg0 <= 36'sb100010010101101001001111011111100101;
            sine_reg0   <= 36'sb110011111111100001110000011110100010;
        end
        9196: begin
            cosine_reg0 <= 36'sb100010010101111100000111001011011101;
            sine_reg0   <= 36'sb110011111110110011001010110001110101;
        end
        9197: begin
            cosine_reg0 <= 36'sb100010010110001111000000000000100001;
            sine_reg0   <= 36'sb110011111110000100100101100010110010;
        end
        9198: begin
            cosine_reg0 <= 36'sb100010010110100001111001111110101111;
            sine_reg0   <= 36'sb110011111101010110000000110001011011;
        end
        9199: begin
            cosine_reg0 <= 36'sb100010010110110100110101000110000110;
            sine_reg0   <= 36'sb110011111100100111011100011101110001;
        end
        9200: begin
            cosine_reg0 <= 36'sb100010010111000111110001010110100111;
            sine_reg0   <= 36'sb110011111011111000111000100111110111;
        end
        9201: begin
            cosine_reg0 <= 36'sb100010010111011010101110110000010001;
            sine_reg0   <= 36'sb110011111011001010010101001111101101;
        end
        9202: begin
            cosine_reg0 <= 36'sb100010010111101101101101010011000001;
            sine_reg0   <= 36'sb110011111010011011110010010101010111;
        end
        9203: begin
            cosine_reg0 <= 36'sb100010011000000000101100111110111001;
            sine_reg0   <= 36'sb110011111001101101001111111000110101;
        end
        9204: begin
            cosine_reg0 <= 36'sb100010011000010011101101110011110111;
            sine_reg0   <= 36'sb110011111000111110101101111010001010;
        end
        9205: begin
            cosine_reg0 <= 36'sb100010011000100110101111110001111011;
            sine_reg0   <= 36'sb110011111000010000001100011001010111;
        end
        9206: begin
            cosine_reg0 <= 36'sb100010011000111001110010111001000011;
            sine_reg0   <= 36'sb110011110111100001101011010110011110;
        end
        9207: begin
            cosine_reg0 <= 36'sb100010011001001100110111001001001111;
            sine_reg0   <= 36'sb110011110110110011001010110001100001;
        end
        9208: begin
            cosine_reg0 <= 36'sb100010011001011111111100100010011110;
            sine_reg0   <= 36'sb110011110110000100101010101010100010;
        end
        9209: begin
            cosine_reg0 <= 36'sb100010011001110011000011000100110000;
            sine_reg0   <= 36'sb110011110101010110001011000001100010;
        end
        9210: begin
            cosine_reg0 <= 36'sb100010011010000110001010110000000011;
            sine_reg0   <= 36'sb110011110100100111101011110110100011;
        end
        9211: begin
            cosine_reg0 <= 36'sb100010011010011001010011100100011000;
            sine_reg0   <= 36'sb110011110011111001001101001001101000;
        end
        9212: begin
            cosine_reg0 <= 36'sb100010011010101100011101100001101101;
            sine_reg0   <= 36'sb110011110011001010101110111010110001;
        end
        9213: begin
            cosine_reg0 <= 36'sb100010011010111111101000101000000001;
            sine_reg0   <= 36'sb110011110010011100010001001010000001;
        end
        9214: begin
            cosine_reg0 <= 36'sb100010011011010010110100110111010100;
            sine_reg0   <= 36'sb110011110001101101110011110111011001;
        end
        9215: begin
            cosine_reg0 <= 36'sb100010011011100110000010001111100110;
            sine_reg0   <= 36'sb110011110000111111010111000010111100;
        end
        9216: begin
            cosine_reg0 <= 36'sb100010011011111001010000110000110100;
            sine_reg0   <= 36'sb110011110000010000111010101100101011;
        end
        9217: begin
            cosine_reg0 <= 36'sb100010011100001100100000011010111111;
            sine_reg0   <= 36'sb110011101111100010011110110100100111;
        end
        9218: begin
            cosine_reg0 <= 36'sb100010011100011111110001001110000110;
            sine_reg0   <= 36'sb110011101110110100000011011010110011;
        end
        9219: begin
            cosine_reg0 <= 36'sb100010011100110011000011001010001001;
            sine_reg0   <= 36'sb110011101110000101101000011111010000;
        end
        9220: begin
            cosine_reg0 <= 36'sb100010011101000110010110001111000101;
            sine_reg0   <= 36'sb110011101101010111001110000010000001;
        end
        9221: begin
            cosine_reg0 <= 36'sb100010011101011001101010011100111011;
            sine_reg0   <= 36'sb110011101100101000110100000011000110;
        end
        9222: begin
            cosine_reg0 <= 36'sb100010011101101100111111110011101010;
            sine_reg0   <= 36'sb110011101011111010011010100010100010;
        end
        9223: begin
            cosine_reg0 <= 36'sb100010011110000000010110010011010001;
            sine_reg0   <= 36'sb110011101011001100000001100000010111;
        end
        9224: begin
            cosine_reg0 <= 36'sb100010011110010011101101111011110000;
            sine_reg0   <= 36'sb110011101010011101101000111100100110;
        end
        9225: begin
            cosine_reg0 <= 36'sb100010011110100111000110101101000101;
            sine_reg0   <= 36'sb110011101001101111010000110111010001;
        end
        9226: begin
            cosine_reg0 <= 36'sb100010011110111010100000100111010000;
            sine_reg0   <= 36'sb110011101001000000111001010000011010;
        end
        9227: begin
            cosine_reg0 <= 36'sb100010011111001101111011101010010000;
            sine_reg0   <= 36'sb110011101000010010100010001000000010;
        end
        9228: begin
            cosine_reg0 <= 36'sb100010011111100001010111110110000100;
            sine_reg0   <= 36'sb110011100111100100001011011110001100;
        end
        9229: begin
            cosine_reg0 <= 36'sb100010011111110100110101001010101100;
            sine_reg0   <= 36'sb110011100110110101110101010010111010;
        end
        9230: begin
            cosine_reg0 <= 36'sb100010100000001000010011101000000111;
            sine_reg0   <= 36'sb110011100110000111011111100110001100;
        end
        9231: begin
            cosine_reg0 <= 36'sb100010100000011011110011001110010100;
            sine_reg0   <= 36'sb110011100101011001001010011000000101;
        end
        9232: begin
            cosine_reg0 <= 36'sb100010100000101111010011111101010011;
            sine_reg0   <= 36'sb110011100100101010110101101000100111;
        end
        9233: begin
            cosine_reg0 <= 36'sb100010100001000010110101110101000010;
            sine_reg0   <= 36'sb110011100011111100100001010111110100;
        end
        9234: begin
            cosine_reg0 <= 36'sb100010100001010110011000110101100001;
            sine_reg0   <= 36'sb110011100011001110001101100101101100;
        end
        9235: begin
            cosine_reg0 <= 36'sb100010100001101001111100111110101111;
            sine_reg0   <= 36'sb110011100010011111111010010010010010;
        end
        9236: begin
            cosine_reg0 <= 36'sb100010100001111101100010010000101011;
            sine_reg0   <= 36'sb110011100001110001100111011101101001;
        end
        9237: begin
            cosine_reg0 <= 36'sb100010100010010001001000101011010101;
            sine_reg0   <= 36'sb110011100001000011010101000111110000;
        end
        9238: begin
            cosine_reg0 <= 36'sb100010100010100100110000001110101100;
            sine_reg0   <= 36'sb110011100000010101000011010000101011;
        end
        9239: begin
            cosine_reg0 <= 36'sb100010100010111000011000111010110000;
            sine_reg0   <= 36'sb110011011111100110110001111000011011;
        end
        9240: begin
            cosine_reg0 <= 36'sb100010100011001100000010101111011110;
            sine_reg0   <= 36'sb110011011110111000100000111111000010;
        end
        9241: begin
            cosine_reg0 <= 36'sb100010100011011111101101101100110111;
            sine_reg0   <= 36'sb110011011110001010010000100100100010;
        end
        9242: begin
            cosine_reg0 <= 36'sb100010100011110011011001110010111010;
            sine_reg0   <= 36'sb110011011101011100000000101000111100;
        end
        9243: begin
            cosine_reg0 <= 36'sb100010100100000111000111000001100110;
            sine_reg0   <= 36'sb110011011100101101110001001100010011;
        end
        9244: begin
            cosine_reg0 <= 36'sb100010100100011010110101011000111010;
            sine_reg0   <= 36'sb110011011011111111100010001110100111;
        end
        9245: begin
            cosine_reg0 <= 36'sb100010100100101110100100111000110110;
            sine_reg0   <= 36'sb110011011011010001010011101111111011;
        end
        9246: begin
            cosine_reg0 <= 36'sb100010100101000010010101100001011000;
            sine_reg0   <= 36'sb110011011010100011000101110000010001;
        end
        9247: begin
            cosine_reg0 <= 36'sb100010100101010110000111010010100001;
            sine_reg0   <= 36'sb110011011001110100111000001111101010;
        end
        9248: begin
            cosine_reg0 <= 36'sb100010100101101001111010001100001110;
            sine_reg0   <= 36'sb110011011001000110101011001110001001;
        end
        9249: begin
            cosine_reg0 <= 36'sb100010100101111101101110001110100001;
            sine_reg0   <= 36'sb110011011000011000011110101011101110;
        end
        9250: begin
            cosine_reg0 <= 36'sb100010100110010001100011011001010111;
            sine_reg0   <= 36'sb110011010111101010010010101000011100;
        end
        9251: begin
            cosine_reg0 <= 36'sb100010100110100101011001101100110000;
            sine_reg0   <= 36'sb110011010110111100000111000100010101;
        end
        9252: begin
            cosine_reg0 <= 36'sb100010100110111001010001001000101011;
            sine_reg0   <= 36'sb110011010110001101111011111111011001;
        end
        9253: begin
            cosine_reg0 <= 36'sb100010100111001101001001101101001000;
            sine_reg0   <= 36'sb110011010101011111110001011001101100;
        end
        9254: begin
            cosine_reg0 <= 36'sb100010100111100001000011011010000101;
            sine_reg0   <= 36'sb110011010100110001100111010011001111;
        end
        9255: begin
            cosine_reg0 <= 36'sb100010100111110100111110001111100010;
            sine_reg0   <= 36'sb110011010100000011011101101100000011;
        end
        9256: begin
            cosine_reg0 <= 36'sb100010101000001000111010001101011111;
            sine_reg0   <= 36'sb110011010011010101010100100100001011;
        end
        9257: begin
            cosine_reg0 <= 36'sb100010101000011100110111010011111010;
            sine_reg0   <= 36'sb110011010010100111001011111011101000;
        end
        9258: begin
            cosine_reg0 <= 36'sb100010101000110000110101100010110010;
            sine_reg0   <= 36'sb110011010001111001000011110010011100;
        end
        9259: begin
            cosine_reg0 <= 36'sb100010101001000100110100111010000111;
            sine_reg0   <= 36'sb110011010001001010111100001000101000;
        end
        9260: begin
            cosine_reg0 <= 36'sb100010101001011000110101011001111000;
            sine_reg0   <= 36'sb110011010000011100110100111110001111;
        end
        9261: begin
            cosine_reg0 <= 36'sb100010101001101100110111000010000101;
            sine_reg0   <= 36'sb110011001111101110101110010011010011;
        end
        9262: begin
            cosine_reg0 <= 36'sb100010101010000000111001110010101100;
            sine_reg0   <= 36'sb110011001111000000101000000111110100;
        end
        9263: begin
            cosine_reg0 <= 36'sb100010101010010100111101101011101101;
            sine_reg0   <= 36'sb110011001110010010100010011011110101;
        end
        9264: begin
            cosine_reg0 <= 36'sb100010101010101001000010101101000111;
            sine_reg0   <= 36'sb110011001101100100011101001111011000;
        end
        9265: begin
            cosine_reg0 <= 36'sb100010101010111101001000110110111001;
            sine_reg0   <= 36'sb110011001100110110011000100010011110;
        end
        9266: begin
            cosine_reg0 <= 36'sb100010101011010001010000001001000010;
            sine_reg0   <= 36'sb110011001100001000010100010101001010;
        end
        9267: begin
            cosine_reg0 <= 36'sb100010101011100101011000100011100010;
            sine_reg0   <= 36'sb110011001011011010010000100111011100;
        end
        9268: begin
            cosine_reg0 <= 36'sb100010101011111001100010000110011000;
            sine_reg0   <= 36'sb110011001010101100001101011001010111;
        end
        9269: begin
            cosine_reg0 <= 36'sb100010101100001101101100110001100011;
            sine_reg0   <= 36'sb110011001001111110001010101010111101;
        end
        9270: begin
            cosine_reg0 <= 36'sb100010101100100001111000100101000010;
            sine_reg0   <= 36'sb110011001001010000001000011100001111;
        end
        9271: begin
            cosine_reg0 <= 36'sb100010101100110110000101100000110101;
            sine_reg0   <= 36'sb110011001000100010000110101101001111;
        end
        9272: begin
            cosine_reg0 <= 36'sb100010101101001010010011100100111011;
            sine_reg0   <= 36'sb110011000111110100000101011101111111;
        end
        9273: begin
            cosine_reg0 <= 36'sb100010101101011110100010110001010010;
            sine_reg0   <= 36'sb110011000111000110000100101110100000;
        end
        9274: begin
            cosine_reg0 <= 36'sb100010101101110010110011000101111011;
            sine_reg0   <= 36'sb110011000110011000000100011110110101;
        end
        9275: begin
            cosine_reg0 <= 36'sb100010101110000111000100100010110100;
            sine_reg0   <= 36'sb110011000101101010000100101110111111;
        end
        9276: begin
            cosine_reg0 <= 36'sb100010101110011011010111000111111101;
            sine_reg0   <= 36'sb110011000100111100000101011110111111;
        end
        9277: begin
            cosine_reg0 <= 36'sb100010101110101111101010110101010101;
            sine_reg0   <= 36'sb110011000100001110000110101110111001;
        end
        9278: begin
            cosine_reg0 <= 36'sb100010101111000011111111101010111011;
            sine_reg0   <= 36'sb110011000011100000001000011110101101;
        end
        9279: begin
            cosine_reg0 <= 36'sb100010101111011000010101101000101110;
            sine_reg0   <= 36'sb110011000010110010001010101110011101;
        end
        9280: begin
            cosine_reg0 <= 36'sb100010101111101100101100101110101101;
            sine_reg0   <= 36'sb110011000010000100001101011110001011;
        end
        9281: begin
            cosine_reg0 <= 36'sb100010110000000001000100111100111001;
            sine_reg0   <= 36'sb110011000001010110010000101101111001;
        end
        9282: begin
            cosine_reg0 <= 36'sb100010110000010101011110010011001111;
            sine_reg0   <= 36'sb110011000000101000010100011101101001;
        end
        9283: begin
            cosine_reg0 <= 36'sb100010110000101001111000110001101111;
            sine_reg0   <= 36'sb110010111111111010011000101101011100;
        end
        9284: begin
            cosine_reg0 <= 36'sb100010110000111110010100011000011001;
            sine_reg0   <= 36'sb110010111111001100011101011101010100;
        end
        9285: begin
            cosine_reg0 <= 36'sb100010110001010010110001000111001011;
            sine_reg0   <= 36'sb110010111110011110100010101101010010;
        end
        9286: begin
            cosine_reg0 <= 36'sb100010110001100111001110111110000110;
            sine_reg0   <= 36'sb110010111101110000101000011101011010;
        end
        9287: begin
            cosine_reg0 <= 36'sb100010110001111011101101111101000111;
            sine_reg0   <= 36'sb110010111101000010101110101101101100;
        end
        9288: begin
            cosine_reg0 <= 36'sb100010110010010000001110000100001110;
            sine_reg0   <= 36'sb110010111100010100110101011110001010;
        end
        9289: begin
            cosine_reg0 <= 36'sb100010110010100100101111010011011011;
            sine_reg0   <= 36'sb110010111011100110111100101110110110;
        end
        9290: begin
            cosine_reg0 <= 36'sb100010110010111001010001101010101100;
            sine_reg0   <= 36'sb110010111010111001000100011111110001;
        end
        9291: begin
            cosine_reg0 <= 36'sb100010110011001101110101001010000001;
            sine_reg0   <= 36'sb110010111010001011001100110000111111;
        end
        9292: begin
            cosine_reg0 <= 36'sb100010110011100010011001110001011001;
            sine_reg0   <= 36'sb110010111001011101010101100010011111;
        end
        9293: begin
            cosine_reg0 <= 36'sb100010110011110110111111100000110100;
            sine_reg0   <= 36'sb110010111000101111011110110100010100;
        end
        9294: begin
            cosine_reg0 <= 36'sb100010110100001011100110011000010000;
            sine_reg0   <= 36'sb110010111000000001101000100110100001;
        end
        9295: begin
            cosine_reg0 <= 36'sb100010110100100000001110010111101100;
            sine_reg0   <= 36'sb110010110111010011110010111001000101;
        end
        9296: begin
            cosine_reg0 <= 36'sb100010110100110100110111011111001001;
            sine_reg0   <= 36'sb110010110110100101111101101100000101;
        end
        9297: begin
            cosine_reg0 <= 36'sb100010110101001001100001101110100100;
            sine_reg0   <= 36'sb110010110101111000001000111111100000;
        end
        9298: begin
            cosine_reg0 <= 36'sb100010110101011110001101000101111110;
            sine_reg0   <= 36'sb110010110101001010010100110011011001;
        end
        9299: begin
            cosine_reg0 <= 36'sb100010110101110010111001100101010101;
            sine_reg0   <= 36'sb110010110100011100100001000111110001;
        end
        9300: begin
            cosine_reg0 <= 36'sb100010110110000111100111001100101001;
            sine_reg0   <= 36'sb110010110011101110101101111100101100;
        end
        9301: begin
            cosine_reg0 <= 36'sb100010110110011100010101111011111001;
            sine_reg0   <= 36'sb110010110011000000111011010010001001;
        end
        9302: begin
            cosine_reg0 <= 36'sb100010110110110001000101110011000100;
            sine_reg0   <= 36'sb110010110010010011001001001000001011;
        end
        9303: begin
            cosine_reg0 <= 36'sb100010110111000101110110110010001001;
            sine_reg0   <= 36'sb110010110001100101010111011110110100;
        end
        9304: begin
            cosine_reg0 <= 36'sb100010110111011010101000111001000111;
            sine_reg0   <= 36'sb110010110000110111100110010110000101;
        end
        9305: begin
            cosine_reg0 <= 36'sb100010110111101111011100000111111111;
            sine_reg0   <= 36'sb110010110000001001110101101110000000;
        end
        9306: begin
            cosine_reg0 <= 36'sb100010111000000100010000011110101110;
            sine_reg0   <= 36'sb110010101111011100000101100110101000;
        end
        9307: begin
            cosine_reg0 <= 36'sb100010111000011001000101111101010100;
            sine_reg0   <= 36'sb110010101110101110010101111111111101;
        end
        9308: begin
            cosine_reg0 <= 36'sb100010111000101101111100100011110001;
            sine_reg0   <= 36'sb110010101110000000100110111010000010;
        end
        9309: begin
            cosine_reg0 <= 36'sb100010111001000010110100010010000011;
            sine_reg0   <= 36'sb110010101101010010111000010100111000;
        end
        9310: begin
            cosine_reg0 <= 36'sb100010111001010111101101001000001001;
            sine_reg0   <= 36'sb110010101100100101001010010000100001;
        end
        9311: begin
            cosine_reg0 <= 36'sb100010111001101100100111000110000100;
            sine_reg0   <= 36'sb110010101011110111011100101100111110;
        end
        9312: begin
            cosine_reg0 <= 36'sb100010111010000001100010001011110001;
            sine_reg0   <= 36'sb110010101011001001101111101010010011;
        end
        9313: begin
            cosine_reg0 <= 36'sb100010111010010110011110011001010001;
            sine_reg0   <= 36'sb110010101010011100000011001000011111;
        end
        9314: begin
            cosine_reg0 <= 36'sb100010111010101011011011101110100010;
            sine_reg0   <= 36'sb110010101001101110010111000111100110;
        end
        9315: begin
            cosine_reg0 <= 36'sb100010111011000000011010001011100100;
            sine_reg0   <= 36'sb110010101001000000101011100111101001;
        end
        9316: begin
            cosine_reg0 <= 36'sb100010111011010101011001110000010110;
            sine_reg0   <= 36'sb110010101000010011000000101000101001;
        end
        9317: begin
            cosine_reg0 <= 36'sb100010111011101010011010011100110111;
            sine_reg0   <= 36'sb110010100111100101010110001010101000;
        end
        9318: begin
            cosine_reg0 <= 36'sb100010111011111111011100010001000101;
            sine_reg0   <= 36'sb110010100110110111101100001101101001;
        end
        9319: begin
            cosine_reg0 <= 36'sb100010111100010100011111001101000010;
            sine_reg0   <= 36'sb110010100110001010000010110001101101;
        end
        9320: begin
            cosine_reg0 <= 36'sb100010111100101001100011010000101010;
            sine_reg0   <= 36'sb110010100101011100011001110110110101;
        end
        9321: begin
            cosine_reg0 <= 36'sb100010111100111110101000011011111111;
            sine_reg0   <= 36'sb110010100100101110110001011101000011;
        end
        9322: begin
            cosine_reg0 <= 36'sb100010111101010011101110101110111111;
            sine_reg0   <= 36'sb110010100100000001001001100100011010;
        end
        9323: begin
            cosine_reg0 <= 36'sb100010111101101000110110001001101000;
            sine_reg0   <= 36'sb110010100011010011100010001100111011;
        end
        9324: begin
            cosine_reg0 <= 36'sb100010111101111101111110101011111011;
            sine_reg0   <= 36'sb110010100010100101111011010110100111;
        end
        9325: begin
            cosine_reg0 <= 36'sb100010111110010011001000010101110111;
            sine_reg0   <= 36'sb110010100001111000010101000001100001;
        end
        9326: begin
            cosine_reg0 <= 36'sb100010111110101000010011000111011010;
            sine_reg0   <= 36'sb110010100001001010101111001101101010;
        end
        9327: begin
            cosine_reg0 <= 36'sb100010111110111101011111000000100100;
            sine_reg0   <= 36'sb110010100000011101001001111011000100;
        end
        9328: begin
            cosine_reg0 <= 36'sb100010111111010010101100000001010100;
            sine_reg0   <= 36'sb110010011111101111100101001001110001;
        end
        9329: begin
            cosine_reg0 <= 36'sb100010111111100111111010001001101010;
            sine_reg0   <= 36'sb110010011111000010000000111001110010;
        end
        9330: begin
            cosine_reg0 <= 36'sb100010111111111101001001011001100011;
            sine_reg0   <= 36'sb110010011110010100011101001011001001;
        end
        9331: begin
            cosine_reg0 <= 36'sb100011000000010010011001110001000001;
            sine_reg0   <= 36'sb110010011101100110111001111101111000;
        end
        9332: begin
            cosine_reg0 <= 36'sb100011000000100111101011010000000001;
            sine_reg0   <= 36'sb110010011100111001010111010010000001;
        end
        9333: begin
            cosine_reg0 <= 36'sb100011000000111100111101110110100011;
            sine_reg0   <= 36'sb110010011100001011110101000111100110;
        end
        9334: begin
            cosine_reg0 <= 36'sb100011000001010010010001100100100111;
            sine_reg0   <= 36'sb110010011011011110010011011110101000;
        end
        9335: begin
            cosine_reg0 <= 36'sb100011000001100111100110011010001010;
            sine_reg0   <= 36'sb110010011010110000110010010111001000;
        end
        9336: begin
            cosine_reg0 <= 36'sb100011000001111100111100010111001101;
            sine_reg0   <= 36'sb110010011010000011010001110001001010;
        end
        9337: begin
            cosine_reg0 <= 36'sb100011000010010010010011011011101111;
            sine_reg0   <= 36'sb110010011001010101110001101100101110;
        end
        9338: begin
            cosine_reg0 <= 36'sb100011000010100111101011100111101111;
            sine_reg0   <= 36'sb110010011000101000010010001001110110;
        end
        9339: begin
            cosine_reg0 <= 36'sb100011000010111101000100111011001100;
            sine_reg0   <= 36'sb110010010111111010110011001000100101;
        end
        9340: begin
            cosine_reg0 <= 36'sb100011000011010010011111010110000100;
            sine_reg0   <= 36'sb110010010111001101010100101000111011;
        end
        9341: begin
            cosine_reg0 <= 36'sb100011000011100111111010111000011001;
            sine_reg0   <= 36'sb110010010110011111110110101010111011;
        end
        9342: begin
            cosine_reg0 <= 36'sb100011000011111101010111100010001000;
            sine_reg0   <= 36'sb110010010101110010011001001110100110;
        end
        9343: begin
            cosine_reg0 <= 36'sb100011000100010010110101010011010000;
            sine_reg0   <= 36'sb110010010101000100111100010011111101;
        end
        9344: begin
            cosine_reg0 <= 36'sb100011000100101000010100001011110010;
            sine_reg0   <= 36'sb110010010100010111011111111011000100;
        end
        9345: begin
            cosine_reg0 <= 36'sb100011000100111101110100001011101011;
            sine_reg0   <= 36'sb110010010011101010000100000011111100;
        end
        9346: begin
            cosine_reg0 <= 36'sb100011000101010011010101010010111100;
            sine_reg0   <= 36'sb110010010010111100101000101110100101;
        end
        9347: begin
            cosine_reg0 <= 36'sb100011000101101000110111100001100011;
            sine_reg0   <= 36'sb110010010010001111001101111011000011;
        end
        9348: begin
            cosine_reg0 <= 36'sb100011000101111110011010110111100000;
            sine_reg0   <= 36'sb110010010001100001110011101001010110;
        end
        9349: begin
            cosine_reg0 <= 36'sb100011000110010011111111010100110010;
            sine_reg0   <= 36'sb110010010000110100011001111001100001;
        end
        9350: begin
            cosine_reg0 <= 36'sb100011000110101001100100111001010111;
            sine_reg0   <= 36'sb110010010000000111000000101011100101;
        end
        9351: begin
            cosine_reg0 <= 36'sb100011000110111111001011100101010000;
            sine_reg0   <= 36'sb110010001111011001100111111111100101;
        end
        9352: begin
            cosine_reg0 <= 36'sb100011000111010100110011011000011010;
            sine_reg0   <= 36'sb110010001110101100001111110101100001;
        end
        9353: begin
            cosine_reg0 <= 36'sb100011000111101010011100010010110111;
            sine_reg0   <= 36'sb110010001101111110111000001101011011;
        end
        9354: begin
            cosine_reg0 <= 36'sb100011001000000000000110010100100100;
            sine_reg0   <= 36'sb110010001101010001100001000111010110;
        end
        9355: begin
            cosine_reg0 <= 36'sb100011001000010101110001011101100000;
            sine_reg0   <= 36'sb110010001100100100001010100011010011;
        end
        9356: begin
            cosine_reg0 <= 36'sb100011001000101011011101101101101100;
            sine_reg0   <= 36'sb110010001011110110110100100001010100;
        end
        9357: begin
            cosine_reg0 <= 36'sb100011001001000001001011000101000101;
            sine_reg0   <= 36'sb110010001011001001011111000001011010;
        end
        9358: begin
            cosine_reg0 <= 36'sb100011001001010110111001100011101100;
            sine_reg0   <= 36'sb110010001010011100001010000011101000;
        end
        9359: begin
            cosine_reg0 <= 36'sb100011001001101100101001001001011111;
            sine_reg0   <= 36'sb110010001001101110110101100111111110;
        end
        9360: begin
            cosine_reg0 <= 36'sb100011001010000010011001110110011110;
            sine_reg0   <= 36'sb110010001001000001100001101110100000;
        end
        9361: begin
            cosine_reg0 <= 36'sb100011001010011000001011101010101000;
            sine_reg0   <= 36'sb110010001000010100001110010111001110;
        end
        9362: begin
            cosine_reg0 <= 36'sb100011001010101101111110100101111011;
            sine_reg0   <= 36'sb110010000111100110111011100010001010;
        end
        9363: begin
            cosine_reg0 <= 36'sb100011001011000011110010101000011000;
            sine_reg0   <= 36'sb110010000110111001101001001111010110;
        end
        9364: begin
            cosine_reg0 <= 36'sb100011001011011001100111110001111100;
            sine_reg0   <= 36'sb110010000110001100010111011110110100;
        end
        9365: begin
            cosine_reg0 <= 36'sb100011001011101111011110000010101000;
            sine_reg0   <= 36'sb110010000101011111000110010000100110;
        end
        9366: begin
            cosine_reg0 <= 36'sb100011001100000101010101011010011011;
            sine_reg0   <= 36'sb110010000100110001110101100100101100;
        end
        9367: begin
            cosine_reg0 <= 36'sb100011001100011011001101111001010011;
            sine_reg0   <= 36'sb110010000100000100100101011011001010;
        end
        9368: begin
            cosine_reg0 <= 36'sb100011001100110001000111011111010000;
            sine_reg0   <= 36'sb110010000011010111010101110100000000;
        end
        9369: begin
            cosine_reg0 <= 36'sb100011001101000111000010001100010001;
            sine_reg0   <= 36'sb110010000010101010000110101111010001;
        end
        9370: begin
            cosine_reg0 <= 36'sb100011001101011100111110000000010110;
            sine_reg0   <= 36'sb110010000001111100111000001100111111;
        end
        9371: begin
            cosine_reg0 <= 36'sb100011001101110010111010111011011100;
            sine_reg0   <= 36'sb110010000001001111101010001101001010;
        end
        9372: begin
            cosine_reg0 <= 36'sb100011001110001000111000111101100100;
            sine_reg0   <= 36'sb110010000000100010011100101111110101;
        end
        9373: begin
            cosine_reg0 <= 36'sb100011001110011110111000000110101101;
            sine_reg0   <= 36'sb110001111111110101001111110101000001;
        end
        9374: begin
            cosine_reg0 <= 36'sb100011001110110100111000010110110101;
            sine_reg0   <= 36'sb110001111111001000000011011100110001;
        end
        9375: begin
            cosine_reg0 <= 36'sb100011001111001010111001101101111100;
            sine_reg0   <= 36'sb110001111110011010110111100111000101;
        end
        9376: begin
            cosine_reg0 <= 36'sb100011001111100000111100001100000010;
            sine_reg0   <= 36'sb110001111101101101101100010100000000;
        end
        9377: begin
            cosine_reg0 <= 36'sb100011001111110110111111110001000100;
            sine_reg0   <= 36'sb110001111101000000100001100011100100;
        end
        9378: begin
            cosine_reg0 <= 36'sb100011010000001101000100011101000011;
            sine_reg0   <= 36'sb110001111100010011010111010101110010;
        end
        9379: begin
            cosine_reg0 <= 36'sb100011010000100011001010001111111110;
            sine_reg0   <= 36'sb110001111011100110001101101010101011;
        end
        9380: begin
            cosine_reg0 <= 36'sb100011010000111001010001001001110011;
            sine_reg0   <= 36'sb110001111010111001000100100010010011;
        end
        9381: begin
            cosine_reg0 <= 36'sb100011010001001111011001001010100010;
            sine_reg0   <= 36'sb110001111010001011111011111100101010;
        end
        9382: begin
            cosine_reg0 <= 36'sb100011010001100101100010010010001001;
            sine_reg0   <= 36'sb110001111001011110110011111001110001;
        end
        9383: begin
            cosine_reg0 <= 36'sb100011010001111011101100100000101001;
            sine_reg0   <= 36'sb110001111000110001101100011001101100;
        end
        9384: begin
            cosine_reg0 <= 36'sb100011010010010001110111110110000001;
            sine_reg0   <= 36'sb110001111000000100100101011100011100;
        end
        9385: begin
            cosine_reg0 <= 36'sb100011010010101000000100010010001110;
            sine_reg0   <= 36'sb110001110111010111011111000010000001;
        end
        9386: begin
            cosine_reg0 <= 36'sb100011010010111110010001110101010001;
            sine_reg0   <= 36'sb110001110110101010011001001010011111;
        end
        9387: begin
            cosine_reg0 <= 36'sb100011010011010100100000011111001001;
            sine_reg0   <= 36'sb110001110101111101010011110101110111;
        end
        9388: begin
            cosine_reg0 <= 36'sb100011010011101010110000001111110101;
            sine_reg0   <= 36'sb110001110101010000001111000100001010;
        end
        9389: begin
            cosine_reg0 <= 36'sb100011010100000001000001000111010100;
            sine_reg0   <= 36'sb110001110100100011001010110101011011;
        end
        9390: begin
            cosine_reg0 <= 36'sb100011010100010111010011000101100100;
            sine_reg0   <= 36'sb110001110011110110000111001001101010;
        end
        9391: begin
            cosine_reg0 <= 36'sb100011010100101101100110001010100110;
            sine_reg0   <= 36'sb110001110011001001000100000000111011;
        end
        9392: begin
            cosine_reg0 <= 36'sb100011010101000011111010010110011001;
            sine_reg0   <= 36'sb110001110010011100000001011011001110;
        end
        9393: begin
            cosine_reg0 <= 36'sb100011010101011010001111101000111011;
            sine_reg0   <= 36'sb110001110001101110111111011000100101;
        end
        9394: begin
            cosine_reg0 <= 36'sb100011010101110000100110000010001011;
            sine_reg0   <= 36'sb110001110001000001111101111001000010;
        end
        9395: begin
            cosine_reg0 <= 36'sb100011010110000110111101100010001010;
            sine_reg0   <= 36'sb110001110000010100111100111100100111;
        end
        9396: begin
            cosine_reg0 <= 36'sb100011010110011101010110001000110101;
            sine_reg0   <= 36'sb110001101111100111111100100011010101;
        end
        9397: begin
            cosine_reg0 <= 36'sb100011010110110011101111110110001100;
            sine_reg0   <= 36'sb110001101110111010111100101101001111;
        end
        9398: begin
            cosine_reg0 <= 36'sb100011010111001010001010101010001111;
            sine_reg0   <= 36'sb110001101110001101111101011010010101;
        end
        9399: begin
            cosine_reg0 <= 36'sb100011010111100000100110100100111100;
            sine_reg0   <= 36'sb110001101101100000111110101010101010;
        end
        9400: begin
            cosine_reg0 <= 36'sb100011010111110111000011100110010010;
            sine_reg0   <= 36'sb110001101100110100000000011110010000;
        end
        9401: begin
            cosine_reg0 <= 36'sb100011011000001101100001101110010010;
            sine_reg0   <= 36'sb110001101100000111000010110101000111;
        end
        9402: begin
            cosine_reg0 <= 36'sb100011011000100100000000111100111000;
            sine_reg0   <= 36'sb110001101011011010000101101111010011;
        end
        9403: begin
            cosine_reg0 <= 36'sb100011011000111010100001010010000110;
            sine_reg0   <= 36'sb110001101010101101001001001100110100;
        end
        9404: begin
            cosine_reg0 <= 36'sb100011011001010001000010101101111010;
            sine_reg0   <= 36'sb110001101010000000001101001101101100;
        end
        9405: begin
            cosine_reg0 <= 36'sb100011011001100111100101010000010011;
            sine_reg0   <= 36'sb110001101001010011010001110001111110;
        end
        9406: begin
            cosine_reg0 <= 36'sb100011011001111110001000111001010000;
            sine_reg0   <= 36'sb110001101000100110010110111001101010;
        end
        9407: begin
            cosine_reg0 <= 36'sb100011011010010100101101101000110001;
            sine_reg0   <= 36'sb110001100111111001011100100100110011;
        end
        9408: begin
            cosine_reg0 <= 36'sb100011011010101011010011011110110100;
            sine_reg0   <= 36'sb110001100111001100100010110011011010;
        end
        9409: begin
            cosine_reg0 <= 36'sb100011011011000001111010011011011001;
            sine_reg0   <= 36'sb110001100110011111101001100101100001;
        end
        9410: begin
            cosine_reg0 <= 36'sb100011011011011000100010011110011110;
            sine_reg0   <= 36'sb110001100101110010110000111011001010;
        end
        9411: begin
            cosine_reg0 <= 36'sb100011011011101111001011101000000100;
            sine_reg0   <= 36'sb110001100101000101111000110100010110;
        end
        9412: begin
            cosine_reg0 <= 36'sb100011011100000101110101111000001001;
            sine_reg0   <= 36'sb110001100100011001000001010001001000;
        end
        9413: begin
            cosine_reg0 <= 36'sb100011011100011100100001001110101011;
            sine_reg0   <= 36'sb110001100011101100001010010001100000;
        end
        9414: begin
            cosine_reg0 <= 36'sb100011011100110011001101101011101100;
            sine_reg0   <= 36'sb110001100010111111010011110101100001;
        end
        9415: begin
            cosine_reg0 <= 36'sb100011011101001001111011001111001000;
            sine_reg0   <= 36'sb110001100010010010011101111101001101;
        end
        9416: begin
            cosine_reg0 <= 36'sb100011011101100000101001111001000000;
            sine_reg0   <= 36'sb110001100001100101101000101000100100;
        end
        9417: begin
            cosine_reg0 <= 36'sb100011011101110111011001101001010011;
            sine_reg0   <= 36'sb110001100000111000110011110111101010;
        end
        9418: begin
            cosine_reg0 <= 36'sb100011011110001110001010100000000000;
            sine_reg0   <= 36'sb110001100000001011111111101010011110;
        end
        9419: begin
            cosine_reg0 <= 36'sb100011011110100100111100011101000101;
            sine_reg0   <= 36'sb110001011111011111001100000001000101;
        end
        9420: begin
            cosine_reg0 <= 36'sb100011011110111011101111100000100011;
            sine_reg0   <= 36'sb110001011110110010011000111011011110;
        end
        9421: begin
            cosine_reg0 <= 36'sb100011011111010010100011101010011000;
            sine_reg0   <= 36'sb110001011110000101100110011001101100;
        end
        9422: begin
            cosine_reg0 <= 36'sb100011011111101001011000111010100011;
            sine_reg0   <= 36'sb110001011101011000110100011011110000;
        end
        9423: begin
            cosine_reg0 <= 36'sb100011100000000000001111010001000011;
            sine_reg0   <= 36'sb110001011100101100000011000001101101;
        end
        9424: begin
            cosine_reg0 <= 36'sb100011100000010111000110101101111000;
            sine_reg0   <= 36'sb110001011011111111010010001011100011;
        end
        9425: begin
            cosine_reg0 <= 36'sb100011100000101101111111010001000001;
            sine_reg0   <= 36'sb110001011011010010100001111001010101;
        end
        9426: begin
            cosine_reg0 <= 36'sb100011100001000100111000111010011100;
            sine_reg0   <= 36'sb110001011010100101110010001011000101;
        end
        9427: begin
            cosine_reg0 <= 36'sb100011100001011011110011101010001001;
            sine_reg0   <= 36'sb110001011001111001000011000000110100;
        end
        9428: begin
            cosine_reg0 <= 36'sb100011100001110010101111100000001000;
            sine_reg0   <= 36'sb110001011001001100010100011010100011;
        end
        9429: begin
            cosine_reg0 <= 36'sb100011100010001001101100011100010110;
            sine_reg0   <= 36'sb110001011000011111100110011000010101;
        end
        9430: begin
            cosine_reg0 <= 36'sb100011100010100000101010011110110100;
            sine_reg0   <= 36'sb110001010111110010111000111010001011;
        end
        9431: begin
            cosine_reg0 <= 36'sb100011100010110111101001100111100000;
            sine_reg0   <= 36'sb110001010111000110001100000000000111;
        end
        9432: begin
            cosine_reg0 <= 36'sb100011100011001110101001110110011001;
            sine_reg0   <= 36'sb110001010110011001011111101010001011;
        end
        9433: begin
            cosine_reg0 <= 36'sb100011100011100101101011001011011111;
            sine_reg0   <= 36'sb110001010101101100110011111000011001;
        end
        9434: begin
            cosine_reg0 <= 36'sb100011100011111100101101100110110001;
            sine_reg0   <= 36'sb110001010101000000001000101010110001;
        end
        9435: begin
            cosine_reg0 <= 36'sb100011100100010011110001001000001101;
            sine_reg0   <= 36'sb110001010100010011011110000001010111;
        end
        9436: begin
            cosine_reg0 <= 36'sb100011100100101010110101101111110100;
            sine_reg0   <= 36'sb110001010011100110110011111100001011;
        end
        9437: begin
            cosine_reg0 <= 36'sb100011100101000001111011011101100011;
            sine_reg0   <= 36'sb110001010010111010001010011011001111;
        end
        9438: begin
            cosine_reg0 <= 36'sb100011100101011001000010010001011011;
            sine_reg0   <= 36'sb110001010010001101100001011110100110;
        end
        9439: begin
            cosine_reg0 <= 36'sb100011100101110000001010001011011010;
            sine_reg0   <= 36'sb110001010001100000111001000110010000;
        end
        9440: begin
            cosine_reg0 <= 36'sb100011100110000111010011001011011111;
            sine_reg0   <= 36'sb110001010000110100010001010010010000;
        end
        9441: begin
            cosine_reg0 <= 36'sb100011100110011110011101010001101001;
            sine_reg0   <= 36'sb110001010000000111101010000010100111;
        end
        9442: begin
            cosine_reg0 <= 36'sb100011100110110101101000011101111001;
            sine_reg0   <= 36'sb110001001111011011000011010111010110;
        end
        9443: begin
            cosine_reg0 <= 36'sb100011100111001100110100110000001011;
            sine_reg0   <= 36'sb110001001110101110011101010000100001;
        end
        9444: begin
            cosine_reg0 <= 36'sb100011100111100100000010001000100001;
            sine_reg0   <= 36'sb110001001110000001110111101110001000;
        end
        9445: begin
            cosine_reg0 <= 36'sb100011100111111011010000100110111000;
            sine_reg0   <= 36'sb110001001101010101010010110000001101;
        end
        9446: begin
            cosine_reg0 <= 36'sb100011101000010010100000001011010001;
            sine_reg0   <= 36'sb110001001100101000101110010110110001;
        end
        9447: begin
            cosine_reg0 <= 36'sb100011101000101001110000110101101001;
            sine_reg0   <= 36'sb110001001011111100001010100001111000;
        end
        9448: begin
            cosine_reg0 <= 36'sb100011101001000001000010100110000001;
            sine_reg0   <= 36'sb110001001011001111100111010001100001;
        end
        9449: begin
            cosine_reg0 <= 36'sb100011101001011000010101011100010111;
            sine_reg0   <= 36'sb110001001010100011000100100101110000;
        end
        9450: begin
            cosine_reg0 <= 36'sb100011101001101111101001011000101011;
            sine_reg0   <= 36'sb110001001001110110100010011110100101;
        end
        9451: begin
            cosine_reg0 <= 36'sb100011101010000110111110011010111011;
            sine_reg0   <= 36'sb110001001001001010000000111100000010;
        end
        9452: begin
            cosine_reg0 <= 36'sb100011101010011110010100100011000110;
            sine_reg0   <= 36'sb110001001000011101011111111110001010;
        end
        9453: begin
            cosine_reg0 <= 36'sb100011101010110101101011110001001100;
            sine_reg0   <= 36'sb110001000111110000111111100100111110;
        end
        9454: begin
            cosine_reg0 <= 36'sb100011101011001101000100000101001100;
            sine_reg0   <= 36'sb110001000111000100011111110000011111;
        end
        9455: begin
            cosine_reg0 <= 36'sb100011101011100100011101011111000101;
            sine_reg0   <= 36'sb110001000110011000000000100000101111;
        end
        9456: begin
            cosine_reg0 <= 36'sb100011101011111011110111111110110110;
            sine_reg0   <= 36'sb110001000101101011100001110101110000;
        end
        9457: begin
            cosine_reg0 <= 36'sb100011101100010011010011100100011110;
            sine_reg0   <= 36'sb110001000100111111000011101111100100;
        end
        9458: begin
            cosine_reg0 <= 36'sb100011101100101010110000001111111100;
            sine_reg0   <= 36'sb110001000100010010100110001110001101;
        end
        9459: begin
            cosine_reg0 <= 36'sb100011101101000010001110000001010000;
            sine_reg0   <= 36'sb110001000011100110001001010001101011;
        end
        9460: begin
            cosine_reg0 <= 36'sb100011101101011001101100111000010111;
            sine_reg0   <= 36'sb110001000010111001101100111010000001;
        end
        9461: begin
            cosine_reg0 <= 36'sb100011101101110001001100110101010011;
            sine_reg0   <= 36'sb110001000010001101010001000111010001;
        end
        9462: begin
            cosine_reg0 <= 36'sb100011101110001000101101111000000001;
            sine_reg0   <= 36'sb110001000001100000110101111001011100;
        end
        9463: begin
            cosine_reg0 <= 36'sb100011101110100000010000000000100000;
            sine_reg0   <= 36'sb110001000000110100011011010000100101;
        end
        9464: begin
            cosine_reg0 <= 36'sb100011101110110111110011001110110000;
            sine_reg0   <= 36'sb110001000000001000000001001100101011;
        end
        9465: begin
            cosine_reg0 <= 36'sb100011101111001111010111100010110001;
            sine_reg0   <= 36'sb110000111111011011100111101101110010;
        end
        9466: begin
            cosine_reg0 <= 36'sb100011101111100110111100111100100000;
            sine_reg0   <= 36'sb110000111110101111001110110011111100;
        end
        9467: begin
            cosine_reg0 <= 36'sb100011101111111110100011011011111101;
            sine_reg0   <= 36'sb110000111110000010110110011111001001;
        end
        9468: begin
            cosine_reg0 <= 36'sb100011110000010110001011000001000111;
            sine_reg0   <= 36'sb110000111101010110011110101111011100;
        end
        9469: begin
            cosine_reg0 <= 36'sb100011110000101101110011101011111101;
            sine_reg0   <= 36'sb110000111100101010000111100100110101;
        end
        9470: begin
            cosine_reg0 <= 36'sb100011110001000101011101011100011111;
            sine_reg0   <= 36'sb110000111011111101110000111111011000;
        end
        9471: begin
            cosine_reg0 <= 36'sb100011110001011101001000010010101011;
            sine_reg0   <= 36'sb110000111011010001011010111111000110;
        end
        9472: begin
            cosine_reg0 <= 36'sb100011110001110100110100001110100001;
            sine_reg0   <= 36'sb110000111010100101000101100100000000;
        end
        9473: begin
            cosine_reg0 <= 36'sb100011110010001100100001001111111111;
            sine_reg0   <= 36'sb110000111001111000110000101110001000;
        end
        9474: begin
            cosine_reg0 <= 36'sb100011110010100100001111010111000101;
            sine_reg0   <= 36'sb110000111001001100011100011101011111;
        end
        9475: begin
            cosine_reg0 <= 36'sb100011110010111011111110100011110001;
            sine_reg0   <= 36'sb110000111000100000001000110010001001;
        end
        9476: begin
            cosine_reg0 <= 36'sb100011110011010011101110110110000011;
            sine_reg0   <= 36'sb110000110111110011110101101100000101;
        end
        9477: begin
            cosine_reg0 <= 36'sb100011110011101011100000001101111011;
            sine_reg0   <= 36'sb110000110111000111100011001011010110;
        end
        9478: begin
            cosine_reg0 <= 36'sb100011110100000011010010101011010110;
            sine_reg0   <= 36'sb110000110110011011010001001111111110;
        end
        9479: begin
            cosine_reg0 <= 36'sb100011110100011011000110001110010100;
            sine_reg0   <= 36'sb110000110101101110111111111001111111;
        end
        9480: begin
            cosine_reg0 <= 36'sb100011110100110010111010110110110100;
            sine_reg0   <= 36'sb110000110101000010101111001001011001;
        end
        9481: begin
            cosine_reg0 <= 36'sb100011110101001010110000100100110110;
            sine_reg0   <= 36'sb110000110100010110011110111110001111;
        end
        9482: begin
            cosine_reg0 <= 36'sb100011110101100010100111011000011000;
            sine_reg0   <= 36'sb110000110011101010001111011000100010;
        end
        9483: begin
            cosine_reg0 <= 36'sb100011110101111010011111010001011001;
            sine_reg0   <= 36'sb110000110010111110000000011000010101;
        end
        9484: begin
            cosine_reg0 <= 36'sb100011110110010010011000001111111001;
            sine_reg0   <= 36'sb110000110010010001110001111101101001;
        end
        9485: begin
            cosine_reg0 <= 36'sb100011110110101010010010010011110110;
            sine_reg0   <= 36'sb110000110001100101100100001000011111;
        end
        9486: begin
            cosine_reg0 <= 36'sb100011110111000010001101011101010000;
            sine_reg0   <= 36'sb110000110000111001010110111000111001;
        end
        9487: begin
            cosine_reg0 <= 36'sb100011110111011010001001101100000110;
            sine_reg0   <= 36'sb110000110000001101001010001110111001;
        end
        9488: begin
            cosine_reg0 <= 36'sb100011110111110010000111000000010111;
            sine_reg0   <= 36'sb110000101111100000111110001010100001;
        end
        9489: begin
            cosine_reg0 <= 36'sb100011111000001010000101011010000001;
            sine_reg0   <= 36'sb110000101110110100110010101011110011;
        end
        9490: begin
            cosine_reg0 <= 36'sb100011111000100010000100111001000100;
            sine_reg0   <= 36'sb110000101110001000100111110010101111;
        end
        9491: begin
            cosine_reg0 <= 36'sb100011111000111010000101011101011111;
            sine_reg0   <= 36'sb110000101101011100011101011111011001;
        end
        9492: begin
            cosine_reg0 <= 36'sb100011111001010010000111000111010010;
            sine_reg0   <= 36'sb110000101100110000010011110001110000;
        end
        9493: begin
            cosine_reg0 <= 36'sb100011111001101010001001110110011010;
            sine_reg0   <= 36'sb110000101100000100001010101001111000;
        end
        9494: begin
            cosine_reg0 <= 36'sb100011111010000010001101101010111000;
            sine_reg0   <= 36'sb110000101011011000000010000111110010;
        end
        9495: begin
            cosine_reg0 <= 36'sb100011111010011010010010100100101010;
            sine_reg0   <= 36'sb110000101010101011111010001011011111;
        end
        9496: begin
            cosine_reg0 <= 36'sb100011111010110010011000100011101111;
            sine_reg0   <= 36'sb110000101001111111110010110101000010;
        end
        9497: begin
            cosine_reg0 <= 36'sb100011111011001010011111101000000111;
            sine_reg0   <= 36'sb110000101001010011101100000100011100;
        end
        9498: begin
            cosine_reg0 <= 36'sb100011111011100010100111110001110000;
            sine_reg0   <= 36'sb110000101000100111100101111001101110;
        end
        9499: begin
            cosine_reg0 <= 36'sb100011111011111010110001000000101010;
            sine_reg0   <= 36'sb110000100111111011100000010100111011;
        end
        9500: begin
            cosine_reg0 <= 36'sb100011111100010010111011010100110100;
            sine_reg0   <= 36'sb110000100111001111011011010110000100;
        end
        9501: begin
            cosine_reg0 <= 36'sb100011111100101011000110101110001100;
            sine_reg0   <= 36'sb110000100110100011010110111101001011;
        end
        9502: begin
            cosine_reg0 <= 36'sb100011111101000011010011001100110010;
            sine_reg0   <= 36'sb110000100101110111010011001010010001;
        end
        9503: begin
            cosine_reg0 <= 36'sb100011111101011011100000110000100101;
            sine_reg0   <= 36'sb110000100101001011001111111101011000;
        end
        9504: begin
            cosine_reg0 <= 36'sb100011111101110011101111011001100100;
            sine_reg0   <= 36'sb110000100100011111001101010110100011;
        end
        9505: begin
            cosine_reg0 <= 36'sb100011111110001011111111000111101110;
            sine_reg0   <= 36'sb110000100011110011001011010101110001;
        end
        9506: begin
            cosine_reg0 <= 36'sb100011111110100100001111111011000010;
            sine_reg0   <= 36'sb110000100011000111001001111011000111;
        end
        9507: begin
            cosine_reg0 <= 36'sb100011111110111100100001110011011111;
            sine_reg0   <= 36'sb110000100010011011001001000110100100;
        end
        9508: begin
            cosine_reg0 <= 36'sb100011111111010100110100110001000100;
            sine_reg0   <= 36'sb110000100001101111001000111000001011;
        end
        9509: begin
            cosine_reg0 <= 36'sb100011111111101101001000110011110001;
            sine_reg0   <= 36'sb110000100001000011001001001111111101;
        end
        9510: begin
            cosine_reg0 <= 36'sb100100000000000101011101111011100100;
            sine_reg0   <= 36'sb110000100000010111001010001101111100;
        end
        9511: begin
            cosine_reg0 <= 36'sb100100000000011101110100001000011100;
            sine_reg0   <= 36'sb110000011111101011001011110010001010;
        end
        9512: begin
            cosine_reg0 <= 36'sb100100000000110110001011011010011000;
            sine_reg0   <= 36'sb110000011110111111001101111100101000;
        end
        9513: begin
            cosine_reg0 <= 36'sb100100000001001110100011110001011001;
            sine_reg0   <= 36'sb110000011110010011010000101101011001;
        end
        9514: begin
            cosine_reg0 <= 36'sb100100000001100110111101001101011011;
            sine_reg0   <= 36'sb110000011101100111010100000100011110;
        end
        9515: begin
            cosine_reg0 <= 36'sb100100000001111111010111101110011111;
            sine_reg0   <= 36'sb110000011100111011011000000001111000;
        end
        9516: begin
            cosine_reg0 <= 36'sb100100000010010111110011010100100100;
            sine_reg0   <= 36'sb110000011100001111011100100101101001;
        end
        9517: begin
            cosine_reg0 <= 36'sb100100000010110000001111111111101001;
            sine_reg0   <= 36'sb110000011011100011100001101111110011;
        end
        9518: begin
            cosine_reg0 <= 36'sb100100000011001000101101101111101101;
            sine_reg0   <= 36'sb110000011010110111100111100000011000;
        end
        9519: begin
            cosine_reg0 <= 36'sb100100000011100001001100100100101110;
            sine_reg0   <= 36'sb110000011010001011101101110111011001;
        end
        9520: begin
            cosine_reg0 <= 36'sb100100000011111001101100011110101100;
            sine_reg0   <= 36'sb110000011001011111110100110100111001;
        end
        9521: begin
            cosine_reg0 <= 36'sb100100000100010010001101011101100110;
            sine_reg0   <= 36'sb110000011000110011111100011000110111;
        end
        9522: begin
            cosine_reg0 <= 36'sb100100000100101010101111100001011011;
            sine_reg0   <= 36'sb110000011000001000000100100011011000;
        end
        9523: begin
            cosine_reg0 <= 36'sb100100000101000011010010101010001011;
            sine_reg0   <= 36'sb110000010111011100001101010100011011;
        end
        9524: begin
            cosine_reg0 <= 36'sb100100000101011011110110110111110011;
            sine_reg0   <= 36'sb110000010110110000010110101100000011;
        end
        9525: begin
            cosine_reg0 <= 36'sb100100000101110100011100001010010011;
            sine_reg0   <= 36'sb110000010110000100100000101010010010;
        end
        9526: begin
            cosine_reg0 <= 36'sb100100000110001101000010100001101011;
            sine_reg0   <= 36'sb110000010101011000101011001111001001;
        end
        9527: begin
            cosine_reg0 <= 36'sb100100000110100101101001111101111001;
            sine_reg0   <= 36'sb110000010100101100110110011010101001;
        end
        9528: begin
            cosine_reg0 <= 36'sb100100000110111110010010011110111101;
            sine_reg0   <= 36'sb110000010100000001000010001100110110;
        end
        9529: begin
            cosine_reg0 <= 36'sb100100000111010110111100000100110100;
            sine_reg0   <= 36'sb110000010011010101001110100101101111;
        end
        9530: begin
            cosine_reg0 <= 36'sb100100000111101111100110101111011111;
            sine_reg0   <= 36'sb110000010010101001011011100101010111;
        end
        9531: begin
            cosine_reg0 <= 36'sb100100001000001000010010011110111101;
            sine_reg0   <= 36'sb110000010001111101101001001011110000;
        end
        9532: begin
            cosine_reg0 <= 36'sb100100001000100000111111010011001100;
            sine_reg0   <= 36'sb110000010001010001110111011000111100;
        end
        9533: begin
            cosine_reg0 <= 36'sb100100001000111001101101001100001100;
            sine_reg0   <= 36'sb110000010000100110000110001100111011;
        end
        9534: begin
            cosine_reg0 <= 36'sb100100001001010010011100001001111011;
            sine_reg0   <= 36'sb110000001111111010010101100111110000;
        end
        9535: begin
            cosine_reg0 <= 36'sb100100001001101011001100001100011001;
            sine_reg0   <= 36'sb110000001111001110100101101001011100;
        end
        9536: begin
            cosine_reg0 <= 36'sb100100001010000011111101010011100101;
            sine_reg0   <= 36'sb110000001110100010110110010010000001;
        end
        9537: begin
            cosine_reg0 <= 36'sb100100001010011100101111011111011101;
            sine_reg0   <= 36'sb110000001101110111000111100001100001;
        end
        9538: begin
            cosine_reg0 <= 36'sb100100001010110101100010110000000010;
            sine_reg0   <= 36'sb110000001101001011011001010111111110;
        end
        9539: begin
            cosine_reg0 <= 36'sb100100001011001110010111000101010001;
            sine_reg0   <= 36'sb110000001100011111101011110101011001;
        end
        9540: begin
            cosine_reg0 <= 36'sb100100001011100111001100011111001010;
            sine_reg0   <= 36'sb110000001011110011111110111001110011;
        end
        9541: begin
            cosine_reg0 <= 36'sb100100001100000000000010111101101100;
            sine_reg0   <= 36'sb110000001011001000010010100101001111;
        end
        9542: begin
            cosine_reg0 <= 36'sb100100001100011000111010100000110110;
            sine_reg0   <= 36'sb110000001010011100100110110111101110;
        end
        9543: begin
            cosine_reg0 <= 36'sb100100001100110001110011001000100111;
            sine_reg0   <= 36'sb110000001001110000111011110001010010;
        end
        9544: begin
            cosine_reg0 <= 36'sb100100001101001010101100110100111110;
            sine_reg0   <= 36'sb110000001001000101010001010001111100;
        end
        9545: begin
            cosine_reg0 <= 36'sb100100001101100011100111100101111010;
            sine_reg0   <= 36'sb110000001000011001100111011001101110;
        end
        9546: begin
            cosine_reg0 <= 36'sb100100001101111100100011011011011010;
            sine_reg0   <= 36'sb110000000111101101111110001000101011;
        end
        9547: begin
            cosine_reg0 <= 36'sb100100001110010101100000010101011101;
            sine_reg0   <= 36'sb110000000111000010010101011110110011;
        end
        9548: begin
            cosine_reg0 <= 36'sb100100001110101110011110010100000011;
            sine_reg0   <= 36'sb110000000110010110101101011100001000;
        end
        9549: begin
            cosine_reg0 <= 36'sb100100001111000111011101010111001010;
            sine_reg0   <= 36'sb110000000101101011000110000000101100;
        end
        9550: begin
            cosine_reg0 <= 36'sb100100001111100000011101011110110001;
            sine_reg0   <= 36'sb110000000100111111011111001100100001;
        end
        9551: begin
            cosine_reg0 <= 36'sb100100001111111001011110101010110111;
            sine_reg0   <= 36'sb110000000100010011111000111111101000;
        end
        9552: begin
            cosine_reg0 <= 36'sb100100010000010010100000111011011100;
            sine_reg0   <= 36'sb110000000011101000010011011010000100;
        end
        9553: begin
            cosine_reg0 <= 36'sb100100010000101011100100010000011110;
            sine_reg0   <= 36'sb110000000010111100101110011011110100;
        end
        9554: begin
            cosine_reg0 <= 36'sb100100010001000100101000101001111101;
            sine_reg0   <= 36'sb110000000010010001001010000100111101;
        end
        9555: begin
            cosine_reg0 <= 36'sb100100010001011101101110000111110111;
            sine_reg0   <= 36'sb110000000001100101100110010101011110;
        end
        9556: begin
            cosine_reg0 <= 36'sb100100010001110110110100101010001011;
            sine_reg0   <= 36'sb110000000000111010000011001101011010;
        end
        9557: begin
            cosine_reg0 <= 36'sb100100010010001111111100010000111001;
            sine_reg0   <= 36'sb110000000000001110100000101100110010;
        end
        9558: begin
            cosine_reg0 <= 36'sb100100010010101001000100111100000000;
            sine_reg0   <= 36'sb101111111111100010111110110011101000;
        end
        9559: begin
            cosine_reg0 <= 36'sb100100010011000010001110101011011110;
            sine_reg0   <= 36'sb101111111110110111011101100001111110;
        end
        9560: begin
            cosine_reg0 <= 36'sb100100010011011011011001011111010011;
            sine_reg0   <= 36'sb101111111110001011111100110111110110;
        end
        9561: begin
            cosine_reg0 <= 36'sb100100010011110100100101010111011110;
            sine_reg0   <= 36'sb101111111101100000011100110101010000;
        end
        9562: begin
            cosine_reg0 <= 36'sb100100010100001101110010010011111101;
            sine_reg0   <= 36'sb101111111100110100111101011010001111;
        end
        9563: begin
            cosine_reg0 <= 36'sb100100010100100111000000010100110000;
            sine_reg0   <= 36'sb101111111100001001011110100110110101;
        end
        9564: begin
            cosine_reg0 <= 36'sb100100010101000000001111011001110101;
            sine_reg0   <= 36'sb101111111011011110000000011011000011;
        end
        9565: begin
            cosine_reg0 <= 36'sb100100010101011001011111100011001101;
            sine_reg0   <= 36'sb101111111010110010100010110110111011;
        end
        9566: begin
            cosine_reg0 <= 36'sb100100010101110010110000110000110101;
            sine_reg0   <= 36'sb101111111010000111000101111010011110;
        end
        9567: begin
            cosine_reg0 <= 36'sb100100010110001100000011000010101101;
            sine_reg0   <= 36'sb101111111001011011101001100101101110;
        end
        9568: begin
            cosine_reg0 <= 36'sb100100010110100101010110011000110011;
            sine_reg0   <= 36'sb101111111000110000001101111000101101;
        end
        9569: begin
            cosine_reg0 <= 36'sb100100010110111110101010110011001000;
            sine_reg0   <= 36'sb101111111000000100110010110011011101;
        end
        9570: begin
            cosine_reg0 <= 36'sb100100010111011000000000010001101010;
            sine_reg0   <= 36'sb101111110111011001011000010101111111;
        end
        9571: begin
            cosine_reg0 <= 36'sb100100010111110001010110110100010111;
            sine_reg0   <= 36'sb101111110110101101111110100000010101;
        end
        9572: begin
            cosine_reg0 <= 36'sb100100011000001010101110011011001111;
            sine_reg0   <= 36'sb101111110110000010100101010010100000;
        end
        9573: begin
            cosine_reg0 <= 36'sb100100011000100100000111000110010010;
            sine_reg0   <= 36'sb101111110101010111001100101100100010;
        end
        9574: begin
            cosine_reg0 <= 36'sb100100011000111101100000110101011101;
            sine_reg0   <= 36'sb101111110100101011110100101110011101;
        end
        9575: begin
            cosine_reg0 <= 36'sb100100011001010110111011101000110000;
            sine_reg0   <= 36'sb101111110100000000011101011000010011;
        end
        9576: begin
            cosine_reg0 <= 36'sb100100011001110000010111100000001011;
            sine_reg0   <= 36'sb101111110011010101000110101010000101;
        end
        9577: begin
            cosine_reg0 <= 36'sb100100011010001001110100011011101011;
            sine_reg0   <= 36'sb101111110010101001110000100011110101;
        end
        9578: begin
            cosine_reg0 <= 36'sb100100011010100011010010011011010000;
            sine_reg0   <= 36'sb101111110001111110011011000101100100;
        end
        9579: begin
            cosine_reg0 <= 36'sb100100011010111100110001011110111010;
            sine_reg0   <= 36'sb101111110001010011000110001111010101;
        end
        9580: begin
            cosine_reg0 <= 36'sb100100011011010110010001100110100110;
            sine_reg0   <= 36'sb101111110000100111110010000001001001;
        end
        9581: begin
            cosine_reg0 <= 36'sb100100011011101111110010110010010101;
            sine_reg0   <= 36'sb101111101111111100011110011011000001;
        end
        9582: begin
            cosine_reg0 <= 36'sb100100011100001001010101000010000101;
            sine_reg0   <= 36'sb101111101111010001001011011100111111;
        end
        9583: begin
            cosine_reg0 <= 36'sb100100011100100010111000010101110101;
            sine_reg0   <= 36'sb101111101110100101111001000111000101;
        end
        9584: begin
            cosine_reg0 <= 36'sb100100011100111100011100101101100100;
            sine_reg0   <= 36'sb101111101101111010100111011001010101;
        end
        9585: begin
            cosine_reg0 <= 36'sb100100011101010110000010001001010001;
            sine_reg0   <= 36'sb101111101101001111010110010011110000;
        end
        9586: begin
            cosine_reg0 <= 36'sb100100011101101111101000101000111011;
            sine_reg0   <= 36'sb101111101100100100000101110110011000;
        end
        9587: begin
            cosine_reg0 <= 36'sb100100011110001001010000001100100010;
            sine_reg0   <= 36'sb101111101011111000110110000001001110;
        end
        9588: begin
            cosine_reg0 <= 36'sb100100011110100010111000110100000100;
            sine_reg0   <= 36'sb101111101011001101100110110100010101;
        end
        9589: begin
            cosine_reg0 <= 36'sb100100011110111100100010011111100000;
            sine_reg0   <= 36'sb101111101010100010011000001111101110;
        end
        9590: begin
            cosine_reg0 <= 36'sb100100011111010110001101001110110101;
            sine_reg0   <= 36'sb101111101001110111001010010011011010;
        end
        9591: begin
            cosine_reg0 <= 36'sb100100011111101111111001000010000010;
            sine_reg0   <= 36'sb101111101001001011111100111111011100;
        end
        9592: begin
            cosine_reg0 <= 36'sb100100100000001001100101111001000111;
            sine_reg0   <= 36'sb101111101000100000110000010011110100;
        end
        9593: begin
            cosine_reg0 <= 36'sb100100100000100011010011110100000010;
            sine_reg0   <= 36'sb101111100111110101100100010000100101;
        end
        9594: begin
            cosine_reg0 <= 36'sb100100100000111101000010110010110010;
            sine_reg0   <= 36'sb101111100111001010011000110101110000;
        end
        9595: begin
            cosine_reg0 <= 36'sb100100100001010110110010110101010111;
            sine_reg0   <= 36'sb101111100110011111001110000011010111;
        end
        9596: begin
            cosine_reg0 <= 36'sb100100100001110000100011111011101110;
            sine_reg0   <= 36'sb101111100101110100000011111001011100;
        end
        9597: begin
            cosine_reg0 <= 36'sb100100100010001010010110000101111001;
            sine_reg0   <= 36'sb101111100101001000111010011000000000;
        end
        9598: begin
            cosine_reg0 <= 36'sb100100100010100100001001010011110100;
            sine_reg0   <= 36'sb101111100100011101110001011111000101;
        end
        9599: begin
            cosine_reg0 <= 36'sb100100100010111101111101100101100000;
            sine_reg0   <= 36'sb101111100011110010101001001110101100;
        end
        9600: begin
            cosine_reg0 <= 36'sb100100100011010111110010111010111011;
            sine_reg0   <= 36'sb101111100011000111100001100110111000;
        end
        9601: begin
            cosine_reg0 <= 36'sb100100100011110001101001010100000100;
            sine_reg0   <= 36'sb101111100010011100011010100111101001;
        end
        9602: begin
            cosine_reg0 <= 36'sb100100100100001011100000110000111010;
            sine_reg0   <= 36'sb101111100001110001010100010001000010;
        end
        9603: begin
            cosine_reg0 <= 36'sb100100100100100101011001010001011101;
            sine_reg0   <= 36'sb101111100001000110001110100011000100;
        end
        9604: begin
            cosine_reg0 <= 36'sb100100100100111111010010110101101011;
            sine_reg0   <= 36'sb101111100000011011001001011101110010;
        end
        9605: begin
            cosine_reg0 <= 36'sb100100100101011001001101011101100100;
            sine_reg0   <= 36'sb101111011111110000000101000001001011;
        end
        9606: begin
            cosine_reg0 <= 36'sb100100100101110011001001001001000110;
            sine_reg0   <= 36'sb101111011111000101000001001101010011;
        end
        9607: begin
            cosine_reg0 <= 36'sb100100100110001101000101111000010000;
            sine_reg0   <= 36'sb101111011110011001111110000010001011;
        end
        9608: begin
            cosine_reg0 <= 36'sb100100100110100111000011101011000001;
            sine_reg0   <= 36'sb101111011101101110111011011111110100;
        end
        9609: begin
            cosine_reg0 <= 36'sb100100100111000001000010100001011001;
            sine_reg0   <= 36'sb101111011101000011111001100110010000;
        end
        9610: begin
            cosine_reg0 <= 36'sb100100100111011011000010011011010110;
            sine_reg0   <= 36'sb101111011100011000111000010101100001;
        end
        9611: begin
            cosine_reg0 <= 36'sb100100100111110101000011011000111000;
            sine_reg0   <= 36'sb101111011011101101110111101101101001;
        end
        9612: begin
            cosine_reg0 <= 36'sb100100101000001111000101011001111100;
            sine_reg0   <= 36'sb101111011011000010110111101110101001;
        end
        9613: begin
            cosine_reg0 <= 36'sb100100101000101001001000011110100011;
            sine_reg0   <= 36'sb101111011010010111111000011000100010;
        end
        9614: begin
            cosine_reg0 <= 36'sb100100101001000011001100100110101100;
            sine_reg0   <= 36'sb101111011001101100111001101011010111;
        end
        9615: begin
            cosine_reg0 <= 36'sb100100101001011101010001110010010100;
            sine_reg0   <= 36'sb101111011001000001111011100111001010;
        end
        9616: begin
            cosine_reg0 <= 36'sb100100101001110111011000000001011100;
            sine_reg0   <= 36'sb101111011000010110111110001011111011;
        end
        9617: begin
            cosine_reg0 <= 36'sb100100101010010001011111010100000011;
            sine_reg0   <= 36'sb101111010111101100000001011001101100;
        end
        9618: begin
            cosine_reg0 <= 36'sb100100101010101011100111101010000110;
            sine_reg0   <= 36'sb101111010111000001000101010000011111;
        end
        9619: begin
            cosine_reg0 <= 36'sb100100101011000101110001000011100110;
            sine_reg0   <= 36'sb101111010110010110001001110000010111;
        end
        9620: begin
            cosine_reg0 <= 36'sb100100101011011111111011100000100001;
            sine_reg0   <= 36'sb101111010101101011001110111001010011;
        end
        9621: begin
            cosine_reg0 <= 36'sb100100101011111010000111000000110110;
            sine_reg0   <= 36'sb101111010101000000010100101011010111;
        end
        9622: begin
            cosine_reg0 <= 36'sb100100101100010100010011100100100101;
            sine_reg0   <= 36'sb101111010100010101011011000110100011;
        end
        9623: begin
            cosine_reg0 <= 36'sb100100101100101110100001001011101011;
            sine_reg0   <= 36'sb101111010011101010100010001010111010;
        end
        9624: begin
            cosine_reg0 <= 36'sb100100101101001000101111110110001001;
            sine_reg0   <= 36'sb101111010010111111101001111000011101;
        end
        9625: begin
            cosine_reg0 <= 36'sb100100101101100010111111100011111101;
            sine_reg0   <= 36'sb101111010010010100110010001111001101;
        end
        9626: begin
            cosine_reg0 <= 36'sb100100101101111101010000010101000111;
            sine_reg0   <= 36'sb101111010001101001111011001111001101;
        end
        9627: begin
            cosine_reg0 <= 36'sb100100101110010111100010001001100100;
            sine_reg0   <= 36'sb101111010000111111000100111000011101;
        end
        9628: begin
            cosine_reg0 <= 36'sb100100101110110001110101000001010101;
            sine_reg0   <= 36'sb101111010000010100001111001011000001;
        end
        9629: begin
            cosine_reg0 <= 36'sb100100101111001100001000111100011000;
            sine_reg0   <= 36'sb101111001111101001011010000110111000;
        end
        9630: begin
            cosine_reg0 <= 36'sb100100101111100110011101111010101100;
            sine_reg0   <= 36'sb101111001110111110100101101100000110;
        end
        9631: begin
            cosine_reg0 <= 36'sb100100110000000000110011111100010000;
            sine_reg0   <= 36'sb101111001110010011110001111010101011;
        end
        9632: begin
            cosine_reg0 <= 36'sb100100110000011011001011000001000100;
            sine_reg0   <= 36'sb101111001101101000111110110010101001;
        end
        9633: begin
            cosine_reg0 <= 36'sb100100110000110101100011001001000101;
            sine_reg0   <= 36'sb101111001100111110001100010100000010;
        end
        9634: begin
            cosine_reg0 <= 36'sb100100110001001111111100010100010011;
            sine_reg0   <= 36'sb101111001100010011011010011110111000;
        end
        9635: begin
            cosine_reg0 <= 36'sb100100110001101010010110100010101110;
            sine_reg0   <= 36'sb101111001011101000101001010011001100;
        end
        9636: begin
            cosine_reg0 <= 36'sb100100110010000100110001110100010100;
            sine_reg0   <= 36'sb101111001010111101111000110001000000;
        end
        9637: begin
            cosine_reg0 <= 36'sb100100110010011111001110001001000011;
            sine_reg0   <= 36'sb101111001010010011001000111000010101;
        end
        9638: begin
            cosine_reg0 <= 36'sb100100110010111001101011100000111100;
            sine_reg0   <= 36'sb101111001001101000011001101001001101;
        end
        9639: begin
            cosine_reg0 <= 36'sb100100110011010100001001111011111100;
            sine_reg0   <= 36'sb101111001000111101101011000011101010;
        end
        9640: begin
            cosine_reg0 <= 36'sb100100110011101110101001011010000100;
            sine_reg0   <= 36'sb101111001000010010111101000111101110;
        end
        9641: begin
            cosine_reg0 <= 36'sb100100110100001001001001111011010010;
            sine_reg0   <= 36'sb101111000111101000001111110101011001;
        end
        9642: begin
            cosine_reg0 <= 36'sb100100110100100011101011011111100100;
            sine_reg0   <= 36'sb101111000110111101100011001100101110;
        end
        9643: begin
            cosine_reg0 <= 36'sb100100110100111110001110000110111010;
            sine_reg0   <= 36'sb101111000110010010110111001101101111;
        end
        9644: begin
            cosine_reg0 <= 36'sb100100110101011000110001110001010100;
            sine_reg0   <= 36'sb101111000101101000001011111000011101;
        end
        9645: begin
            cosine_reg0 <= 36'sb100100110101110011010110011110101111;
            sine_reg0   <= 36'sb101111000100111101100001001100111001;
        end
        9646: begin
            cosine_reg0 <= 36'sb100100110110001101111100001111001011;
            sine_reg0   <= 36'sb101111000100010010110111001011000101;
        end
        9647: begin
            cosine_reg0 <= 36'sb100100110110101000100011000010100110;
            sine_reg0   <= 36'sb101111000011101000001101110011000100;
        end
        9648: begin
            cosine_reg0 <= 36'sb100100110111000011001010111001000001;
            sine_reg0   <= 36'sb101111000010111101100101000100110110;
        end
        9649: begin
            cosine_reg0 <= 36'sb100100110111011101110011110010011001;
            sine_reg0   <= 36'sb101111000010010010111101000000011101;
        end
        9650: begin
            cosine_reg0 <= 36'sb100100110111111000011101101110101110;
            sine_reg0   <= 36'sb101111000001101000010101100101111011;
        end
        9651: begin
            cosine_reg0 <= 36'sb100100111000010011001000101101111111;
            sine_reg0   <= 36'sb101111000000111101101110110101010010;
        end
        9652: begin
            cosine_reg0 <= 36'sb100100111000101101110100110000001010;
            sine_reg0   <= 36'sb101111000000010011001000101110100011;
        end
        9653: begin
            cosine_reg0 <= 36'sb100100111001001000100001110101001111;
            sine_reg0   <= 36'sb101110111111101000100011010001101111;
        end
        9654: begin
            cosine_reg0 <= 36'sb100100111001100011001111111101001101;
            sine_reg0   <= 36'sb101110111110111101111110011110111001;
        end
        9655: begin
            cosine_reg0 <= 36'sb100100111001111101111111001000000010;
            sine_reg0   <= 36'sb101110111110010011011010010110000011;
        end
        9656: begin
            cosine_reg0 <= 36'sb100100111010011000101111010101101110;
            sine_reg0   <= 36'sb101110111101101000110110110111001100;
        end
        9657: begin
            cosine_reg0 <= 36'sb100100111010110011100000100110001111;
            sine_reg0   <= 36'sb101110111100111110010100000010011001;
        end
        9658: begin
            cosine_reg0 <= 36'sb100100111011001110010010111001100101;
            sine_reg0   <= 36'sb101110111100010011110001110111101001;
        end
        9659: begin
            cosine_reg0 <= 36'sb100100111011101001000110001111101110;
            sine_reg0   <= 36'sb101110111011101001010000010110111111;
        end
        9660: begin
            cosine_reg0 <= 36'sb100100111100000011111010101000101010;
            sine_reg0   <= 36'sb101110111010111110101111100000011100;
        end
        9661: begin
            cosine_reg0 <= 36'sb100100111100011110110000000100010111;
            sine_reg0   <= 36'sb101110111010010100001111010100000010;
        end
        9662: begin
            cosine_reg0 <= 36'sb100100111100111001100110100010110100;
            sine_reg0   <= 36'sb101110111001101001101111110001110010;
        end
        9663: begin
            cosine_reg0 <= 36'sb100100111101010100011110000100000001;
            sine_reg0   <= 36'sb101110111000111111010000111001101111;
        end
        9664: begin
            cosine_reg0 <= 36'sb100100111101101111010110100111111100;
            sine_reg0   <= 36'sb101110111000010100110010101011111010;
        end
        9665: begin
            cosine_reg0 <= 36'sb100100111110001010010000001110100100;
            sine_reg0   <= 36'sb101110110111101010010101001000010100;
        end
        9666: begin
            cosine_reg0 <= 36'sb100100111110100101001010110111111000;
            sine_reg0   <= 36'sb101110110110111111111000001110111111;
        end
        9667: begin
            cosine_reg0 <= 36'sb100100111111000000000110100011111000;
            sine_reg0   <= 36'sb101110110110010101011011111111111101;
        end
        9668: begin
            cosine_reg0 <= 36'sb100100111111011011000011010010100010;
            sine_reg0   <= 36'sb101110110101101011000000011011001111;
        end
        9669: begin
            cosine_reg0 <= 36'sb100100111111110110000001000011110100;
            sine_reg0   <= 36'sb101110110101000000100101100000111000;
        end
        9670: begin
            cosine_reg0 <= 36'sb100101000000010000111111110111101111;
            sine_reg0   <= 36'sb101110110100010110001011010000111000;
        end
        9671: begin
            cosine_reg0 <= 36'sb100101000000101011111111101110010001;
            sine_reg0   <= 36'sb101110110011101011110001101011010001;
        end
        9672: begin
            cosine_reg0 <= 36'sb100101000001000111000000100111011001;
            sine_reg0   <= 36'sb101110110011000001011000110000000101;
        end
        9673: begin
            cosine_reg0 <= 36'sb100101000001100010000010100011000110;
            sine_reg0   <= 36'sb101110110010010111000000011111010110;
        end
        9674: begin
            cosine_reg0 <= 36'sb100101000001111101000101100001010110;
            sine_reg0   <= 36'sb101110110001101100101000111001000101;
        end
        9675: begin
            cosine_reg0 <= 36'sb100101000010011000001001100010001010;
            sine_reg0   <= 36'sb101110110001000010010001111101010011;
        end
        9676: begin
            cosine_reg0 <= 36'sb100101000010110011001110100101011111;
            sine_reg0   <= 36'sb101110110000010111111011101100000100;
        end
        9677: begin
            cosine_reg0 <= 36'sb100101000011001110010100101011010101;
            sine_reg0   <= 36'sb101110101111101101100110000101010111;
        end
        9678: begin
            cosine_reg0 <= 36'sb100101000011101001011011110011101011;
            sine_reg0   <= 36'sb101110101111000011010001001001001111;
        end
        9679: begin
            cosine_reg0 <= 36'sb100101000100000100100011111110100000;
            sine_reg0   <= 36'sb101110101110011000111100110111101101;
        end
        9680: begin
            cosine_reg0 <= 36'sb100101000100011111101101001011110010;
            sine_reg0   <= 36'sb101110101101101110101001010000110100;
        end
        9681: begin
            cosine_reg0 <= 36'sb100101000100111010110111011011100000;
            sine_reg0   <= 36'sb101110101101000100010110010100100100;
        end
        9682: begin
            cosine_reg0 <= 36'sb100101000101010110000010101101101011;
            sine_reg0   <= 36'sb101110101100011010000100000010111111;
        end
        9683: begin
            cosine_reg0 <= 36'sb100101000101110001001111000010001111;
            sine_reg0   <= 36'sb101110101011101111110010011100000111;
        end
        9684: begin
            cosine_reg0 <= 36'sb100101000110001100011100011001001110;
            sine_reg0   <= 36'sb101110101011000101100001011111111110;
        end
        9685: begin
            cosine_reg0 <= 36'sb100101000110100111101010110010100100;
            sine_reg0   <= 36'sb101110101010011011010001001110100100;
        end
        9686: begin
            cosine_reg0 <= 36'sb100101000111000010111010001110010010;
            sine_reg0   <= 36'sb101110101001110001000001100111111101;
        end
        9687: begin
            cosine_reg0 <= 36'sb100101000111011110001010101100010110;
            sine_reg0   <= 36'sb101110101001000110110010101100001001;
        end
        9688: begin
            cosine_reg0 <= 36'sb100101000111111001011100001100101111;
            sine_reg0   <= 36'sb101110101000011100100100011011001010;
        end
        9689: begin
            cosine_reg0 <= 36'sb100101001000010100101110101111011101;
            sine_reg0   <= 36'sb101110100111110010010110110101000001;
        end
        9690: begin
            cosine_reg0 <= 36'sb100101001000110000000010010100011110;
            sine_reg0   <= 36'sb101110100111001000001001111001110001;
        end
        9691: begin
            cosine_reg0 <= 36'sb100101001001001011010110111011110000;
            sine_reg0   <= 36'sb101110100110011101111101101001011011;
        end
        9692: begin
            cosine_reg0 <= 36'sb100101001001100110101100100101010100;
            sine_reg0   <= 36'sb101110100101110011110010000100000000;
        end
        9693: begin
            cosine_reg0 <= 36'sb100101001010000010000011010001001000;
            sine_reg0   <= 36'sb101110100101001001100111001001100010;
        end
        9694: begin
            cosine_reg0 <= 36'sb100101001010011101011010111111001011;
            sine_reg0   <= 36'sb101110100100011111011100111010000100;
        end
        9695: begin
            cosine_reg0 <= 36'sb100101001010111000110011101111011011;
            sine_reg0   <= 36'sb101110100011110101010011010101100101;
        end
        9696: begin
            cosine_reg0 <= 36'sb100101001011010100001101100001111000;
            sine_reg0   <= 36'sb101110100011001011001010011100001001;
        end
        9697: begin
            cosine_reg0 <= 36'sb100101001011101111101000010110100001;
            sine_reg0   <= 36'sb101110100010100001000010001101110000;
        end
        9698: begin
            cosine_reg0 <= 36'sb100101001100001011000100001101010101;
            sine_reg0   <= 36'sb101110100001110110111010101010011101;
        end
        9699: begin
            cosine_reg0 <= 36'sb100101001100100110100001000110010011;
            sine_reg0   <= 36'sb101110100001001100110011110010010000;
        end
        9700: begin
            cosine_reg0 <= 36'sb100101001101000001111111000001011001;
            sine_reg0   <= 36'sb101110100000100010101101100101001100;
        end
        9701: begin
            cosine_reg0 <= 36'sb100101001101011101011101111110100110;
            sine_reg0   <= 36'sb101110011111111000101000000011010010;
        end
        9702: begin
            cosine_reg0 <= 36'sb100101001101111000111101111101111010;
            sine_reg0   <= 36'sb101110011111001110100011001100100100;
        end
        9703: begin
            cosine_reg0 <= 36'sb100101001110010100011110111111010011;
            sine_reg0   <= 36'sb101110011110100100011111000001000100;
        end
        9704: begin
            cosine_reg0 <= 36'sb100101001110110000000001000010110001;
            sine_reg0   <= 36'sb101110011101111010011011100000110010;
        end
        9705: begin
            cosine_reg0 <= 36'sb100101001111001011100100001000010010;
            sine_reg0   <= 36'sb101110011101010000011000101011110001;
        end
        9706: begin
            cosine_reg0 <= 36'sb100101001111100111001000001111110101;
            sine_reg0   <= 36'sb101110011100100110010110100010000010;
        end
        9707: begin
            cosine_reg0 <= 36'sb100101010000000010101101011001011010;
            sine_reg0   <= 36'sb101110011011111100010101000011100111;
        end
        9708: begin
            cosine_reg0 <= 36'sb100101010000011110010011100100111110;
            sine_reg0   <= 36'sb101110011011010010010100010000100010;
        end
        9709: begin
            cosine_reg0 <= 36'sb100101010000111001111010110010100001;
            sine_reg0   <= 36'sb101110011010101000010100001000110100;
        end
        9710: begin
            cosine_reg0 <= 36'sb100101010001010101100011000010000011;
            sine_reg0   <= 36'sb101110011001111110010100101100011110;
        end
        9711: begin
            cosine_reg0 <= 36'sb100101010001110001001100010011100001;
            sine_reg0   <= 36'sb101110011001010100010101111011100011;
        end
        9712: begin
            cosine_reg0 <= 36'sb100101010010001100110110100110111011;
            sine_reg0   <= 36'sb101110011000101010010111110110000100;
        end
        9713: begin
            cosine_reg0 <= 36'sb100101010010101000100001111100010000;
            sine_reg0   <= 36'sb101110011000000000011010011100000010;
        end
        9714: begin
            cosine_reg0 <= 36'sb100101010011000100001110010011011111;
            sine_reg0   <= 36'sb101110010111010110011101101101100000;
        end
        9715: begin
            cosine_reg0 <= 36'sb100101010011011111111011101100100110;
            sine_reg0   <= 36'sb101110010110101100100001101010011110;
        end
        9716: begin
            cosine_reg0 <= 36'sb100101010011111011101010000111100100;
            sine_reg0   <= 36'sb101110010110000010100110010010111111;
        end
        9717: begin
            cosine_reg0 <= 36'sb100101010100010111011001100100011010;
            sine_reg0   <= 36'sb101110010101011000101011100111000100;
        end
        9718: begin
            cosine_reg0 <= 36'sb100101010100110011001010000011000100;
            sine_reg0   <= 36'sb101110010100101110110001100110101111;
        end
        9719: begin
            cosine_reg0 <= 36'sb100101010101001110111011100011100011;
            sine_reg0   <= 36'sb101110010100000100111000010010000001;
        end
        9720: begin
            cosine_reg0 <= 36'sb100101010101101010101110000101110110;
            sine_reg0   <= 36'sb101110010011011010111111101000111100;
        end
        9721: begin
            cosine_reg0 <= 36'sb100101010110000110100001101001111010;
            sine_reg0   <= 36'sb101110010010110001000111101011100001;
        end
        9722: begin
            cosine_reg0 <= 36'sb100101010110100010010110001111110000;
            sine_reg0   <= 36'sb101110010010000111010000011001110011;
        end
        9723: begin
            cosine_reg0 <= 36'sb100101010110111110001011110111010101;
            sine_reg0   <= 36'sb101110010001011101011001110011110010;
        end
        9724: begin
            cosine_reg0 <= 36'sb100101010111011010000010100000101010;
            sine_reg0   <= 36'sb101110010000110011100011111001100000;
        end
        9725: begin
            cosine_reg0 <= 36'sb100101010111110101111010001011101101;
            sine_reg0   <= 36'sb101110010000001001101110101011000000;
        end
        9726: begin
            cosine_reg0 <= 36'sb100101011000010001110010111000011100;
            sine_reg0   <= 36'sb101110001111011111111010001000010010;
        end
        9727: begin
            cosine_reg0 <= 36'sb100101011000101101101100100110110111;
            sine_reg0   <= 36'sb101110001110110110000110010001011001;
        end
        9728: begin
            cosine_reg0 <= 36'sb100101011001001001100111010110111101;
            sine_reg0   <= 36'sb101110001110001100010011000110010101;
        end
        9729: begin
            cosine_reg0 <= 36'sb100101011001100101100011001000101101;
            sine_reg0   <= 36'sb101110001101100010100000100111001001;
        end
        9730: begin
            cosine_reg0 <= 36'sb100101011010000001011111111100000101;
            sine_reg0   <= 36'sb101110001100111000101110110011110101;
        end
        9731: begin
            cosine_reg0 <= 36'sb100101011010011101011101110001000100;
            sine_reg0   <= 36'sb101110001100001110111101101100011101;
        end
        9732: begin
            cosine_reg0 <= 36'sb100101011010111001011100100111101010;
            sine_reg0   <= 36'sb101110001011100101001101010001000000;
        end
        9733: begin
            cosine_reg0 <= 36'sb100101011011010101011100011111110101;
            sine_reg0   <= 36'sb101110001010111011011101100001100010;
        end
        9734: begin
            cosine_reg0 <= 36'sb100101011011110001011101011001100101;
            sine_reg0   <= 36'sb101110001010010001101110011110000011;
        end
        9735: begin
            cosine_reg0 <= 36'sb100101011100001101011111010100110111;
            sine_reg0   <= 36'sb101110001001101000000000000110100101;
        end
        9736: begin
            cosine_reg0 <= 36'sb100101011100101001100010010001101100;
            sine_reg0   <= 36'sb101110001000111110010010011011001001;
        end
        9737: begin
            cosine_reg0 <= 36'sb100101011101000101100110010000000001;
            sine_reg0   <= 36'sb101110001000010100100101011011110011;
        end
        9738: begin
            cosine_reg0 <= 36'sb100101011101100001101011001111110111;
            sine_reg0   <= 36'sb101110000111101010111001001000100001;
        end
        9739: begin
            cosine_reg0 <= 36'sb100101011101111101110001010001001011;
            sine_reg0   <= 36'sb101110000111000001001101100001011000;
        end
        9740: begin
            cosine_reg0 <= 36'sb100101011110011001111000010011111101;
            sine_reg0   <= 36'sb101110000110010111100010100110011000;
        end
        9741: begin
            cosine_reg0 <= 36'sb100101011110110110000000011000001100;
            sine_reg0   <= 36'sb101110000101101101111000010111100010;
        end
        9742: begin
            cosine_reg0 <= 36'sb100101011111010010001001011101110110;
            sine_reg0   <= 36'sb101110000101000100001110110100111001;
        end
        9743: begin
            cosine_reg0 <= 36'sb100101011111101110010011100100111011;
            sine_reg0   <= 36'sb101110000100011010100101111110011101;
        end
        9744: begin
            cosine_reg0 <= 36'sb100101100000001010011110101101011001;
            sine_reg0   <= 36'sb101110000011110000111101110100010001;
        end
        9745: begin
            cosine_reg0 <= 36'sb100101100000100110101010110111001111;
            sine_reg0   <= 36'sb101110000011000111010110010110010111;
        end
        9746: begin
            cosine_reg0 <= 36'sb100101100001000010111000000010011101;
            sine_reg0   <= 36'sb101110000010011101101111100100101111;
        end
        9747: begin
            cosine_reg0 <= 36'sb100101100001011111000110001111000001;
            sine_reg0   <= 36'sb101110000001110100001001011111011011;
        end
        9748: begin
            cosine_reg0 <= 36'sb100101100001111011010101011100111010;
            sine_reg0   <= 36'sb101110000001001010100100000110011110;
        end
        9749: begin
            cosine_reg0 <= 36'sb100101100010010111100101101100000110;
            sine_reg0   <= 36'sb101110000000100000111111011001111000;
        end
        9750: begin
            cosine_reg0 <= 36'sb100101100010110011110110111100100110;
            sine_reg0   <= 36'sb101101111111110111011011011001101011;
        end
        9751: begin
            cosine_reg0 <= 36'sb100101100011010000001001001110010111;
            sine_reg0   <= 36'sb101101111111001101111000000101111001;
        end
        9752: begin
            cosine_reg0 <= 36'sb100101100011101100011100100001011001;
            sine_reg0   <= 36'sb101101111110100100010101011110100011;
        end
        9753: begin
            cosine_reg0 <= 36'sb100101100100001000110000110101101011;
            sine_reg0   <= 36'sb101101111101111010110011100011101100;
        end
        9754: begin
            cosine_reg0 <= 36'sb100101100100100101000110001011001011;
            sine_reg0   <= 36'sb101101111101010001010010010101010011;
        end
        9755: begin
            cosine_reg0 <= 36'sb100101100101000001011100100001111001;
            sine_reg0   <= 36'sb101101111100100111110001110011011100;
        end
        9756: begin
            cosine_reg0 <= 36'sb100101100101011101110011111001110011;
            sine_reg0   <= 36'sb101101111011111110010001111110001000;
        end
        9757: begin
            cosine_reg0 <= 36'sb100101100101111010001100010010111000;
            sine_reg0   <= 36'sb101101111011010100110010110101011001;
        end
        9758: begin
            cosine_reg0 <= 36'sb100101100110010110100101101101000111;
            sine_reg0   <= 36'sb101101111010101011010100011001001111;
        end
        9759: begin
            cosine_reg0 <= 36'sb100101100110110011000000001000100000;
            sine_reg0   <= 36'sb101101111010000001110110101001101101;
        end
        9760: begin
            cosine_reg0 <= 36'sb100101100111001111011011100101000000;
            sine_reg0   <= 36'sb101101111001011000011001100110110100;
        end
        9761: begin
            cosine_reg0 <= 36'sb100101100111101011111000000010100111;
            sine_reg0   <= 36'sb101101111000101110111101010000100101;
        end
        9762: begin
            cosine_reg0 <= 36'sb100101101000001000010101100001010100;
            sine_reg0   <= 36'sb101101111000000101100001100111000011;
        end
        9763: begin
            cosine_reg0 <= 36'sb100101101000100100110100000001000110;
            sine_reg0   <= 36'sb101101110111011100000110101010010000;
        end
        9764: begin
            cosine_reg0 <= 36'sb100101101001000001010011100001111011;
            sine_reg0   <= 36'sb101101110110110010101100011010001011;
        end
        9765: begin
            cosine_reg0 <= 36'sb100101101001011101110100000011110010;
            sine_reg0   <= 36'sb101101110110001001010010110110111000;
        end
        9766: begin
            cosine_reg0 <= 36'sb100101101001111010010101100110101011;
            sine_reg0   <= 36'sb101101110101011111111010000000011000;
        end
        9767: begin
            cosine_reg0 <= 36'sb100101101010010110111000001010100100;
            sine_reg0   <= 36'sb101101110100110110100001110110101100;
        end
        9768: begin
            cosine_reg0 <= 36'sb100101101010110011011011101111011101;
            sine_reg0   <= 36'sb101101110100001101001010011001110110;
        end
        9769: begin
            cosine_reg0 <= 36'sb100101101011010000000000010101010011;
            sine_reg0   <= 36'sb101101110011100011110011101001110111;
        end
        9770: begin
            cosine_reg0 <= 36'sb100101101011101100100101111100000110;
            sine_reg0   <= 36'sb101101110010111010011101100110110010;
        end
        9771: begin
            cosine_reg0 <= 36'sb100101101100001001001100100011110101;
            sine_reg0   <= 36'sb101101110010010001001000010000100111;
        end
        9772: begin
            cosine_reg0 <= 36'sb100101101100100101110100001100011111;
            sine_reg0   <= 36'sb101101110001100111110011100111011001;
        end
        9773: begin
            cosine_reg0 <= 36'sb100101101101000010011100110110000011;
            sine_reg0   <= 36'sb101101110000111110011111101011001000;
        end
        9774: begin
            cosine_reg0 <= 36'sb100101101101011111000110100000011111;
            sine_reg0   <= 36'sb101101110000010101001100011011110111;
        end
        9775: begin
            cosine_reg0 <= 36'sb100101101101111011110001001011110011;
            sine_reg0   <= 36'sb101101101111101011111001111001100111;
        end
        9776: begin
            cosine_reg0 <= 36'sb100101101110011000011100110111111100;
            sine_reg0   <= 36'sb101101101111000010101000000100011010;
        end
        9777: begin
            cosine_reg0 <= 36'sb100101101110110101001001100100111100;
            sine_reg0   <= 36'sb101101101110011001010110111100010010;
        end
        9778: begin
            cosine_reg0 <= 36'sb100101101111010001110111010010101111;
            sine_reg0   <= 36'sb101101101101110000000110100001001111;
        end
        9779: begin
            cosine_reg0 <= 36'sb100101101111101110100110000001010101;
            sine_reg0   <= 36'sb101101101101000110110110110011010011;
        end
        9780: begin
            cosine_reg0 <= 36'sb100101110000001011010101110000101101;
            sine_reg0   <= 36'sb101101101100011101100111110010100001;
        end
        9781: begin
            cosine_reg0 <= 36'sb100101110000101000000110100000110110;
            sine_reg0   <= 36'sb101101101011110100011001011110111001;
        end
        9782: begin
            cosine_reg0 <= 36'sb100101110001000100111000010001101111;
            sine_reg0   <= 36'sb101101101011001011001011111000011110;
        end
        9783: begin
            cosine_reg0 <= 36'sb100101110001100001101011000011010110;
            sine_reg0   <= 36'sb101101101010100001111110111111010000;
        end
        9784: begin
            cosine_reg0 <= 36'sb100101110001111110011110110101101011;
            sine_reg0   <= 36'sb101101101001111000110010110011010010;
        end
        9785: begin
            cosine_reg0 <= 36'sb100101110010011011010011101000101100;
            sine_reg0   <= 36'sb101101101001001111100111010100100100;
        end
        9786: begin
            cosine_reg0 <= 36'sb100101110010111000001001011100011000;
            sine_reg0   <= 36'sb101101101000100110011100100011001010;
        end
        9787: begin
            cosine_reg0 <= 36'sb100101110011010101000000010000101110;
            sine_reg0   <= 36'sb101101100111111101010010011111000011;
        end
        9788: begin
            cosine_reg0 <= 36'sb100101110011110001111000000101101110;
            sine_reg0   <= 36'sb101101100111010100001001001000010011;
        end
        9789: begin
            cosine_reg0 <= 36'sb100101110100001110110000111011010101;
            sine_reg0   <= 36'sb101101100110101011000000011110111001;
        end
        9790: begin
            cosine_reg0 <= 36'sb100101110100101011101010110001100011;
            sine_reg0   <= 36'sb101101100110000001111000100010111001;
        end
        9791: begin
            cosine_reg0 <= 36'sb100101110101001000100101101000010111;
            sine_reg0   <= 36'sb101101100101011000110001010100010011;
        end
        9792: begin
            cosine_reg0 <= 36'sb100101110101100101100001011111101111;
            sine_reg0   <= 36'sb101101100100101111101010110011001001;
        end
        9793: begin
            cosine_reg0 <= 36'sb100101110110000010011110010111101011;
            sine_reg0   <= 36'sb101101100100000110100100111111011101;
        end
        9794: begin
            cosine_reg0 <= 36'sb100101110110011111011100010000001001;
            sine_reg0   <= 36'sb101101100011011101011111111001010000;
        end
        9795: begin
            cosine_reg0 <= 36'sb100101110110111100011011001001001001;
            sine_reg0   <= 36'sb101101100010110100011011100000100101;
        end
        9796: begin
            cosine_reg0 <= 36'sb100101110111011001011011000010101000;
            sine_reg0   <= 36'sb101101100010001011010111110101011011;
        end
        9797: begin
            cosine_reg0 <= 36'sb100101110111110110011011111100100111;
            sine_reg0   <= 36'sb101101100001100010010100110111110110;
        end
        9798: begin
            cosine_reg0 <= 36'sb100101111000010011011101110111000011;
            sine_reg0   <= 36'sb101101100000111001010010100111110110;
        end
        9799: begin
            cosine_reg0 <= 36'sb100101111000110000100000110001111100;
            sine_reg0   <= 36'sb101101100000010000010001000101011101;
        end
        9800: begin
            cosine_reg0 <= 36'sb100101111001001101100100101101010001;
            sine_reg0   <= 36'sb101101011111100111010000010000101101;
        end
        9801: begin
            cosine_reg0 <= 36'sb100101111001101010101001101001000000;
            sine_reg0   <= 36'sb101101011110111110010000001001101000;
        end
        9802: begin
            cosine_reg0 <= 36'sb100101111010000111101111100101001000;
            sine_reg0   <= 36'sb101101011110010101010000110000001110;
        end
        9803: begin
            cosine_reg0 <= 36'sb100101111010100100110110100001101001;
            sine_reg0   <= 36'sb101101011101101100010010000100100010;
        end
        9804: begin
            cosine_reg0 <= 36'sb100101111011000001111110011110100001;
            sine_reg0   <= 36'sb101101011101000011010100000110100101;
        end
        9805: begin
            cosine_reg0 <= 36'sb100101111011011111000111011011101111;
            sine_reg0   <= 36'sb101101011100011010010110110110011001;
        end
        9806: begin
            cosine_reg0 <= 36'sb100101111011111100010001011001010010;
            sine_reg0   <= 36'sb101101011011110001011010010011111111;
        end
        9807: begin
            cosine_reg0 <= 36'sb100101111100011001011100010111001001;
            sine_reg0   <= 36'sb101101011011001000011110011111011001;
        end
        9808: begin
            cosine_reg0 <= 36'sb100101111100110110101000010101010010;
            sine_reg0   <= 36'sb101101011010011111100011011000101000;
        end
        9809: begin
            cosine_reg0 <= 36'sb100101111101010011110101010011101101;
            sine_reg0   <= 36'sb101101011001110110101000111111101110;
        end
        9810: begin
            cosine_reg0 <= 36'sb100101111101110001000011010010011000;
            sine_reg0   <= 36'sb101101011001001101101111010100101101;
        end
        9811: begin
            cosine_reg0 <= 36'sb100101111110001110010010010001010011;
            sine_reg0   <= 36'sb101101011000100100110110010111100110;
        end
        9812: begin
            cosine_reg0 <= 36'sb100101111110101011100010010000011011;
            sine_reg0   <= 36'sb101101010111111011111110001000011011;
        end
        9813: begin
            cosine_reg0 <= 36'sb100101111111001000110011001111110001;
            sine_reg0   <= 36'sb101101010111010011000110100111001100;
        end
        9814: begin
            cosine_reg0 <= 36'sb100101111111100110000101001111010010;
            sine_reg0   <= 36'sb101101010110101010001111110011111101;
        end
        9815: begin
            cosine_reg0 <= 36'sb100110000000000011011000001110111111;
            sine_reg0   <= 36'sb101101010110000001011001101110101111;
        end
        9816: begin
            cosine_reg0 <= 36'sb100110000000100000101100001110110100;
            sine_reg0   <= 36'sb101101010101011000100100010111100010;
        end
        9817: begin
            cosine_reg0 <= 36'sb100110000000111110000001001110110011;
            sine_reg0   <= 36'sb101101010100101111101111101110011001;
        end
        9818: begin
            cosine_reg0 <= 36'sb100110000001011011010111001110111001;
            sine_reg0   <= 36'sb101101010100000110111011110011010101;
        end
        9819: begin
            cosine_reg0 <= 36'sb100110000001111000101110001111000101;
            sine_reg0   <= 36'sb101101010011011110001000100110011000;
        end
        9820: begin
            cosine_reg0 <= 36'sb100110000010010110000110001111010110;
            sine_reg0   <= 36'sb101101010010110101010110000111100011;
        end
        9821: begin
            cosine_reg0 <= 36'sb100110000010110011011111001111101011;
            sine_reg0   <= 36'sb101101010010001100100100010110111000;
        end
        9822: begin
            cosine_reg0 <= 36'sb100110000011010000111001010000000011;
            sine_reg0   <= 36'sb101101010001100011110011010100011000;
        end
        9823: begin
            cosine_reg0 <= 36'sb100110000011101110010100010000011100;
            sine_reg0   <= 36'sb101101010000111011000011000000000110;
        end
        9824: begin
            cosine_reg0 <= 36'sb100110000100001011110000010000110110;
            sine_reg0   <= 36'sb101101010000010010010011011010000010;
        end
        9825: begin
            cosine_reg0 <= 36'sb100110000100101001001101010001010000;
            sine_reg0   <= 36'sb101101001111101001100100100010001110;
        end
        9826: begin
            cosine_reg0 <= 36'sb100110000101000110101011010001101000;
            sine_reg0   <= 36'sb101101001111000000110110011000101100;
        end
        9827: begin
            cosine_reg0 <= 36'sb100110000101100100001010010001111101;
            sine_reg0   <= 36'sb101101001110011000001000111101011110;
        end
        9828: begin
            cosine_reg0 <= 36'sb100110000110000001101010010010001110;
            sine_reg0   <= 36'sb101101001101101111011100010000100100;
        end
        9829: begin
            cosine_reg0 <= 36'sb100110000110011111001011010010011010;
            sine_reg0   <= 36'sb101101001101000110110000010010000000;
        end
        9830: begin
            cosine_reg0 <= 36'sb100110000110111100101101010010100000;
            sine_reg0   <= 36'sb101101001100011110000101000001110101;
        end
        9831: begin
            cosine_reg0 <= 36'sb100110000111011010010000010010011110;
            sine_reg0   <= 36'sb101101001011110101011010100000000011;
        end
        9832: begin
            cosine_reg0 <= 36'sb100110000111110111110100010010010100;
            sine_reg0   <= 36'sb101101001011001100110000101100101101;
        end
        9833: begin
            cosine_reg0 <= 36'sb100110001000010101011001010010000000;
            sine_reg0   <= 36'sb101101001010100100000111100111110011;
        end
        9834: begin
            cosine_reg0 <= 36'sb100110001000110010111111010001100001;
            sine_reg0   <= 36'sb101101001001111011011111010001011000;
        end
        9835: begin
            cosine_reg0 <= 36'sb100110001001010000100110010000110111;
            sine_reg0   <= 36'sb101101001001010010110111101001011100;
        end
        9836: begin
            cosine_reg0 <= 36'sb100110001001101110001110001111111111;
            sine_reg0   <= 36'sb101101001000101010010000110000000010;
        end
        9837: begin
            cosine_reg0 <= 36'sb100110001010001011110111001110111001;
            sine_reg0   <= 36'sb101101001000000001101010100101001010;
        end
        9838: begin
            cosine_reg0 <= 36'sb100110001010101001100001001101100100;
            sine_reg0   <= 36'sb101101000111011001000101001000111000;
        end
        9839: begin
            cosine_reg0 <= 36'sb100110001011000111001100001011111110;
            sine_reg0   <= 36'sb101101000110110000100000011011001011;
        end
        9840: begin
            cosine_reg0 <= 36'sb100110001011100100111000001010000110;
            sine_reg0   <= 36'sb101101000110000111111100011100000110;
        end
        9841: begin
            cosine_reg0 <= 36'sb100110001100000010100101000111111100;
            sine_reg0   <= 36'sb101101000101011111011001001011101011;
        end
        9842: begin
            cosine_reg0 <= 36'sb100110001100100000010011000101011110;
            sine_reg0   <= 36'sb101101000100110110110110101001111010;
        end
        9843: begin
            cosine_reg0 <= 36'sb100110001100111110000010000010101010;
            sine_reg0   <= 36'sb101101000100001110010100110110110101;
        end
        9844: begin
            cosine_reg0 <= 36'sb100110001101011011110001111111100001;
            sine_reg0   <= 36'sb101101000011100101110011110010011111;
        end
        9845: begin
            cosine_reg0 <= 36'sb100110001101111001100010111100000000;
            sine_reg0   <= 36'sb101101000010111101010011011100111000;
        end
        9846: begin
            cosine_reg0 <= 36'sb100110001110010111010100111000000110;
            sine_reg0   <= 36'sb101101000010010100110011110110000010;
        end
        9847: begin
            cosine_reg0 <= 36'sb100110001110110101000111110011110011;
            sine_reg0   <= 36'sb101101000001101100010100111101111111;
        end
        9848: begin
            cosine_reg0 <= 36'sb100110001111010010111011101111000101;
            sine_reg0   <= 36'sb101101000001000011110110110100110000;
        end
        9849: begin
            cosine_reg0 <= 36'sb100110001111110000110000101001111011;
            sine_reg0   <= 36'sb101101000000011011011001011010010110;
        end
        9850: begin
            cosine_reg0 <= 36'sb100110010000001110100110100100010011;
            sine_reg0   <= 36'sb101100111111110010111100101110110100;
        end
        9851: begin
            cosine_reg0 <= 36'sb100110010000101100011101011110001110;
            sine_reg0   <= 36'sb101100111111001010100000110010001011;
        end
        9852: begin
            cosine_reg0 <= 36'sb100110010001001010010101010111101001;
            sine_reg0   <= 36'sb101100111110100010000101100100011100;
        end
        9853: begin
            cosine_reg0 <= 36'sb100110010001101000001110010000100100;
            sine_reg0   <= 36'sb101100111101111001101011000101101001;
        end
        9854: begin
            cosine_reg0 <= 36'sb100110010010000110001000001000111100;
            sine_reg0   <= 36'sb101100111101010001010001010101110100;
        end
        9855: begin
            cosine_reg0 <= 36'sb100110010010100100000011000000110010;
            sine_reg0   <= 36'sb101100111100101000111000010100111110;
        end
        9856: begin
            cosine_reg0 <= 36'sb100110010011000001111110111000000100;
            sine_reg0   <= 36'sb101100111100000000100000000011001000;
        end
        9857: begin
            cosine_reg0 <= 36'sb100110010011011111111011101110110001;
            sine_reg0   <= 36'sb101100111011011000001000100000010101;
        end
        9858: begin
            cosine_reg0 <= 36'sb100110010011111101111001100100110111;
            sine_reg0   <= 36'sb101100111010101111110001101100100101;
        end
        9859: begin
            cosine_reg0 <= 36'sb100110010100011011111000011010010110;
            sine_reg0   <= 36'sb101100111010000111011011100111111011;
        end
        9860: begin
            cosine_reg0 <= 36'sb100110010100111001111000001111001100;
            sine_reg0   <= 36'sb101100111001011111000110010010011000;
        end
        9861: begin
            cosine_reg0 <= 36'sb100110010101010111111001000011011000;
            sine_reg0   <= 36'sb101100111000110110110001101011111101;
        end
        9862: begin
            cosine_reg0 <= 36'sb100110010101110101111010110110111001;
            sine_reg0   <= 36'sb101100111000001110011101110100101100;
        end
        9863: begin
            cosine_reg0 <= 36'sb100110010110010011111101101001101110;
            sine_reg0   <= 36'sb101100110111100110001010101100100110;
        end
        9864: begin
            cosine_reg0 <= 36'sb100110010110110010000001011011110110;
            sine_reg0   <= 36'sb101100110110111101111000010011101110;
        end
        9865: begin
            cosine_reg0 <= 36'sb100110010111010000000110001101001111;
            sine_reg0   <= 36'sb101100110110010101100110101010000101;
        end
        9866: begin
            cosine_reg0 <= 36'sb100110010111101110001011111101111001;
            sine_reg0   <= 36'sb101100110101101101010101101111101011;
        end
        9867: begin
            cosine_reg0 <= 36'sb100110011000001100010010101101110010;
            sine_reg0   <= 36'sb101100110101000101000101100100100011;
        end
        9868: begin
            cosine_reg0 <= 36'sb100110011000101010011010011100111001;
            sine_reg0   <= 36'sb101100110100011100110110001000101111;
        end
        9869: begin
            cosine_reg0 <= 36'sb100110011001001000100011001011001101;
            sine_reg0   <= 36'sb101100110011110100100111011100001111;
        end
        9870: begin
            cosine_reg0 <= 36'sb100110011001100110101100111000101101;
            sine_reg0   <= 36'sb101100110011001100011001011111000110;
        end
        9871: begin
            cosine_reg0 <= 36'sb100110011010000100110111100101010111;
            sine_reg0   <= 36'sb101100110010100100001100010001010101;
        end
        9872: begin
            cosine_reg0 <= 36'sb100110011010100011000011010001001011;
            sine_reg0   <= 36'sb101100110001111011111111110010111101;
        end
        9873: begin
            cosine_reg0 <= 36'sb100110011011000001001111111100000111;
            sine_reg0   <= 36'sb101100110001010011110100000100000001;
        end
        9874: begin
            cosine_reg0 <= 36'sb100110011011011111011101100110001010;
            sine_reg0   <= 36'sb101100110000101011101001000100100001;
        end
        9875: begin
            cosine_reg0 <= 36'sb100110011011111101101100001111010011;
            sine_reg0   <= 36'sb101100110000000011011110110100011111;
        end
        9876: begin
            cosine_reg0 <= 36'sb100110011100011011111011110111100000;
            sine_reg0   <= 36'sb101100101111011011010101010011111101;
        end
        9877: begin
            cosine_reg0 <= 36'sb100110011100111010001100011110110010;
            sine_reg0   <= 36'sb101100101110110011001100100010111100;
        end
        9878: begin
            cosine_reg0 <= 36'sb100110011101011000011110000101000101;
            sine_reg0   <= 36'sb101100101110001011000100100001011110;
        end
        9879: begin
            cosine_reg0 <= 36'sb100110011101110110110000101010011010;
            sine_reg0   <= 36'sb101100101101100010111101001111100100;
        end
        9880: begin
            cosine_reg0 <= 36'sb100110011110010101000100001110101111;
            sine_reg0   <= 36'sb101100101100111010110110101101010000;
        end
        9881: begin
            cosine_reg0 <= 36'sb100110011110110011011000110010000011;
            sine_reg0   <= 36'sb101100101100010010110000111010100100;
        end
        9882: begin
            cosine_reg0 <= 36'sb100110011111010001101110010100010101;
            sine_reg0   <= 36'sb101100101011101010101011110111100000;
        end
        9883: begin
            cosine_reg0 <= 36'sb100110011111110000000100110101100011;
            sine_reg0   <= 36'sb101100101011000010100111100100001000;
        end
        9884: begin
            cosine_reg0 <= 36'sb100110100000001110011100010101101101;
            sine_reg0   <= 36'sb101100101010011010100100000000011011;
        end
        9885: begin
            cosine_reg0 <= 36'sb100110100000101100110100110100110001;
            sine_reg0   <= 36'sb101100101001110010100001001100011011;
        end
        9886: begin
            cosine_reg0 <= 36'sb100110100001001011001110010010101110;
            sine_reg0   <= 36'sb101100101001001010011111001000001011;
        end
        9887: begin
            cosine_reg0 <= 36'sb100110100001101001101000101111100011;
            sine_reg0   <= 36'sb101100101000100010011101110011101100;
        end
        9888: begin
            cosine_reg0 <= 36'sb100110100010001000000100001011001111;
            sine_reg0   <= 36'sb101100100111111010011101001110111111;
        end
        9889: begin
            cosine_reg0 <= 36'sb100110100010100110100000100101110000;
            sine_reg0   <= 36'sb101100100111010010011101011010000110;
        end
        9890: begin
            cosine_reg0 <= 36'sb100110100011000100111101111111000110;
            sine_reg0   <= 36'sb101100100110101010011110010101000010;
        end
        9891: begin
            cosine_reg0 <= 36'sb100110100011100011011100010111001110;
            sine_reg0   <= 36'sb101100100110000010011111111111110101;
        end
        9892: begin
            cosine_reg0 <= 36'sb100110100100000001111011101110001001;
            sine_reg0   <= 36'sb101100100101011010100010011010100000;
        end
        9893: begin
            cosine_reg0 <= 36'sb100110100100100000011100000011110101;
            sine_reg0   <= 36'sb101100100100110010100101100101000101;
        end
        9894: begin
            cosine_reg0 <= 36'sb100110100100111110111101011000010000;
            sine_reg0   <= 36'sb101100100100001010101001011111100110;
        end
        9895: begin
            cosine_reg0 <= 36'sb100110100101011101011111101011011010;
            sine_reg0   <= 36'sb101100100011100010101110001010000100;
        end
        9896: begin
            cosine_reg0 <= 36'sb100110100101111100000010111101010001;
            sine_reg0   <= 36'sb101100100010111010110011100100100000;
        end
        9897: begin
            cosine_reg0 <= 36'sb100110100110011010100111001101110101;
            sine_reg0   <= 36'sb101100100010010010111001101110111101;
        end
        9898: begin
            cosine_reg0 <= 36'sb100110100110111001001100011101000011;
            sine_reg0   <= 36'sb101100100001101011000000101001011011;
        end
        9899: begin
            cosine_reg0 <= 36'sb100110100111010111110010101010111011;
            sine_reg0   <= 36'sb101100100001000011001000010011111100;
        end
        9900: begin
            cosine_reg0 <= 36'sb100110100111110110011001110111011100;
            sine_reg0   <= 36'sb101100100000011011010000101110100010;
        end
        9901: begin
            cosine_reg0 <= 36'sb100110101000010101000010000010100100;
            sine_reg0   <= 36'sb101100011111110011011001111001001111;
        end
        9902: begin
            cosine_reg0 <= 36'sb100110101000110011101011001100010010;
            sine_reg0   <= 36'sb101100011111001011100011110100000011;
        end
        9903: begin
            cosine_reg0 <= 36'sb100110101001010010010101010100100110;
            sine_reg0   <= 36'sb101100011110100011101110011111000000;
        end
        9904: begin
            cosine_reg0 <= 36'sb100110101001110001000000011011011101;
            sine_reg0   <= 36'sb101100011101111011111001111010001001;
        end
        9905: begin
            cosine_reg0 <= 36'sb100110101010001111101100100000110111;
            sine_reg0   <= 36'sb101100011101010100000110000101011101;
        end
        9906: begin
            cosine_reg0 <= 36'sb100110101010101110011001100100110011;
            sine_reg0   <= 36'sb101100011100101100010011000001000000;
        end
        9907: begin
            cosine_reg0 <= 36'sb100110101011001101000111100111001111;
            sine_reg0   <= 36'sb101100011100000100100000101100110010;
        end
        9908: begin
            cosine_reg0 <= 36'sb100110101011101011110110101000001010;
            sine_reg0   <= 36'sb101100011011011100101111001000110101;
        end
        9909: begin
            cosine_reg0 <= 36'sb100110101100001010100110100111100011;
            sine_reg0   <= 36'sb101100011010110100111110010101001011;
        end
        9910: begin
            cosine_reg0 <= 36'sb100110101100101001010111100101011001;
            sine_reg0   <= 36'sb101100011010001101001110010001110101;
        end
        9911: begin
            cosine_reg0 <= 36'sb100110101101001000001001100001101010;
            sine_reg0   <= 36'sb101100011001100101011110111110110100;
        end
        9912: begin
            cosine_reg0 <= 36'sb100110101101100110111100011100010110;
            sine_reg0   <= 36'sb101100011000111101110000011100001011;
        end
        9913: begin
            cosine_reg0 <= 36'sb100110101110000101110000010101011011;
            sine_reg0   <= 36'sb101100011000010110000010101001111010;
        end
        9914: begin
            cosine_reg0 <= 36'sb100110101110100100100101001100111000;
            sine_reg0   <= 36'sb101100010111101110010101101000000100;
        end
        9915: begin
            cosine_reg0 <= 36'sb100110101111000011011011000010101100;
            sine_reg0   <= 36'sb101100010111000110101001010110101001;
        end
        9916: begin
            cosine_reg0 <= 36'sb100110101111100010010001110110110101;
            sine_reg0   <= 36'sb101100010110011110111101110101101011;
        end
        9917: begin
            cosine_reg0 <= 36'sb100110110000000001001001101001010011;
            sine_reg0   <= 36'sb101100010101110111010011000101001101;
        end
        9918: begin
            cosine_reg0 <= 36'sb100110110000100000000010011010000101;
            sine_reg0   <= 36'sb101100010101001111101001000101001110;
        end
        9919: begin
            cosine_reg0 <= 36'sb100110110000111110111100001001001000;
            sine_reg0   <= 36'sb101100010100100111111111110101110010;
        end
        9920: begin
            cosine_reg0 <= 36'sb100110110001011101110110110110011100;
            sine_reg0   <= 36'sb101100010100000000010111010110111001;
        end
        9921: begin
            cosine_reg0 <= 36'sb100110110001111100110010100010000000;
            sine_reg0   <= 36'sb101100010011011000101111101000100100;
        end
        9922: begin
            cosine_reg0 <= 36'sb100110110010011011101111001011110011;
            sine_reg0   <= 36'sb101100010010110001001000101010110110;
        end
        9923: begin
            cosine_reg0 <= 36'sb100110110010111010101100110011110010;
            sine_reg0   <= 36'sb101100010010001001100010011101110001;
        end
        9924: begin
            cosine_reg0 <= 36'sb100110110011011001101011011001111110;
            sine_reg0   <= 36'sb101100010001100001111101000001010100;
        end
        9925: begin
            cosine_reg0 <= 36'sb100110110011111000101010111110010101;
            sine_reg0   <= 36'sb101100010000111010011000010101100011;
        end
        9926: begin
            cosine_reg0 <= 36'sb100110110100010111101011100000110110;
            sine_reg0   <= 36'sb101100010000010010110100011010011110;
        end
        9927: begin
            cosine_reg0 <= 36'sb100110110100110110101101000001011111;
            sine_reg0   <= 36'sb101100001111101011010001010000000111;
        end
        9928: begin
            cosine_reg0 <= 36'sb100110110101010101101111100000001111;
            sine_reg0   <= 36'sb101100001111000011101110110110100000;
        end
        9929: begin
            cosine_reg0 <= 36'sb100110110101110100110010111101000110;
            sine_reg0   <= 36'sb101100001110011100001101001101101010;
        end
        9930: begin
            cosine_reg0 <= 36'sb100110110110010011110111011000000010;
            sine_reg0   <= 36'sb101100001101110100101100010101100111;
        end
        9931: begin
            cosine_reg0 <= 36'sb100110110110110010111100110001000001;
            sine_reg0   <= 36'sb101100001101001101001100001110011000;
        end
        9932: begin
            cosine_reg0 <= 36'sb100110110111010010000011001000000011;
            sine_reg0   <= 36'sb101100001100100101101100110111111110;
        end
        9933: begin
            cosine_reg0 <= 36'sb100110110111110001001010011101000110;
            sine_reg0   <= 36'sb101100001011111110001110010010011100;
        end
        9934: begin
            cosine_reg0 <= 36'sb100110111000010000010010110000001001;
            sine_reg0   <= 36'sb101100001011010110110000011101110010;
        end
        9935: begin
            cosine_reg0 <= 36'sb100110111000101111011100000001001100;
            sine_reg0   <= 36'sb101100001010101111010011011010000011;
        end
        9936: begin
            cosine_reg0 <= 36'sb100110111001001110100110010000001100;
            sine_reg0   <= 36'sb101100001010000111110111000111001111;
        end
        9937: begin
            cosine_reg0 <= 36'sb100110111001101101110001011101001000;
            sine_reg0   <= 36'sb101100001001100000011011100101011001;
        end
        9938: begin
            cosine_reg0 <= 36'sb100110111010001100111101101000000000;
            sine_reg0   <= 36'sb101100001000111001000000110100100010;
        end
        9939: begin
            cosine_reg0 <= 36'sb100110111010101100001010110000110010;
            sine_reg0   <= 36'sb101100001000010001100110110100101010;
        end
        9940: begin
            cosine_reg0 <= 36'sb100110111011001011011000110111011101;
            sine_reg0   <= 36'sb101100000111101010001101100101110101;
        end
        9941: begin
            cosine_reg0 <= 36'sb100110111011101010100111111100000000;
            sine_reg0   <= 36'sb101100000111000010110101001000000011;
        end
        9942: begin
            cosine_reg0 <= 36'sb100110111100001001110111111110011001;
            sine_reg0   <= 36'sb101100000110011011011101011011010110;
        end
        9943: begin
            cosine_reg0 <= 36'sb100110111100101001001000111110101000;
            sine_reg0   <= 36'sb101100000101110100000110011111110000;
        end
        9944: begin
            cosine_reg0 <= 36'sb100110111101001000011010111100101011;
            sine_reg0   <= 36'sb101100000101001100110000010101010001;
        end
        9945: begin
            cosine_reg0 <= 36'sb100110111101100111101101111000100001;
            sine_reg0   <= 36'sb101100000100100101011010111011111100;
        end
        9946: begin
            cosine_reg0 <= 36'sb100110111110000111000001110010001000;
            sine_reg0   <= 36'sb101100000011111110000110010011110010;
        end
        9947: begin
            cosine_reg0 <= 36'sb100110111110100110010110101001100000;
            sine_reg0   <= 36'sb101100000011010110110010011100110100;
        end
        9948: begin
            cosine_reg0 <= 36'sb100110111111000101101100011110100111;
            sine_reg0   <= 36'sb101100000010101111011111010111000100;
        end
        9949: begin
            cosine_reg0 <= 36'sb100110111111100101000011010001011101;
            sine_reg0   <= 36'sb101100000010001000001101000010100100;
        end
        9950: begin
            cosine_reg0 <= 36'sb100111000000000100011011000001111111;
            sine_reg0   <= 36'sb101100000001100000111011011111010101;
        end
        9951: begin
            cosine_reg0 <= 36'sb100111000000100011110011110000001101;
            sine_reg0   <= 36'sb101100000000111001101010101101011000;
        end
        9952: begin
            cosine_reg0 <= 36'sb100111000001000011001101011100000101;
            sine_reg0   <= 36'sb101100000000010010011010101100101111;
        end
        9953: begin
            cosine_reg0 <= 36'sb100111000001100010101000000101100110;
            sine_reg0   <= 36'sb101011111111101011001011011101011100;
        end
        9954: begin
            cosine_reg0 <= 36'sb100111000010000010000011101100110000;
            sine_reg0   <= 36'sb101011111111000011111100111111100000;
        end
        9955: begin
            cosine_reg0 <= 36'sb100111000010100001100000010001100001;
            sine_reg0   <= 36'sb101011111110011100101111010010111101;
        end
        9956: begin
            cosine_reg0 <= 36'sb100111000011000000111101110011110111;
            sine_reg0   <= 36'sb101011111101110101100010010111110011;
        end
        9957: begin
            cosine_reg0 <= 36'sb100111000011100000011100010011110001;
            sine_reg0   <= 36'sb101011111101001110010110001110000110;
        end
        9958: begin
            cosine_reg0 <= 36'sb100111000011111111111011110001001111;
            sine_reg0   <= 36'sb101011111100100111001010110101110101;
        end
        9959: begin
            cosine_reg0 <= 36'sb100111000100011111011100001100001110;
            sine_reg0   <= 36'sb101011111100000000000000001111000011;
        end
        9960: begin
            cosine_reg0 <= 36'sb100111000100111110111101100100101111;
            sine_reg0   <= 36'sb101011111011011000110110011001110001;
        end
        9961: begin
            cosine_reg0 <= 36'sb100111000101011110011111111010101111;
            sine_reg0   <= 36'sb101011111010110001101101010110000001;
        end
        9962: begin
            cosine_reg0 <= 36'sb100111000101111110000011001110001101;
            sine_reg0   <= 36'sb101011111010001010100101000011110100;
        end
        9963: begin
            cosine_reg0 <= 36'sb100111000110011101100111011111001000;
            sine_reg0   <= 36'sb101011111001100011011101100011001100;
        end
        9964: begin
            cosine_reg0 <= 36'sb100111000110111101001100101101011111;
            sine_reg0   <= 36'sb101011111000111100010110110100001010;
        end
        9965: begin
            cosine_reg0 <= 36'sb100111000111011100110010111001010001;
            sine_reg0   <= 36'sb101011111000010101010000110110101111;
        end
        9966: begin
            cosine_reg0 <= 36'sb100111000111111100011010000010011101;
            sine_reg0   <= 36'sb101011110111101110001011101010111110;
        end
        9967: begin
            cosine_reg0 <= 36'sb100111001000011100000010001001000000;
            sine_reg0   <= 36'sb101011110111000111000111010000110111;
        end
        9968: begin
            cosine_reg0 <= 36'sb100111001000111011101011001100111011;
            sine_reg0   <= 36'sb101011110110100000000011101000011101;
        end
        9969: begin
            cosine_reg0 <= 36'sb100111001001011011010101001110001100;
            sine_reg0   <= 36'sb101011110101111001000000110001110000;
        end
        9970: begin
            cosine_reg0 <= 36'sb100111001001111011000000001100110001;
            sine_reg0   <= 36'sb101011110101010001111110101100110011;
        end
        9971: begin
            cosine_reg0 <= 36'sb100111001010011010101100001000101001;
            sine_reg0   <= 36'sb101011110100101010111101011001100110;
        end
        9972: begin
            cosine_reg0 <= 36'sb100111001010111010011001000001110100;
            sine_reg0   <= 36'sb101011110100000011111100111000001100;
        end
        9973: begin
            cosine_reg0 <= 36'sb100111001011011010000110111000001111;
            sine_reg0   <= 36'sb101011110011011100111101001000100101;
        end
        9974: begin
            cosine_reg0 <= 36'sb100111001011111001110101101011111010;
            sine_reg0   <= 36'sb101011110010110101111110001010110011;
        end
        9975: begin
            cosine_reg0 <= 36'sb100111001100011001100101011100110100;
            sine_reg0   <= 36'sb101011110010001110111111111110111001;
        end
        9976: begin
            cosine_reg0 <= 36'sb100111001100111001010110001010111011;
            sine_reg0   <= 36'sb101011110001101000000010100100110110;
        end
        9977: begin
            cosine_reg0 <= 36'sb100111001101011001000111110110001110;
            sine_reg0   <= 36'sb101011110001000001000101111100101101;
        end
        9978: begin
            cosine_reg0 <= 36'sb100111001101111000111010011110101011;
            sine_reg0   <= 36'sb101011110000011010001010000110100000;
        end
        9979: begin
            cosine_reg0 <= 36'sb100111001110011000101110000100010011;
            sine_reg0   <= 36'sb101011101111110011001111000010001111;
        end
        9980: begin
            cosine_reg0 <= 36'sb100111001110111000100010100111000010;
            sine_reg0   <= 36'sb101011101111001100010100101111111100;
        end
        9981: begin
            cosine_reg0 <= 36'sb100111001111011000011000000110111001;
            sine_reg0   <= 36'sb101011101110100101011011001111101001;
        end
        9982: begin
            cosine_reg0 <= 36'sb100111001111111000001110100011110110;
            sine_reg0   <= 36'sb101011101101111110100010100001011000;
        end
        9983: begin
            cosine_reg0 <= 36'sb100111010000011000000101111101110111;
            sine_reg0   <= 36'sb101011101101010111101010100101001001;
        end
        9984: begin
            cosine_reg0 <= 36'sb100111010000110111111110010100111100;
            sine_reg0   <= 36'sb101011101100110000110011011010111110;
        end
        9985: begin
            cosine_reg0 <= 36'sb100111010001010111110111101001000010;
            sine_reg0   <= 36'sb101011101100001001111101000010111001;
        end
        9986: begin
            cosine_reg0 <= 36'sb100111010001110111110001111010001010;
            sine_reg0   <= 36'sb101011101011100011000111011100111100;
        end
        9987: begin
            cosine_reg0 <= 36'sb100111010010010111101101001000010010;
            sine_reg0   <= 36'sb101011101010111100010010101001000111;
        end
        9988: begin
            cosine_reg0 <= 36'sb100111010010110111101001010011011000;
            sine_reg0   <= 36'sb101011101010010101011110100111011100;
        end
        9989: begin
            cosine_reg0 <= 36'sb100111010011010111100110011011011100;
            sine_reg0   <= 36'sb101011101001101110101011010111111101;
        end
        9990: begin
            cosine_reg0 <= 36'sb100111010011110111100100100000011011;
            sine_reg0   <= 36'sb101011101001000111111000111010101100;
        end
        9991: begin
            cosine_reg0 <= 36'sb100111010100010111100011100010010101;
            sine_reg0   <= 36'sb101011101000100001000111001111101001;
        end
        9992: begin
            cosine_reg0 <= 36'sb100111010100110111100011100001001001;
            sine_reg0   <= 36'sb101011100111111010010110010110110110;
        end
        9993: begin
            cosine_reg0 <= 36'sb100111010101010111100100011100110101;
            sine_reg0   <= 36'sb101011100111010011100110010000010101;
        end
        9994: begin
            cosine_reg0 <= 36'sb100111010101110111100110010101011001;
            sine_reg0   <= 36'sb101011100110101100110110111100000111;
        end
        9995: begin
            cosine_reg0 <= 36'sb100111010110010111101001001010110010;
            sine_reg0   <= 36'sb101011100110000110001000011010001110;
        end
        9996: begin
            cosine_reg0 <= 36'sb100111010110110111101100111101000000;
            sine_reg0   <= 36'sb101011100101011111011010101010101011;
        end
        9997: begin
            cosine_reg0 <= 36'sb100111010111010111110001101100000001;
            sine_reg0   <= 36'sb101011100100111000101101101101011111;
        end
        9998: begin
            cosine_reg0 <= 36'sb100111010111110111110111010111110101;
            sine_reg0   <= 36'sb101011100100010010000001100010101101;
        end
        9999: begin
            cosine_reg0 <= 36'sb100111011000010111111110000000011001;
            sine_reg0   <= 36'sb101011100011101011010110001010010110;
        end
        10000: begin
            cosine_reg0 <= 36'sb100111011000111000000101100101101101;
            sine_reg0   <= 36'sb101011100011000100101011100100011011;
        end
        10001: begin
            cosine_reg0 <= 36'sb100111011001011000001110000111110000;
            sine_reg0   <= 36'sb101011100010011110000001110000111101;
        end
        10002: begin
            cosine_reg0 <= 36'sb100111011001111000010111100110100000;
            sine_reg0   <= 36'sb101011100001110111011000101111111110;
        end
        10003: begin
            cosine_reg0 <= 36'sb100111011010011000100010000001111011;
            sine_reg0   <= 36'sb101011100001010000110000100001100000;
        end
        10004: begin
            cosine_reg0 <= 36'sb100111011010111000101101011010000010;
            sine_reg0   <= 36'sb101011100000101010001001000101100101;
        end
        10005: begin
            cosine_reg0 <= 36'sb100111011011011000111001101110110010;
            sine_reg0   <= 36'sb101011100000000011100010011100001101;
        end
        10006: begin
            cosine_reg0 <= 36'sb100111011011111001000111000000001010;
            sine_reg0   <= 36'sb101011011111011100111100100101011001;
        end
        10007: begin
            cosine_reg0 <= 36'sb100111011100011001010101001110001010;
            sine_reg0   <= 36'sb101011011110110110010111100001001101;
        end
        10008: begin
            cosine_reg0 <= 36'sb100111011100111001100100011000101111;
            sine_reg0   <= 36'sb101011011110001111110011001111101000;
        end
        10009: begin
            cosine_reg0 <= 36'sb100111011101011001110100011111111000;
            sine_reg0   <= 36'sb101011011101101001001111110000101110;
        end
        10010: begin
            cosine_reg0 <= 36'sb100111011101111010000101100011100101;
            sine_reg0   <= 36'sb101011011101000010101101000100011110;
        end
        10011: begin
            cosine_reg0 <= 36'sb100111011110011010010111100011110100;
            sine_reg0   <= 36'sb101011011100011100001011001010111010;
        end
        10012: begin
            cosine_reg0 <= 36'sb100111011110111010101010100000100100;
            sine_reg0   <= 36'sb101011011011110101101010000100000101;
        end
        10013: begin
            cosine_reg0 <= 36'sb100111011111011010111110011001110011;
            sine_reg0   <= 36'sb101011011011001111001001101111111111;
        end
        10014: begin
            cosine_reg0 <= 36'sb100111011111111011010011001111100001;
            sine_reg0   <= 36'sb101011011010101000101010001110101011;
        end
        10015: begin
            cosine_reg0 <= 36'sb100111100000011011101001000001101100;
            sine_reg0   <= 36'sb101011011010000010001011100000001000;
        end
        10016: begin
            cosine_reg0 <= 36'sb100111100000111011111111110000010010;
            sine_reg0   <= 36'sb101011011001011011101101100100011010;
        end
        10017: begin
            cosine_reg0 <= 36'sb100111100001011100010111011011010011;
            sine_reg0   <= 36'sb101011011000110101010000011011100001;
        end
        10018: begin
            cosine_reg0 <= 36'sb100111100001111100110000000010101110;
            sine_reg0   <= 36'sb101011011000001110110100000101011111;
        end
        10019: begin
            cosine_reg0 <= 36'sb100111100010011101001001100110100000;
            sine_reg0   <= 36'sb101011010111101000011000100010010101;
        end
        10020: begin
            cosine_reg0 <= 36'sb100111100010111101100100000110101010;
            sine_reg0   <= 36'sb101011010111000001111101110010000101;
        end
        10021: begin
            cosine_reg0 <= 36'sb100111100011011101111111100011001000;
            sine_reg0   <= 36'sb101011010110011011100011110100110001;
        end
        10022: begin
            cosine_reg0 <= 36'sb100111100011111110011011111011111100;
            sine_reg0   <= 36'sb101011010101110101001010101010011010;
        end
        10023: begin
            cosine_reg0 <= 36'sb100111100100011110111001010001000010;
            sine_reg0   <= 36'sb101011010101001110110010010011000000;
        end
        10024: begin
            cosine_reg0 <= 36'sb100111100100111111010111100010011010;
            sine_reg0   <= 36'sb101011010100101000011010101110100111;
        end
        10025: begin
            cosine_reg0 <= 36'sb100111100101011111110110110000000011;
            sine_reg0   <= 36'sb101011010100000010000011111101001111;
        end
        10026: begin
            cosine_reg0 <= 36'sb100111100110000000010110111001111011;
            sine_reg0   <= 36'sb101011010011011011101101111110111001;
        end
        10027: begin
            cosine_reg0 <= 36'sb100111100110100000111000000000000001;
            sine_reg0   <= 36'sb101011010010110101011000110011101000;
        end
        10028: begin
            cosine_reg0 <= 36'sb100111100111000001011010000010010100;
            sine_reg0   <= 36'sb101011010010001111000100011011011101;
        end
        10029: begin
            cosine_reg0 <= 36'sb100111100111100001111101000000110010;
            sine_reg0   <= 36'sb101011010001101000110000110110011000;
        end
        10030: begin
            cosine_reg0 <= 36'sb100111101000000010100000111011011011;
            sine_reg0   <= 36'sb101011010001000010011110000100011101;
        end
        10031: begin
            cosine_reg0 <= 36'sb100111101000100011000101110010001101;
            sine_reg0   <= 36'sb101011010000011100001100000101101011;
        end
        10032: begin
            cosine_reg0 <= 36'sb100111101001000011101011100101000110;
            sine_reg0   <= 36'sb101011001111110101111010111010000110;
        end
        10033: begin
            cosine_reg0 <= 36'sb100111101001100100010010010100000111;
            sine_reg0   <= 36'sb101011001111001111101010100001101101;
        end
        10034: begin
            cosine_reg0 <= 36'sb100111101010000100111001111111001100;
            sine_reg0   <= 36'sb101011001110101001011010111100100011;
        end
        10035: begin
            cosine_reg0 <= 36'sb100111101010100101100010100110010101;
            sine_reg0   <= 36'sb101011001110000011001100001010101001;
        end
        10036: begin
            cosine_reg0 <= 36'sb100111101011000110001100001001100010;
            sine_reg0   <= 36'sb101011001101011100111110001100000000;
        end
        10037: begin
            cosine_reg0 <= 36'sb100111101011100110110110101000101111;
            sine_reg0   <= 36'sb101011001100110110110001000000101011;
        end
        10038: begin
            cosine_reg0 <= 36'sb100111101100000111100010000011111101;
            sine_reg0   <= 36'sb101011001100010000100100101000101001;
        end
        10039: begin
            cosine_reg0 <= 36'sb100111101100101000001110011011001010;
            sine_reg0   <= 36'sb101011001011101010011001000011111110;
        end
        10040: begin
            cosine_reg0 <= 36'sb100111101101001000111011101110010101;
            sine_reg0   <= 36'sb101011001011000100001110010010101010;
        end
        10041: begin
            cosine_reg0 <= 36'sb100111101101101001101001111101011100;
            sine_reg0   <= 36'sb101011001010011110000100010100110000;
        end
        10042: begin
            cosine_reg0 <= 36'sb100111101110001010011001001000011110;
            sine_reg0   <= 36'sb101011001001110111111011001010001111;
        end
        10043: begin
            cosine_reg0 <= 36'sb100111101110101011001001001111011011;
            sine_reg0   <= 36'sb101011001001010001110010110011001010;
        end
        10044: begin
            cosine_reg0 <= 36'sb100111101111001011111010010010010000;
            sine_reg0   <= 36'sb101011001000101011101011001111100011;
        end
        10045: begin
            cosine_reg0 <= 36'sb100111101111101100101100010000111100;
            sine_reg0   <= 36'sb101011001000000101100100011111011010;
        end
        10046: begin
            cosine_reg0 <= 36'sb100111110000001101011111001011011110;
            sine_reg0   <= 36'sb101011000111011111011110100010110010;
        end
        10047: begin
            cosine_reg0 <= 36'sb100111110000101110010011000001110110;
            sine_reg0   <= 36'sb101011000110111001011001011001101011;
        end
        10048: begin
            cosine_reg0 <= 36'sb100111110001001111000111110100000001;
            sine_reg0   <= 36'sb101011000110010011010101000100001000;
        end
        10049: begin
            cosine_reg0 <= 36'sb100111110001101111111101100001111110;
            sine_reg0   <= 36'sb101011000101101101010001100010001001;
        end
        10050: begin
            cosine_reg0 <= 36'sb100111110010010000110100001011101101;
            sine_reg0   <= 36'sb101011000101000111001110110011110000;
        end
        10051: begin
            cosine_reg0 <= 36'sb100111110010110001101011110001001011;
            sine_reg0   <= 36'sb101011000100100001001100111000111111;
        end
        10052: begin
            cosine_reg0 <= 36'sb100111110011010010100100010010011000;
            sine_reg0   <= 36'sb101011000011111011001011110001110111;
        end
        10053: begin
            cosine_reg0 <= 36'sb100111110011110011011101101111010010;
            sine_reg0   <= 36'sb101011000011010101001011011110011001;
        end
        10054: begin
            cosine_reg0 <= 36'sb100111110100010100011000000111111000;
            sine_reg0   <= 36'sb101011000010101111001011111110100111;
        end
        10055: begin
            cosine_reg0 <= 36'sb100111110100110101010011011100001001;
            sine_reg0   <= 36'sb101011000010001001001101010010100011;
        end
        10056: begin
            cosine_reg0 <= 36'sb100111110101010110001111101100000011;
            sine_reg0   <= 36'sb101011000001100011001111011010001101;
        end
        10057: begin
            cosine_reg0 <= 36'sb100111110101110111001100110111100110;
            sine_reg0   <= 36'sb101011000000111101010010010101101000;
        end
        10058: begin
            cosine_reg0 <= 36'sb100111110110011000001010111110110000;
            sine_reg0   <= 36'sb101011000000010111010110000100110101;
        end
        10059: begin
            cosine_reg0 <= 36'sb100111110110111001001010000001011111;
            sine_reg0   <= 36'sb101010111111110001011010100111110101;
        end
        10060: begin
            cosine_reg0 <= 36'sb100111110111011010001001111111110010;
            sine_reg0   <= 36'sb101010111111001011011111111110101010;
        end
        10061: begin
            cosine_reg0 <= 36'sb100111110111111011001010111001101001;
            sine_reg0   <= 36'sb101010111110100101100110001001010101;
        end
        10062: begin
            cosine_reg0 <= 36'sb100111111000011100001100101111000010;
            sine_reg0   <= 36'sb101010111101111111101101000111111000;
        end
        10063: begin
            cosine_reg0 <= 36'sb100111111000111101001111011111111011;
            sine_reg0   <= 36'sb101010111101011001110100111010010100;
        end
        10064: begin
            cosine_reg0 <= 36'sb100111111001011110010011001100010011;
            sine_reg0   <= 36'sb101010111100110011111101100000101010;
        end
        10065: begin
            cosine_reg0 <= 36'sb100111111001111111010111110100001010;
            sine_reg0   <= 36'sb101010111100001110000110111010111101;
        end
        10066: begin
            cosine_reg0 <= 36'sb100111111010100000011101010111011101;
            sine_reg0   <= 36'sb101010111011101000010001001001001101;
        end
        10067: begin
            cosine_reg0 <= 36'sb100111111011000001100011110110001100;
            sine_reg0   <= 36'sb101010111011000010011100001011011100;
        end
        10068: begin
            cosine_reg0 <= 36'sb100111111011100010101011010000010101;
            sine_reg0   <= 36'sb101010111010011100101000000001101011;
        end
        10069: begin
            cosine_reg0 <= 36'sb100111111100000011110011100101110111;
            sine_reg0   <= 36'sb101010111001110110110100101011111100;
        end
        10070: begin
            cosine_reg0 <= 36'sb100111111100100100111100110110110000;
            sine_reg0   <= 36'sb101010111001010001000010001010010001;
        end
        10071: begin
            cosine_reg0 <= 36'sb100111111101000110000111000011000000;
            sine_reg0   <= 36'sb101010111000101011010000011100101011;
        end
        10072: begin
            cosine_reg0 <= 36'sb100111111101100111010010001010100101;
            sine_reg0   <= 36'sb101010111000000101011111100011001010;
        end
        10073: begin
            cosine_reg0 <= 36'sb100111111110001000011110001101011110;
            sine_reg0   <= 36'sb101010110111011111101111011101110010;
        end
        10074: begin
            cosine_reg0 <= 36'sb100111111110101001101011001011101001;
            sine_reg0   <= 36'sb101010110110111010000000001100100010;
        end
        10075: begin
            cosine_reg0 <= 36'sb100111111111001010111001000101000110;
            sine_reg0   <= 36'sb101010110110010100010001101111011101;
        end
        10076: begin
            cosine_reg0 <= 36'sb100111111111101100000111111001110011;
            sine_reg0   <= 36'sb101010110101101110100100000110100101;
        end
        10077: begin
            cosine_reg0 <= 36'sb101000000000001101010111101001101110;
            sine_reg0   <= 36'sb101010110101001000110111010001111010;
        end
        10078: begin
            cosine_reg0 <= 36'sb101000000000101110101000010100110110;
            sine_reg0   <= 36'sb101010110100100011001011010001011101;
        end
        10079: begin
            cosine_reg0 <= 36'sb101000000001001111111001111011001011;
            sine_reg0   <= 36'sb101010110011111101100000000101010010;
        end
        10080: begin
            cosine_reg0 <= 36'sb101000000001110001001100011100101011;
            sine_reg0   <= 36'sb101010110011010111110101101101011000;
        end
        10081: begin
            cosine_reg0 <= 36'sb101000000010010010011111111001010100;
            sine_reg0   <= 36'sb101010110010110010001100001001110001;
        end
        10082: begin
            cosine_reg0 <= 36'sb101000000010110011110100010001000110;
            sine_reg0   <= 36'sb101010110010001100100011011010100000;
        end
        10083: begin
            cosine_reg0 <= 36'sb101000000011010101001001100011111110;
            sine_reg0   <= 36'sb101010110001100110111011011111100100;
        end
        10084: begin
            cosine_reg0 <= 36'sb101000000011110110011111110001111100;
            sine_reg0   <= 36'sb101010110001000001010100011001000000;
        end
        10085: begin
            cosine_reg0 <= 36'sb101000000100010111110110111010111111;
            sine_reg0   <= 36'sb101010110000011011101110000110110110;
        end
        10086: begin
            cosine_reg0 <= 36'sb101000000100111001001110111111000101;
            sine_reg0   <= 36'sb101010101111110110001000101001000110;
        end
        10087: begin
            cosine_reg0 <= 36'sb101000000101011010100111111110001100;
            sine_reg0   <= 36'sb101010101111010000100011111111110010;
        end
        10088: begin
            cosine_reg0 <= 36'sb101000000101111100000001111000010101;
            sine_reg0   <= 36'sb101010101110101011000000001010111011;
        end
        10089: begin
            cosine_reg0 <= 36'sb101000000110011101011100101101011100;
            sine_reg0   <= 36'sb101010101110000101011101001010100100;
        end
        10090: begin
            cosine_reg0 <= 36'sb101000000110111110111000011101100010;
            sine_reg0   <= 36'sb101010101101011111111010111110101101;
        end
        10091: begin
            cosine_reg0 <= 36'sb101000000111100000010101001000100100;
            sine_reg0   <= 36'sb101010101100111010011001100111010111;
        end
        10092: begin
            cosine_reg0 <= 36'sb101000001000000001110010101110100001;
            sine_reg0   <= 36'sb101010101100010100111001000100100101;
        end
        10093: begin
            cosine_reg0 <= 36'sb101000001000100011010001001111011001;
            sine_reg0   <= 36'sb101010101011101111011001010110011000;
        end
        10094: begin
            cosine_reg0 <= 36'sb101000001001000100110000101011001010;
            sine_reg0   <= 36'sb101010101011001001111010011100110001;
        end
        10095: begin
            cosine_reg0 <= 36'sb101000001001100110010001000001110010;
            sine_reg0   <= 36'sb101010101010100100011100010111110001;
        end
        10096: begin
            cosine_reg0 <= 36'sb101000001010000111110010010011010000;
            sine_reg0   <= 36'sb101010101001111110111111000111011011;
        end
        10097: begin
            cosine_reg0 <= 36'sb101000001010101001010100011111100011;
            sine_reg0   <= 36'sb101010101001011001100010101011101111;
        end
        10098: begin
            cosine_reg0 <= 36'sb101000001011001010110111100110101010;
            sine_reg0   <= 36'sb101010101000110100000111000100101111;
        end
        10099: begin
            cosine_reg0 <= 36'sb101000001011101100011011101000100011;
            sine_reg0   <= 36'sb101010101000001110101100010010011100;
        end
        10100: begin
            cosine_reg0 <= 36'sb101000001100001110000000100101001110;
            sine_reg0   <= 36'sb101010100111101001010010010100111001;
        end
        10101: begin
            cosine_reg0 <= 36'sb101000001100101111100110011100101000;
            sine_reg0   <= 36'sb101010100111000011111001001100000101;
        end
        10102: begin
            cosine_reg0 <= 36'sb101000001101010001001101001110110001;
            sine_reg0   <= 36'sb101010100110011110100000111000000011;
        end
        10103: begin
            cosine_reg0 <= 36'sb101000001101110010110100111011100110;
            sine_reg0   <= 36'sb101010100101111001001001011000110101;
        end
        10104: begin
            cosine_reg0 <= 36'sb101000001110010100011101100011001000;
            sine_reg0   <= 36'sb101010100101010011110010101110011011;
        end
        10105: begin
            cosine_reg0 <= 36'sb101000001110110110000111000101010100;
            sine_reg0   <= 36'sb101010100100101110011100111000110111;
        end
        10106: begin
            cosine_reg0 <= 36'sb101000001111010111110001100010001010;
            sine_reg0   <= 36'sb101010100100001001000111111000001010;
        end
        10107: begin
            cosine_reg0 <= 36'sb101000001111111001011100111001101000;
            sine_reg0   <= 36'sb101010100011100011110011101100010111;
        end
        10108: begin
            cosine_reg0 <= 36'sb101000010000011011001001001011101100;
            sine_reg0   <= 36'sb101010100010111110100000010101011110;
        end
        10109: begin
            cosine_reg0 <= 36'sb101000010000111100110110011000010110;
            sine_reg0   <= 36'sb101010100010011001001101110011100000;
        end
        10110: begin
            cosine_reg0 <= 36'sb101000010001011110100100011111100011;
            sine_reg0   <= 36'sb101010100001110011111100000110100000;
        end
        10111: begin
            cosine_reg0 <= 36'sb101000010010000000010011100001010100;
            sine_reg0   <= 36'sb101010100001001110101011001110011111;
        end
        10112: begin
            cosine_reg0 <= 36'sb101000010010100010000011011101100110;
            sine_reg0   <= 36'sb101010100000101001011011001011011101;
        end
        10113: begin
            cosine_reg0 <= 36'sb101000010011000011110100010100011000;
            sine_reg0   <= 36'sb101010100000000100001011111101011110;
        end
        10114: begin
            cosine_reg0 <= 36'sb101000010011100101100110000101101010;
            sine_reg0   <= 36'sb101010011111011110111101100100100001;
        end
        10115: begin
            cosine_reg0 <= 36'sb101000010100000111011000110001011000;
            sine_reg0   <= 36'sb101010011110111001110000000000101000;
        end
        10116: begin
            cosine_reg0 <= 36'sb101000010100101001001100010111100100;
            sine_reg0   <= 36'sb101010011110010100100011010001110110;
        end
        10117: begin
            cosine_reg0 <= 36'sb101000010101001011000000111000001010;
            sine_reg0   <= 36'sb101010011101101111010111011000001011;
        end
        10118: begin
            cosine_reg0 <= 36'sb101000010101101100110110010011001001;
            sine_reg0   <= 36'sb101010011101001010001100010011101000;
        end
        10119: begin
            cosine_reg0 <= 36'sb101000010110001110101100101000100010;
            sine_reg0   <= 36'sb101010011100100101000010000100010000;
        end
        10120: begin
            cosine_reg0 <= 36'sb101000010110110000100011111000010001;
            sine_reg0   <= 36'sb101010011011111111111000101010000011;
        end
        10121: begin
            cosine_reg0 <= 36'sb101000010111010010011100000010010110;
            sine_reg0   <= 36'sb101010011011011010110000000101000011;
        end
        10122: begin
            cosine_reg0 <= 36'sb101000010111110100010101000110101111;
            sine_reg0   <= 36'sb101010011010110101101000010101010010;
        end
        10123: begin
            cosine_reg0 <= 36'sb101000011000010110001111000101011100;
            sine_reg0   <= 36'sb101010011010010000100001011010110000;
        end
        10124: begin
            cosine_reg0 <= 36'sb101000011000111000001001111110011011;
            sine_reg0   <= 36'sb101010011001101011011011010101100000;
        end
        10125: begin
            cosine_reg0 <= 36'sb101000011001011010000101110001101010;
            sine_reg0   <= 36'sb101010011001000110010110000101100011;
        end
        10126: begin
            cosine_reg0 <= 36'sb101000011001111100000010011111001000;
            sine_reg0   <= 36'sb101010011000100001010001101010111010;
        end
        10127: begin
            cosine_reg0 <= 36'sb101000011010011110000000000110110100;
            sine_reg0   <= 36'sb101010010111111100001110000101100110;
        end
        10128: begin
            cosine_reg0 <= 36'sb101000011010111111111110101000101101;
            sine_reg0   <= 36'sb101010010111010111001011010101101001;
        end
        10129: begin
            cosine_reg0 <= 36'sb101000011011100001111110000100110001;
            sine_reg0   <= 36'sb101010010110110010001001011011000101;
        end
        10130: begin
            cosine_reg0 <= 36'sb101000011100000011111110011010111111;
            sine_reg0   <= 36'sb101010010110001101001000010101111011;
        end
        10131: begin
            cosine_reg0 <= 36'sb101000011100100101111111101011010110;
            sine_reg0   <= 36'sb101010010101101000001000000110001100;
        end
        10132: begin
            cosine_reg0 <= 36'sb101000011101001000000001110101110100;
            sine_reg0   <= 36'sb101010010101000011001000101011111010;
        end
        10133: begin
            cosine_reg0 <= 36'sb101000011101101010000100111010011000;
            sine_reg0   <= 36'sb101010010100011110001010000111000110;
        end
        10134: begin
            cosine_reg0 <= 36'sb101000011110001100001000111001000010;
            sine_reg0   <= 36'sb101010010011111001001100010111110001;
        end
        10135: begin
            cosine_reg0 <= 36'sb101000011110101110001101110001101110;
            sine_reg0   <= 36'sb101010010011010100001111011101111110;
        end
        10136: begin
            cosine_reg0 <= 36'sb101000011111010000010011100100011101;
            sine_reg0   <= 36'sb101010010010101111010011011001101101;
        end
        10137: begin
            cosine_reg0 <= 36'sb101000011111110010011010010001001100;
            sine_reg0   <= 36'sb101010010010001010011000001011000000;
        end
        10138: begin
            cosine_reg0 <= 36'sb101000100000010100100001110111111011;
            sine_reg0   <= 36'sb101010010001100101011101110001111000;
        end
        10139: begin
            cosine_reg0 <= 36'sb101000100000110110101010011000101000;
            sine_reg0   <= 36'sb101010010001000000100100001110010111;
        end
        10140: begin
            cosine_reg0 <= 36'sb101000100001011000110011110011010010;
            sine_reg0   <= 36'sb101010010000011011101011100000011110;
        end
        10141: begin
            cosine_reg0 <= 36'sb101000100001111010111110000111110111;
            sine_reg0   <= 36'sb101010001111110110110011101000001110;
        end
        10142: begin
            cosine_reg0 <= 36'sb101000100010011101001001010110010111;
            sine_reg0   <= 36'sb101010001111010001111100100101101010;
        end
        10143: begin
            cosine_reg0 <= 36'sb101000100010111111010101011110110000;
            sine_reg0   <= 36'sb101010001110101101000110011000110010;
        end
        10144: begin
            cosine_reg0 <= 36'sb101000100011100001100010100001000000;
            sine_reg0   <= 36'sb101010001110001000010001000001100111;
        end
        10145: begin
            cosine_reg0 <= 36'sb101000100100000011110000011101000110;
            sine_reg0   <= 36'sb101010001101100011011100100000001100;
        end
        10146: begin
            cosine_reg0 <= 36'sb101000100100100101111111010011000010;
            sine_reg0   <= 36'sb101010001100111110101000110100100010;
        end
        10147: begin
            cosine_reg0 <= 36'sb101000100101001000001111000010110001;
            sine_reg0   <= 36'sb101010001100011001110101111110101010;
        end
        10148: begin
            cosine_reg0 <= 36'sb101000100101101010011111101100010010;
            sine_reg0   <= 36'sb101010001011110101000011111110100101;
        end
        10149: begin
            cosine_reg0 <= 36'sb101000100110001100110001001111100101;
            sine_reg0   <= 36'sb101010001011010000010010110100010101;
        end
        10150: begin
            cosine_reg0 <= 36'sb101000100110101111000011101100100111;
            sine_reg0   <= 36'sb101010001010101011100010011111111100;
        end
        10151: begin
            cosine_reg0 <= 36'sb101000100111010001010111000011010111;
            sine_reg0   <= 36'sb101010001010000110110011000001011010;
        end
        10152: begin
            cosine_reg0 <= 36'sb101000100111110011101011010011110101;
            sine_reg0   <= 36'sb101010001001100010000100011000110001;
        end
        10153: begin
            cosine_reg0 <= 36'sb101000101000010110000000011101111110;
            sine_reg0   <= 36'sb101010001000111101010110100110000011;
        end
        10154: begin
            cosine_reg0 <= 36'sb101000101000111000010110100001110001;
            sine_reg0   <= 36'sb101010001000011000101001101001010001;
        end
        10155: begin
            cosine_reg0 <= 36'sb101000101001011010101101011111001110;
            sine_reg0   <= 36'sb101010000111110011111101100010011100;
        end
        10156: begin
            cosine_reg0 <= 36'sb101000101001111101000101010110010010;
            sine_reg0   <= 36'sb101010000111001111010010010001100111;
        end
        10157: begin
            cosine_reg0 <= 36'sb101000101010011111011110000110111101;
            sine_reg0   <= 36'sb101010000110101010100111110110110001;
        end
        10158: begin
            cosine_reg0 <= 36'sb101000101011000001110111110001001101;
            sine_reg0   <= 36'sb101010000110000101111110010001111101;
        end
        10159: begin
            cosine_reg0 <= 36'sb101000101011100100010010010101000000;
            sine_reg0   <= 36'sb101010000101100001010101100011001100;
        end
        10160: begin
            cosine_reg0 <= 36'sb101000101100000110101101110010010111;
            sine_reg0   <= 36'sb101010000100111100101101101010100000;
        end
        10161: begin
            cosine_reg0 <= 36'sb101000101100101001001010001001001110;
            sine_reg0   <= 36'sb101010000100011000000110100111111001;
        end
        10162: begin
            cosine_reg0 <= 36'sb101000101101001011100111011001100101;
            sine_reg0   <= 36'sb101010000011110011100000011011011010;
        end
        10163: begin
            cosine_reg0 <= 36'sb101000101101101110000101100011011010;
            sine_reg0   <= 36'sb101010000011001110111011000101000100;
        end
        10164: begin
            cosine_reg0 <= 36'sb101000101110010000100100100110101100;
            sine_reg0   <= 36'sb101010000010101010010110100100110111;
        end
        10165: begin
            cosine_reg0 <= 36'sb101000101110110011000100100011011011;
            sine_reg0   <= 36'sb101010000010000101110010111010110111;
        end
        10166: begin
            cosine_reg0 <= 36'sb101000101111010101100101011001100011;
            sine_reg0   <= 36'sb101010000001100001010000000111000011;
        end
        10167: begin
            cosine_reg0 <= 36'sb101000101111111000000111001001000101;
            sine_reg0   <= 36'sb101010000000111100101110001001011101;
        end
        10168: begin
            cosine_reg0 <= 36'sb101000110000011010101001110001111111;
            sine_reg0   <= 36'sb101010000000011000001101000010000111;
        end
        10169: begin
            cosine_reg0 <= 36'sb101000110000111101001101010100001111;
            sine_reg0   <= 36'sb101001111111110011101100110001000011;
        end
        10170: begin
            cosine_reg0 <= 36'sb101000110001011111110001101111110100;
            sine_reg0   <= 36'sb101001111111001111001101010110010001;
        end
        10171: begin
            cosine_reg0 <= 36'sb101000110010000010010111000100101101;
            sine_reg0   <= 36'sb101001111110101010101110110001110011;
        end
        10172: begin
            cosine_reg0 <= 36'sb101000110010100100111101010010111001;
            sine_reg0   <= 36'sb101001111110000110010001000011101010;
        end
        10173: begin
            cosine_reg0 <= 36'sb101000110011000111100100011010010101;
            sine_reg0   <= 36'sb101001111101100001110100001011111000;
        end
        10174: begin
            cosine_reg0 <= 36'sb101000110011101010001100011011000010;
            sine_reg0   <= 36'sb101001111100111101011000001010011110;
        end
        10175: begin
            cosine_reg0 <= 36'sb101000110100001100110101010100111101;
            sine_reg0   <= 36'sb101001111100011000111100111111011110;
        end
        10176: begin
            cosine_reg0 <= 36'sb101000110100101111011111001000000101;
            sine_reg0   <= 36'sb101001111011110100100010101010111001;
        end
        10177: begin
            cosine_reg0 <= 36'sb101000110101010010001001110100011001;
            sine_reg0   <= 36'sb101001111011010000001001001100110001;
        end
        10178: begin
            cosine_reg0 <= 36'sb101000110101110100110101011001110111;
            sine_reg0   <= 36'sb101001111010101011110000100101000110;
        end
        10179: begin
            cosine_reg0 <= 36'sb101000110110010111100001111000011110;
            sine_reg0   <= 36'sb101001111010000111011000110011111010;
        end
        10180: begin
            cosine_reg0 <= 36'sb101000110110111010001111010000001101;
            sine_reg0   <= 36'sb101001111001100011000001111001001111;
        end
        10181: begin
            cosine_reg0 <= 36'sb101000110111011100111101100001000011;
            sine_reg0   <= 36'sb101001111000111110101011110101000110;
        end
        10182: begin
            cosine_reg0 <= 36'sb101000110111111111101100101010111110;
            sine_reg0   <= 36'sb101001111000011010010110100111100001;
        end
        10183: begin
            cosine_reg0 <= 36'sb101000111000100010011100101101111100;
            sine_reg0   <= 36'sb101001110111110110000010010000100000;
        end
        10184: begin
            cosine_reg0 <= 36'sb101000111001000101001101101001111101;
            sine_reg0   <= 36'sb101001110111010001101110110000000110;
        end
        10185: begin
            cosine_reg0 <= 36'sb101000111001100111111111011110111111;
            sine_reg0   <= 36'sb101001110110101101011100000110010011;
        end
        10186: begin
            cosine_reg0 <= 36'sb101000111010001010110010001101000001;
            sine_reg0   <= 36'sb101001110110001001001010010011001001;
        end
        10187: begin
            cosine_reg0 <= 36'sb101000111010101101100101110100000001;
            sine_reg0   <= 36'sb101001110101100100111001010110101010;
        end
        10188: begin
            cosine_reg0 <= 36'sb101000111011010000011010010011111110;
            sine_reg0   <= 36'sb101001110101000000101001010000110110;
        end
        10189: begin
            cosine_reg0 <= 36'sb101000111011110011001111101100110111;
            sine_reg0   <= 36'sb101001110100011100011010000001110000;
        end
        10190: begin
            cosine_reg0 <= 36'sb101000111100010110000101111110101011;
            sine_reg0   <= 36'sb101001110011111000001011101001011000;
        end
        10191: begin
            cosine_reg0 <= 36'sb101000111100111000111101001001010111;
            sine_reg0   <= 36'sb101001110011010011111110000111110000;
        end
        10192: begin
            cosine_reg0 <= 36'sb101000111101011011110101001100111011;
            sine_reg0   <= 36'sb101001110010101111110001011100111010;
        end
        10193: begin
            cosine_reg0 <= 36'sb101000111101111110101110001001010101;
            sine_reg0   <= 36'sb101001110010001011100101101000110110;
        end
        10194: begin
            cosine_reg0 <= 36'sb101000111110100001100111111110100101;
            sine_reg0   <= 36'sb101001110001100111011010101011100111;
        end
        10195: begin
            cosine_reg0 <= 36'sb101000111111000100100010101100101000;
            sine_reg0   <= 36'sb101001110001000011010000100101001101;
        end
        10196: begin
            cosine_reg0 <= 36'sb101000111111100111011110010011011101;
            sine_reg0   <= 36'sb101001110000011111000111010101101010;
        end
        10197: begin
            cosine_reg0 <= 36'sb101001000000001010011010110011000011;
            sine_reg0   <= 36'sb101001101111111010111110111101000000;
        end
        10198: begin
            cosine_reg0 <= 36'sb101001000000101101011000001011011001;
            sine_reg0   <= 36'sb101001101111010110110111011011001111;
        end
        10199: begin
            cosine_reg0 <= 36'sb101001000001010000010110011100011101;
            sine_reg0   <= 36'sb101001101110110010110000110000011010;
        end
        10200: begin
            cosine_reg0 <= 36'sb101001000001110011010101100110001110;
            sine_reg0   <= 36'sb101001101110001110101010111100100001;
        end
        10201: begin
            cosine_reg0 <= 36'sb101001000010010110010101101000101011;
            sine_reg0   <= 36'sb101001101101101010100101111111100110;
        end
        10202: begin
            cosine_reg0 <= 36'sb101001000010111001010110100011110010;
            sine_reg0   <= 36'sb101001101101000110100001111001101010;
        end
        10203: begin
            cosine_reg0 <= 36'sb101001000011011100011000010111100010;
            sine_reg0   <= 36'sb101001101100100010011110101010101111;
        end
        10204: begin
            cosine_reg0 <= 36'sb101001000011111111011011000011111001;
            sine_reg0   <= 36'sb101001101011111110011100010010110111;
        end
        10205: begin
            cosine_reg0 <= 36'sb101001000100100010011110101000110110;
            sine_reg0   <= 36'sb101001101011011010011010110010000001;
        end
        10206: begin
            cosine_reg0 <= 36'sb101001000101000101100011000110011001;
            sine_reg0   <= 36'sb101001101010110110011010001000010001;
        end
        10207: begin
            cosine_reg0 <= 36'sb101001000101101000101000011100011110;
            sine_reg0   <= 36'sb101001101010010010011010010101100111;
        end
        10208: begin
            cosine_reg0 <= 36'sb101001000110001011101110101011000110;
            sine_reg0   <= 36'sb101001101001101110011011011010000101;
        end
        10209: begin
            cosine_reg0 <= 36'sb101001000110101110110101110010001111;
            sine_reg0   <= 36'sb101001101001001010011101010101101011;
        end
        10210: begin
            cosine_reg0 <= 36'sb101001000111010001111101110001110111;
            sine_reg0   <= 36'sb101001101000100110100000001000011100;
        end
        10211: begin
            cosine_reg0 <= 36'sb101001000111110101000110101001111101;
            sine_reg0   <= 36'sb101001101000000010100011110010011001;
        end
        10212: begin
            cosine_reg0 <= 36'sb101001001000011000010000011010011111;
            sine_reg0   <= 36'sb101001100111011110101000010011100011;
        end
        10213: begin
            cosine_reg0 <= 36'sb101001001000111011011011000011011101;
            sine_reg0   <= 36'sb101001100110111010101101101011111100;
        end
        10214: begin
            cosine_reg0 <= 36'sb101001001001011110100110100100110101;
            sine_reg0   <= 36'sb101001100110010110110011111011100101;
        end
        10215: begin
            cosine_reg0 <= 36'sb101001001010000001110010111110100110;
            sine_reg0   <= 36'sb101001100101110010111011000010011111;
        end
        10216: begin
            cosine_reg0 <= 36'sb101001001010100101000000010000101110;
            sine_reg0   <= 36'sb101001100101001111000011000000101100;
        end
        10217: begin
            cosine_reg0 <= 36'sb101001001011001000001110011011001100;
            sine_reg0   <= 36'sb101001100100101011001011110110001101;
        end
        10218: begin
            cosine_reg0 <= 36'sb101001001011101011011101011101111110;
            sine_reg0   <= 36'sb101001100100000111010101100011000100;
        end
        10219: begin
            cosine_reg0 <= 36'sb101001001100001110101101011001000100;
            sine_reg0   <= 36'sb101001100011100011100000000111010001;
        end
        10220: begin
            cosine_reg0 <= 36'sb101001001100110001111110001100011011;
            sine_reg0   <= 36'sb101001100010111111101011100010110111;
        end
        10221: begin
            cosine_reg0 <= 36'sb101001001101010101001111111000000011;
            sine_reg0   <= 36'sb101001100010011011110111110101110110;
        end
        10222: begin
            cosine_reg0 <= 36'sb101001001101111000100010011011111010;
            sine_reg0   <= 36'sb101001100001111000000101000000010001;
        end
        10223: begin
            cosine_reg0 <= 36'sb101001001110011011110101110111111111;
            sine_reg0   <= 36'sb101001100001010100010011000010001000;
        end
        10224: begin
            cosine_reg0 <= 36'sb101001001110111111001010001100010000;
            sine_reg0   <= 36'sb101001100000110000100001111011011100;
        end
        10225: begin
            cosine_reg0 <= 36'sb101001001111100010011111011000101101;
            sine_reg0   <= 36'sb101001100000001100110001101100010000;
        end
        10226: begin
            cosine_reg0 <= 36'sb101001010000000101110101011101010010;
            sine_reg0   <= 36'sb101001011111101001000010010100100101;
        end
        10227: begin
            cosine_reg0 <= 36'sb101001010000101001001100011010000001;
            sine_reg0   <= 36'sb101001011111000101010011110100011011;
        end
        10228: begin
            cosine_reg0 <= 36'sb101001010001001100100100001110110110;
            sine_reg0   <= 36'sb101001011110100001100110001011110101;
        end
        10229: begin
            cosine_reg0 <= 36'sb101001010001101111111100111011110001;
            sine_reg0   <= 36'sb101001011101111101111001011010110011;
        end
        10230: begin
            cosine_reg0 <= 36'sb101001010010010011010110100000110000;
            sine_reg0   <= 36'sb101001011101011010001101100001011000;
        end
        10231: begin
            cosine_reg0 <= 36'sb101001010010110110110000111101110001;
            sine_reg0   <= 36'sb101001011100110110100010011111100100;
        end
        10232: begin
            cosine_reg0 <= 36'sb101001010011011010001100010010110101;
            sine_reg0   <= 36'sb101001011100010010111000010101011000;
        end
        10233: begin
            cosine_reg0 <= 36'sb101001010011111101101000011111111000;
            sine_reg0   <= 36'sb101001011011101111001111000010110111;
        end
        10234: begin
            cosine_reg0 <= 36'sb101001010100100001000101100100111010;
            sine_reg0   <= 36'sb101001011011001011100110101000000010;
        end
        10235: begin
            cosine_reg0 <= 36'sb101001010101000100100011100001111010;
            sine_reg0   <= 36'sb101001011010100111111111000100111001;
        end
        10236: begin
            cosine_reg0 <= 36'sb101001010101101000000010010110110110;
            sine_reg0   <= 36'sb101001011010000100011000011001011111;
        end
        10237: begin
            cosine_reg0 <= 36'sb101001010110001011100010000011101100;
            sine_reg0   <= 36'sb101001011001100000110010100101110101;
        end
        10238: begin
            cosine_reg0 <= 36'sb101001010110101111000010101000011011;
            sine_reg0   <= 36'sb101001011000111101001101101001111011;
        end
        10239: begin
            cosine_reg0 <= 36'sb101001010111010010100100000101000011;
            sine_reg0   <= 36'sb101001011000011001101001100101110100;
        end
        10240: begin
            cosine_reg0 <= 36'sb101001010111110110000110011001100001;
            sine_reg0   <= 36'sb101001010111110110000110011001100001;
        end
        10241: begin
            cosine_reg0 <= 36'sb101001011000011001101001100101110100;
            sine_reg0   <= 36'sb101001010111010010100100000101000011;
        end
        10242: begin
            cosine_reg0 <= 36'sb101001011000111101001101101001111011;
            sine_reg0   <= 36'sb101001010110101111000010101000011011;
        end
        10243: begin
            cosine_reg0 <= 36'sb101001011001100000110010100101110101;
            sine_reg0   <= 36'sb101001010110001011100010000011101100;
        end
        10244: begin
            cosine_reg0 <= 36'sb101001011010000100011000011001011111;
            sine_reg0   <= 36'sb101001010101101000000010010110110110;
        end
        10245: begin
            cosine_reg0 <= 36'sb101001011010100111111111000100111001;
            sine_reg0   <= 36'sb101001010101000100100011100001111010;
        end
        10246: begin
            cosine_reg0 <= 36'sb101001011011001011100110101000000010;
            sine_reg0   <= 36'sb101001010100100001000101100100111010;
        end
        10247: begin
            cosine_reg0 <= 36'sb101001011011101111001111000010110111;
            sine_reg0   <= 36'sb101001010011111101101000011111111000;
        end
        10248: begin
            cosine_reg0 <= 36'sb101001011100010010111000010101011000;
            sine_reg0   <= 36'sb101001010011011010001100010010110101;
        end
        10249: begin
            cosine_reg0 <= 36'sb101001011100110110100010011111100100;
            sine_reg0   <= 36'sb101001010010110110110000111101110001;
        end
        10250: begin
            cosine_reg0 <= 36'sb101001011101011010001101100001011000;
            sine_reg0   <= 36'sb101001010010010011010110100000110000;
        end
        10251: begin
            cosine_reg0 <= 36'sb101001011101111101111001011010110011;
            sine_reg0   <= 36'sb101001010001101111111100111011110001;
        end
        10252: begin
            cosine_reg0 <= 36'sb101001011110100001100110001011110101;
            sine_reg0   <= 36'sb101001010001001100100100001110110110;
        end
        10253: begin
            cosine_reg0 <= 36'sb101001011111000101010011110100011011;
            sine_reg0   <= 36'sb101001010000101001001100011010000001;
        end
        10254: begin
            cosine_reg0 <= 36'sb101001011111101001000010010100100101;
            sine_reg0   <= 36'sb101001010000000101110101011101010010;
        end
        10255: begin
            cosine_reg0 <= 36'sb101001100000001100110001101100010000;
            sine_reg0   <= 36'sb101001001111100010011111011000101101;
        end
        10256: begin
            cosine_reg0 <= 36'sb101001100000110000100001111011011100;
            sine_reg0   <= 36'sb101001001110111111001010001100010000;
        end
        10257: begin
            cosine_reg0 <= 36'sb101001100001010100010011000010001000;
            sine_reg0   <= 36'sb101001001110011011110101110111111111;
        end
        10258: begin
            cosine_reg0 <= 36'sb101001100001111000000101000000010001;
            sine_reg0   <= 36'sb101001001101111000100010011011111010;
        end
        10259: begin
            cosine_reg0 <= 36'sb101001100010011011110111110101110110;
            sine_reg0   <= 36'sb101001001101010101001111111000000011;
        end
        10260: begin
            cosine_reg0 <= 36'sb101001100010111111101011100010110111;
            sine_reg0   <= 36'sb101001001100110001111110001100011011;
        end
        10261: begin
            cosine_reg0 <= 36'sb101001100011100011100000000111010001;
            sine_reg0   <= 36'sb101001001100001110101101011001000100;
        end
        10262: begin
            cosine_reg0 <= 36'sb101001100100000111010101100011000100;
            sine_reg0   <= 36'sb101001001011101011011101011101111110;
        end
        10263: begin
            cosine_reg0 <= 36'sb101001100100101011001011110110001101;
            sine_reg0   <= 36'sb101001001011001000001110011011001100;
        end
        10264: begin
            cosine_reg0 <= 36'sb101001100101001111000011000000101100;
            sine_reg0   <= 36'sb101001001010100101000000010000101110;
        end
        10265: begin
            cosine_reg0 <= 36'sb101001100101110010111011000010011111;
            sine_reg0   <= 36'sb101001001010000001110010111110100110;
        end
        10266: begin
            cosine_reg0 <= 36'sb101001100110010110110011111011100101;
            sine_reg0   <= 36'sb101001001001011110100110100100110101;
        end
        10267: begin
            cosine_reg0 <= 36'sb101001100110111010101101101011111100;
            sine_reg0   <= 36'sb101001001000111011011011000011011101;
        end
        10268: begin
            cosine_reg0 <= 36'sb101001100111011110101000010011100011;
            sine_reg0   <= 36'sb101001001000011000010000011010011111;
        end
        10269: begin
            cosine_reg0 <= 36'sb101001101000000010100011110010011001;
            sine_reg0   <= 36'sb101001000111110101000110101001111101;
        end
        10270: begin
            cosine_reg0 <= 36'sb101001101000100110100000001000011100;
            sine_reg0   <= 36'sb101001000111010001111101110001110111;
        end
        10271: begin
            cosine_reg0 <= 36'sb101001101001001010011101010101101011;
            sine_reg0   <= 36'sb101001000110101110110101110010001111;
        end
        10272: begin
            cosine_reg0 <= 36'sb101001101001101110011011011010000101;
            sine_reg0   <= 36'sb101001000110001011101110101011000110;
        end
        10273: begin
            cosine_reg0 <= 36'sb101001101010010010011010010101100111;
            sine_reg0   <= 36'sb101001000101101000101000011100011110;
        end
        10274: begin
            cosine_reg0 <= 36'sb101001101010110110011010001000010001;
            sine_reg0   <= 36'sb101001000101000101100011000110011001;
        end
        10275: begin
            cosine_reg0 <= 36'sb101001101011011010011010110010000001;
            sine_reg0   <= 36'sb101001000100100010011110101000110110;
        end
        10276: begin
            cosine_reg0 <= 36'sb101001101011111110011100010010110111;
            sine_reg0   <= 36'sb101001000011111111011011000011111001;
        end
        10277: begin
            cosine_reg0 <= 36'sb101001101100100010011110101010101111;
            sine_reg0   <= 36'sb101001000011011100011000010111100010;
        end
        10278: begin
            cosine_reg0 <= 36'sb101001101101000110100001111001101010;
            sine_reg0   <= 36'sb101001000010111001010110100011110010;
        end
        10279: begin
            cosine_reg0 <= 36'sb101001101101101010100101111111100110;
            sine_reg0   <= 36'sb101001000010010110010101101000101011;
        end
        10280: begin
            cosine_reg0 <= 36'sb101001101110001110101010111100100001;
            sine_reg0   <= 36'sb101001000001110011010101100110001110;
        end
        10281: begin
            cosine_reg0 <= 36'sb101001101110110010110000110000011010;
            sine_reg0   <= 36'sb101001000001010000010110011100011101;
        end
        10282: begin
            cosine_reg0 <= 36'sb101001101111010110110111011011001111;
            sine_reg0   <= 36'sb101001000000101101011000001011011001;
        end
        10283: begin
            cosine_reg0 <= 36'sb101001101111111010111110111101000000;
            sine_reg0   <= 36'sb101001000000001010011010110011000011;
        end
        10284: begin
            cosine_reg0 <= 36'sb101001110000011111000111010101101010;
            sine_reg0   <= 36'sb101000111111100111011110010011011101;
        end
        10285: begin
            cosine_reg0 <= 36'sb101001110001000011010000100101001101;
            sine_reg0   <= 36'sb101000111111000100100010101100101000;
        end
        10286: begin
            cosine_reg0 <= 36'sb101001110001100111011010101011100111;
            sine_reg0   <= 36'sb101000111110100001100111111110100101;
        end
        10287: begin
            cosine_reg0 <= 36'sb101001110010001011100101101000110110;
            sine_reg0   <= 36'sb101000111101111110101110001001010101;
        end
        10288: begin
            cosine_reg0 <= 36'sb101001110010101111110001011100111010;
            sine_reg0   <= 36'sb101000111101011011110101001100111011;
        end
        10289: begin
            cosine_reg0 <= 36'sb101001110011010011111110000111110000;
            sine_reg0   <= 36'sb101000111100111000111101001001010111;
        end
        10290: begin
            cosine_reg0 <= 36'sb101001110011111000001011101001011000;
            sine_reg0   <= 36'sb101000111100010110000101111110101011;
        end
        10291: begin
            cosine_reg0 <= 36'sb101001110100011100011010000001110000;
            sine_reg0   <= 36'sb101000111011110011001111101100110111;
        end
        10292: begin
            cosine_reg0 <= 36'sb101001110101000000101001010000110110;
            sine_reg0   <= 36'sb101000111011010000011010010011111110;
        end
        10293: begin
            cosine_reg0 <= 36'sb101001110101100100111001010110101010;
            sine_reg0   <= 36'sb101000111010101101100101110100000001;
        end
        10294: begin
            cosine_reg0 <= 36'sb101001110110001001001010010011001001;
            sine_reg0   <= 36'sb101000111010001010110010001101000001;
        end
        10295: begin
            cosine_reg0 <= 36'sb101001110110101101011100000110010011;
            sine_reg0   <= 36'sb101000111001100111111111011110111111;
        end
        10296: begin
            cosine_reg0 <= 36'sb101001110111010001101110110000000110;
            sine_reg0   <= 36'sb101000111001000101001101101001111101;
        end
        10297: begin
            cosine_reg0 <= 36'sb101001110111110110000010010000100000;
            sine_reg0   <= 36'sb101000111000100010011100101101111100;
        end
        10298: begin
            cosine_reg0 <= 36'sb101001111000011010010110100111100001;
            sine_reg0   <= 36'sb101000110111111111101100101010111110;
        end
        10299: begin
            cosine_reg0 <= 36'sb101001111000111110101011110101000110;
            sine_reg0   <= 36'sb101000110111011100111101100001000011;
        end
        10300: begin
            cosine_reg0 <= 36'sb101001111001100011000001111001001111;
            sine_reg0   <= 36'sb101000110110111010001111010000001101;
        end
        10301: begin
            cosine_reg0 <= 36'sb101001111010000111011000110011111010;
            sine_reg0   <= 36'sb101000110110010111100001111000011110;
        end
        10302: begin
            cosine_reg0 <= 36'sb101001111010101011110000100101000110;
            sine_reg0   <= 36'sb101000110101110100110101011001110111;
        end
        10303: begin
            cosine_reg0 <= 36'sb101001111011010000001001001100110001;
            sine_reg0   <= 36'sb101000110101010010001001110100011001;
        end
        10304: begin
            cosine_reg0 <= 36'sb101001111011110100100010101010111001;
            sine_reg0   <= 36'sb101000110100101111011111001000000101;
        end
        10305: begin
            cosine_reg0 <= 36'sb101001111100011000111100111111011110;
            sine_reg0   <= 36'sb101000110100001100110101010100111101;
        end
        10306: begin
            cosine_reg0 <= 36'sb101001111100111101011000001010011110;
            sine_reg0   <= 36'sb101000110011101010001100011011000010;
        end
        10307: begin
            cosine_reg0 <= 36'sb101001111101100001110100001011111000;
            sine_reg0   <= 36'sb101000110011000111100100011010010101;
        end
        10308: begin
            cosine_reg0 <= 36'sb101001111110000110010001000011101010;
            sine_reg0   <= 36'sb101000110010100100111101010010111001;
        end
        10309: begin
            cosine_reg0 <= 36'sb101001111110101010101110110001110011;
            sine_reg0   <= 36'sb101000110010000010010111000100101101;
        end
        10310: begin
            cosine_reg0 <= 36'sb101001111111001111001101010110010001;
            sine_reg0   <= 36'sb101000110001011111110001101111110100;
        end
        10311: begin
            cosine_reg0 <= 36'sb101001111111110011101100110001000011;
            sine_reg0   <= 36'sb101000110000111101001101010100001111;
        end
        10312: begin
            cosine_reg0 <= 36'sb101010000000011000001101000010000111;
            sine_reg0   <= 36'sb101000110000011010101001110001111111;
        end
        10313: begin
            cosine_reg0 <= 36'sb101010000000111100101110001001011101;
            sine_reg0   <= 36'sb101000101111111000000111001001000101;
        end
        10314: begin
            cosine_reg0 <= 36'sb101010000001100001010000000111000011;
            sine_reg0   <= 36'sb101000101111010101100101011001100011;
        end
        10315: begin
            cosine_reg0 <= 36'sb101010000010000101110010111010110111;
            sine_reg0   <= 36'sb101000101110110011000100100011011011;
        end
        10316: begin
            cosine_reg0 <= 36'sb101010000010101010010110100100110111;
            sine_reg0   <= 36'sb101000101110010000100100100110101100;
        end
        10317: begin
            cosine_reg0 <= 36'sb101010000011001110111011000101000100;
            sine_reg0   <= 36'sb101000101101101110000101100011011010;
        end
        10318: begin
            cosine_reg0 <= 36'sb101010000011110011100000011011011010;
            sine_reg0   <= 36'sb101000101101001011100111011001100101;
        end
        10319: begin
            cosine_reg0 <= 36'sb101010000100011000000110100111111001;
            sine_reg0   <= 36'sb101000101100101001001010001001001110;
        end
        10320: begin
            cosine_reg0 <= 36'sb101010000100111100101101101010100000;
            sine_reg0   <= 36'sb101000101100000110101101110010010111;
        end
        10321: begin
            cosine_reg0 <= 36'sb101010000101100001010101100011001100;
            sine_reg0   <= 36'sb101000101011100100010010010101000000;
        end
        10322: begin
            cosine_reg0 <= 36'sb101010000110000101111110010001111101;
            sine_reg0   <= 36'sb101000101011000001110111110001001101;
        end
        10323: begin
            cosine_reg0 <= 36'sb101010000110101010100111110110110001;
            sine_reg0   <= 36'sb101000101010011111011110000110111101;
        end
        10324: begin
            cosine_reg0 <= 36'sb101010000111001111010010010001100111;
            sine_reg0   <= 36'sb101000101001111101000101010110010010;
        end
        10325: begin
            cosine_reg0 <= 36'sb101010000111110011111101100010011100;
            sine_reg0   <= 36'sb101000101001011010101101011111001110;
        end
        10326: begin
            cosine_reg0 <= 36'sb101010001000011000101001101001010001;
            sine_reg0   <= 36'sb101000101000111000010110100001110001;
        end
        10327: begin
            cosine_reg0 <= 36'sb101010001000111101010110100110000011;
            sine_reg0   <= 36'sb101000101000010110000000011101111110;
        end
        10328: begin
            cosine_reg0 <= 36'sb101010001001100010000100011000110001;
            sine_reg0   <= 36'sb101000100111110011101011010011110101;
        end
        10329: begin
            cosine_reg0 <= 36'sb101010001010000110110011000001011010;
            sine_reg0   <= 36'sb101000100111010001010111000011010111;
        end
        10330: begin
            cosine_reg0 <= 36'sb101010001010101011100010011111111100;
            sine_reg0   <= 36'sb101000100110101111000011101100100111;
        end
        10331: begin
            cosine_reg0 <= 36'sb101010001011010000010010110100010101;
            sine_reg0   <= 36'sb101000100110001100110001001111100101;
        end
        10332: begin
            cosine_reg0 <= 36'sb101010001011110101000011111110100101;
            sine_reg0   <= 36'sb101000100101101010011111101100010010;
        end
        10333: begin
            cosine_reg0 <= 36'sb101010001100011001110101111110101010;
            sine_reg0   <= 36'sb101000100101001000001111000010110001;
        end
        10334: begin
            cosine_reg0 <= 36'sb101010001100111110101000110100100010;
            sine_reg0   <= 36'sb101000100100100101111111010011000010;
        end
        10335: begin
            cosine_reg0 <= 36'sb101010001101100011011100100000001100;
            sine_reg0   <= 36'sb101000100100000011110000011101000110;
        end
        10336: begin
            cosine_reg0 <= 36'sb101010001110001000010001000001100111;
            sine_reg0   <= 36'sb101000100011100001100010100001000000;
        end
        10337: begin
            cosine_reg0 <= 36'sb101010001110101101000110011000110010;
            sine_reg0   <= 36'sb101000100010111111010101011110110000;
        end
        10338: begin
            cosine_reg0 <= 36'sb101010001111010001111100100101101010;
            sine_reg0   <= 36'sb101000100010011101001001010110010111;
        end
        10339: begin
            cosine_reg0 <= 36'sb101010001111110110110011101000001110;
            sine_reg0   <= 36'sb101000100001111010111110000111110111;
        end
        10340: begin
            cosine_reg0 <= 36'sb101010010000011011101011100000011110;
            sine_reg0   <= 36'sb101000100001011000110011110011010010;
        end
        10341: begin
            cosine_reg0 <= 36'sb101010010001000000100100001110010111;
            sine_reg0   <= 36'sb101000100000110110101010011000101000;
        end
        10342: begin
            cosine_reg0 <= 36'sb101010010001100101011101110001111000;
            sine_reg0   <= 36'sb101000100000010100100001110111111011;
        end
        10343: begin
            cosine_reg0 <= 36'sb101010010010001010011000001011000000;
            sine_reg0   <= 36'sb101000011111110010011010010001001100;
        end
        10344: begin
            cosine_reg0 <= 36'sb101010010010101111010011011001101101;
            sine_reg0   <= 36'sb101000011111010000010011100100011101;
        end
        10345: begin
            cosine_reg0 <= 36'sb101010010011010100001111011101111110;
            sine_reg0   <= 36'sb101000011110101110001101110001101110;
        end
        10346: begin
            cosine_reg0 <= 36'sb101010010011111001001100010111110001;
            sine_reg0   <= 36'sb101000011110001100001000111001000010;
        end
        10347: begin
            cosine_reg0 <= 36'sb101010010100011110001010000111000110;
            sine_reg0   <= 36'sb101000011101101010000100111010011000;
        end
        10348: begin
            cosine_reg0 <= 36'sb101010010101000011001000101011111010;
            sine_reg0   <= 36'sb101000011101001000000001110101110100;
        end
        10349: begin
            cosine_reg0 <= 36'sb101010010101101000001000000110001100;
            sine_reg0   <= 36'sb101000011100100101111111101011010110;
        end
        10350: begin
            cosine_reg0 <= 36'sb101010010110001101001000010101111011;
            sine_reg0   <= 36'sb101000011100000011111110011010111111;
        end
        10351: begin
            cosine_reg0 <= 36'sb101010010110110010001001011011000101;
            sine_reg0   <= 36'sb101000011011100001111110000100110001;
        end
        10352: begin
            cosine_reg0 <= 36'sb101010010111010111001011010101101001;
            sine_reg0   <= 36'sb101000011010111111111110101000101101;
        end
        10353: begin
            cosine_reg0 <= 36'sb101010010111111100001110000101100110;
            sine_reg0   <= 36'sb101000011010011110000000000110110100;
        end
        10354: begin
            cosine_reg0 <= 36'sb101010011000100001010001101010111010;
            sine_reg0   <= 36'sb101000011001111100000010011111001000;
        end
        10355: begin
            cosine_reg0 <= 36'sb101010011001000110010110000101100011;
            sine_reg0   <= 36'sb101000011001011010000101110001101010;
        end
        10356: begin
            cosine_reg0 <= 36'sb101010011001101011011011010101100000;
            sine_reg0   <= 36'sb101000011000111000001001111110011011;
        end
        10357: begin
            cosine_reg0 <= 36'sb101010011010010000100001011010110000;
            sine_reg0   <= 36'sb101000011000010110001111000101011100;
        end
        10358: begin
            cosine_reg0 <= 36'sb101010011010110101101000010101010010;
            sine_reg0   <= 36'sb101000010111110100010101000110101111;
        end
        10359: begin
            cosine_reg0 <= 36'sb101010011011011010110000000101000011;
            sine_reg0   <= 36'sb101000010111010010011100000010010110;
        end
        10360: begin
            cosine_reg0 <= 36'sb101010011011111111111000101010000011;
            sine_reg0   <= 36'sb101000010110110000100011111000010001;
        end
        10361: begin
            cosine_reg0 <= 36'sb101010011100100101000010000100010000;
            sine_reg0   <= 36'sb101000010110001110101100101000100010;
        end
        10362: begin
            cosine_reg0 <= 36'sb101010011101001010001100010011101000;
            sine_reg0   <= 36'sb101000010101101100110110010011001001;
        end
        10363: begin
            cosine_reg0 <= 36'sb101010011101101111010111011000001011;
            sine_reg0   <= 36'sb101000010101001011000000111000001010;
        end
        10364: begin
            cosine_reg0 <= 36'sb101010011110010100100011010001110110;
            sine_reg0   <= 36'sb101000010100101001001100010111100100;
        end
        10365: begin
            cosine_reg0 <= 36'sb101010011110111001110000000000101000;
            sine_reg0   <= 36'sb101000010100000111011000110001011000;
        end
        10366: begin
            cosine_reg0 <= 36'sb101010011111011110111101100100100001;
            sine_reg0   <= 36'sb101000010011100101100110000101101010;
        end
        10367: begin
            cosine_reg0 <= 36'sb101010100000000100001011111101011110;
            sine_reg0   <= 36'sb101000010011000011110100010100011000;
        end
        10368: begin
            cosine_reg0 <= 36'sb101010100000101001011011001011011101;
            sine_reg0   <= 36'sb101000010010100010000011011101100110;
        end
        10369: begin
            cosine_reg0 <= 36'sb101010100001001110101011001110011111;
            sine_reg0   <= 36'sb101000010010000000010011100001010100;
        end
        10370: begin
            cosine_reg0 <= 36'sb101010100001110011111100000110100000;
            sine_reg0   <= 36'sb101000010001011110100100011111100011;
        end
        10371: begin
            cosine_reg0 <= 36'sb101010100010011001001101110011100000;
            sine_reg0   <= 36'sb101000010000111100110110011000010110;
        end
        10372: begin
            cosine_reg0 <= 36'sb101010100010111110100000010101011110;
            sine_reg0   <= 36'sb101000010000011011001001001011101100;
        end
        10373: begin
            cosine_reg0 <= 36'sb101010100011100011110011101100010111;
            sine_reg0   <= 36'sb101000001111111001011100111001101000;
        end
        10374: begin
            cosine_reg0 <= 36'sb101010100100001001000111111000001010;
            sine_reg0   <= 36'sb101000001111010111110001100010001010;
        end
        10375: begin
            cosine_reg0 <= 36'sb101010100100101110011100111000110111;
            sine_reg0   <= 36'sb101000001110110110000111000101010100;
        end
        10376: begin
            cosine_reg0 <= 36'sb101010100101010011110010101110011011;
            sine_reg0   <= 36'sb101000001110010100011101100011001000;
        end
        10377: begin
            cosine_reg0 <= 36'sb101010100101111001001001011000110101;
            sine_reg0   <= 36'sb101000001101110010110100111011100110;
        end
        10378: begin
            cosine_reg0 <= 36'sb101010100110011110100000111000000011;
            sine_reg0   <= 36'sb101000001101010001001101001110110001;
        end
        10379: begin
            cosine_reg0 <= 36'sb101010100111000011111001001100000101;
            sine_reg0   <= 36'sb101000001100101111100110011100101000;
        end
        10380: begin
            cosine_reg0 <= 36'sb101010100111101001010010010100111001;
            sine_reg0   <= 36'sb101000001100001110000000100101001110;
        end
        10381: begin
            cosine_reg0 <= 36'sb101010101000001110101100010010011100;
            sine_reg0   <= 36'sb101000001011101100011011101000100011;
        end
        10382: begin
            cosine_reg0 <= 36'sb101010101000110100000111000100101111;
            sine_reg0   <= 36'sb101000001011001010110111100110101010;
        end
        10383: begin
            cosine_reg0 <= 36'sb101010101001011001100010101011101111;
            sine_reg0   <= 36'sb101000001010101001010100011111100011;
        end
        10384: begin
            cosine_reg0 <= 36'sb101010101001111110111111000111011011;
            sine_reg0   <= 36'sb101000001010000111110010010011010000;
        end
        10385: begin
            cosine_reg0 <= 36'sb101010101010100100011100010111110001;
            sine_reg0   <= 36'sb101000001001100110010001000001110010;
        end
        10386: begin
            cosine_reg0 <= 36'sb101010101011001001111010011100110001;
            sine_reg0   <= 36'sb101000001001000100110000101011001010;
        end
        10387: begin
            cosine_reg0 <= 36'sb101010101011101111011001010110011000;
            sine_reg0   <= 36'sb101000001000100011010001001111011001;
        end
        10388: begin
            cosine_reg0 <= 36'sb101010101100010100111001000100100101;
            sine_reg0   <= 36'sb101000001000000001110010101110100001;
        end
        10389: begin
            cosine_reg0 <= 36'sb101010101100111010011001100111010111;
            sine_reg0   <= 36'sb101000000111100000010101001000100100;
        end
        10390: begin
            cosine_reg0 <= 36'sb101010101101011111111010111110101101;
            sine_reg0   <= 36'sb101000000110111110111000011101100010;
        end
        10391: begin
            cosine_reg0 <= 36'sb101010101110000101011101001010100100;
            sine_reg0   <= 36'sb101000000110011101011100101101011100;
        end
        10392: begin
            cosine_reg0 <= 36'sb101010101110101011000000001010111011;
            sine_reg0   <= 36'sb101000000101111100000001111000010101;
        end
        10393: begin
            cosine_reg0 <= 36'sb101010101111010000100011111111110010;
            sine_reg0   <= 36'sb101000000101011010100111111110001100;
        end
        10394: begin
            cosine_reg0 <= 36'sb101010101111110110001000101001000110;
            sine_reg0   <= 36'sb101000000100111001001110111111000101;
        end
        10395: begin
            cosine_reg0 <= 36'sb101010110000011011101110000110110110;
            sine_reg0   <= 36'sb101000000100010111110110111010111111;
        end
        10396: begin
            cosine_reg0 <= 36'sb101010110001000001010100011001000000;
            sine_reg0   <= 36'sb101000000011110110011111110001111100;
        end
        10397: begin
            cosine_reg0 <= 36'sb101010110001100110111011011111100100;
            sine_reg0   <= 36'sb101000000011010101001001100011111110;
        end
        10398: begin
            cosine_reg0 <= 36'sb101010110010001100100011011010100000;
            sine_reg0   <= 36'sb101000000010110011110100010001000110;
        end
        10399: begin
            cosine_reg0 <= 36'sb101010110010110010001100001001110001;
            sine_reg0   <= 36'sb101000000010010010011111111001010100;
        end
        10400: begin
            cosine_reg0 <= 36'sb101010110011010111110101101101011000;
            sine_reg0   <= 36'sb101000000001110001001100011100101011;
        end
        10401: begin
            cosine_reg0 <= 36'sb101010110011111101100000000101010010;
            sine_reg0   <= 36'sb101000000001001111111001111011001011;
        end
        10402: begin
            cosine_reg0 <= 36'sb101010110100100011001011010001011101;
            sine_reg0   <= 36'sb101000000000101110101000010100110110;
        end
        10403: begin
            cosine_reg0 <= 36'sb101010110101001000110111010001111010;
            sine_reg0   <= 36'sb101000000000001101010111101001101110;
        end
        10404: begin
            cosine_reg0 <= 36'sb101010110101101110100100000110100101;
            sine_reg0   <= 36'sb100111111111101100000111111001110011;
        end
        10405: begin
            cosine_reg0 <= 36'sb101010110110010100010001101111011101;
            sine_reg0   <= 36'sb100111111111001010111001000101000110;
        end
        10406: begin
            cosine_reg0 <= 36'sb101010110110111010000000001100100010;
            sine_reg0   <= 36'sb100111111110101001101011001011101001;
        end
        10407: begin
            cosine_reg0 <= 36'sb101010110111011111101111011101110010;
            sine_reg0   <= 36'sb100111111110001000011110001101011110;
        end
        10408: begin
            cosine_reg0 <= 36'sb101010111000000101011111100011001010;
            sine_reg0   <= 36'sb100111111101100111010010001010100101;
        end
        10409: begin
            cosine_reg0 <= 36'sb101010111000101011010000011100101011;
            sine_reg0   <= 36'sb100111111101000110000111000011000000;
        end
        10410: begin
            cosine_reg0 <= 36'sb101010111001010001000010001010010001;
            sine_reg0   <= 36'sb100111111100100100111100110110110000;
        end
        10411: begin
            cosine_reg0 <= 36'sb101010111001110110110100101011111100;
            sine_reg0   <= 36'sb100111111100000011110011100101110111;
        end
        10412: begin
            cosine_reg0 <= 36'sb101010111010011100101000000001101011;
            sine_reg0   <= 36'sb100111111011100010101011010000010101;
        end
        10413: begin
            cosine_reg0 <= 36'sb101010111011000010011100001011011100;
            sine_reg0   <= 36'sb100111111011000001100011110110001100;
        end
        10414: begin
            cosine_reg0 <= 36'sb101010111011101000010001001001001101;
            sine_reg0   <= 36'sb100111111010100000011101010111011101;
        end
        10415: begin
            cosine_reg0 <= 36'sb101010111100001110000110111010111101;
            sine_reg0   <= 36'sb100111111001111111010111110100001010;
        end
        10416: begin
            cosine_reg0 <= 36'sb101010111100110011111101100000101010;
            sine_reg0   <= 36'sb100111111001011110010011001100010011;
        end
        10417: begin
            cosine_reg0 <= 36'sb101010111101011001110100111010010100;
            sine_reg0   <= 36'sb100111111000111101001111011111111011;
        end
        10418: begin
            cosine_reg0 <= 36'sb101010111101111111101101000111111000;
            sine_reg0   <= 36'sb100111111000011100001100101111000010;
        end
        10419: begin
            cosine_reg0 <= 36'sb101010111110100101100110001001010101;
            sine_reg0   <= 36'sb100111110111111011001010111001101001;
        end
        10420: begin
            cosine_reg0 <= 36'sb101010111111001011011111111110101010;
            sine_reg0   <= 36'sb100111110111011010001001111111110010;
        end
        10421: begin
            cosine_reg0 <= 36'sb101010111111110001011010100111110101;
            sine_reg0   <= 36'sb100111110110111001001010000001011111;
        end
        10422: begin
            cosine_reg0 <= 36'sb101011000000010111010110000100110101;
            sine_reg0   <= 36'sb100111110110011000001010111110110000;
        end
        10423: begin
            cosine_reg0 <= 36'sb101011000000111101010010010101101000;
            sine_reg0   <= 36'sb100111110101110111001100110111100110;
        end
        10424: begin
            cosine_reg0 <= 36'sb101011000001100011001111011010001101;
            sine_reg0   <= 36'sb100111110101010110001111101100000011;
        end
        10425: begin
            cosine_reg0 <= 36'sb101011000010001001001101010010100011;
            sine_reg0   <= 36'sb100111110100110101010011011100001001;
        end
        10426: begin
            cosine_reg0 <= 36'sb101011000010101111001011111110100111;
            sine_reg0   <= 36'sb100111110100010100011000000111111000;
        end
        10427: begin
            cosine_reg0 <= 36'sb101011000011010101001011011110011001;
            sine_reg0   <= 36'sb100111110011110011011101101111010010;
        end
        10428: begin
            cosine_reg0 <= 36'sb101011000011111011001011110001110111;
            sine_reg0   <= 36'sb100111110011010010100100010010011000;
        end
        10429: begin
            cosine_reg0 <= 36'sb101011000100100001001100111000111111;
            sine_reg0   <= 36'sb100111110010110001101011110001001011;
        end
        10430: begin
            cosine_reg0 <= 36'sb101011000101000111001110110011110000;
            sine_reg0   <= 36'sb100111110010010000110100001011101101;
        end
        10431: begin
            cosine_reg0 <= 36'sb101011000101101101010001100010001001;
            sine_reg0   <= 36'sb100111110001101111111101100001111110;
        end
        10432: begin
            cosine_reg0 <= 36'sb101011000110010011010101000100001000;
            sine_reg0   <= 36'sb100111110001001111000111110100000001;
        end
        10433: begin
            cosine_reg0 <= 36'sb101011000110111001011001011001101011;
            sine_reg0   <= 36'sb100111110000101110010011000001110110;
        end
        10434: begin
            cosine_reg0 <= 36'sb101011000111011111011110100010110010;
            sine_reg0   <= 36'sb100111110000001101011111001011011110;
        end
        10435: begin
            cosine_reg0 <= 36'sb101011001000000101100100011111011010;
            sine_reg0   <= 36'sb100111101111101100101100010000111100;
        end
        10436: begin
            cosine_reg0 <= 36'sb101011001000101011101011001111100011;
            sine_reg0   <= 36'sb100111101111001011111010010010010000;
        end
        10437: begin
            cosine_reg0 <= 36'sb101011001001010001110010110011001010;
            sine_reg0   <= 36'sb100111101110101011001001001111011011;
        end
        10438: begin
            cosine_reg0 <= 36'sb101011001001110111111011001010001111;
            sine_reg0   <= 36'sb100111101110001010011001001000011110;
        end
        10439: begin
            cosine_reg0 <= 36'sb101011001010011110000100010100110000;
            sine_reg0   <= 36'sb100111101101101001101001111101011100;
        end
        10440: begin
            cosine_reg0 <= 36'sb101011001011000100001110010010101010;
            sine_reg0   <= 36'sb100111101101001000111011101110010101;
        end
        10441: begin
            cosine_reg0 <= 36'sb101011001011101010011001000011111110;
            sine_reg0   <= 36'sb100111101100101000001110011011001010;
        end
        10442: begin
            cosine_reg0 <= 36'sb101011001100010000100100101000101001;
            sine_reg0   <= 36'sb100111101100000111100010000011111101;
        end
        10443: begin
            cosine_reg0 <= 36'sb101011001100110110110001000000101011;
            sine_reg0   <= 36'sb100111101011100110110110101000101111;
        end
        10444: begin
            cosine_reg0 <= 36'sb101011001101011100111110001100000000;
            sine_reg0   <= 36'sb100111101011000110001100001001100010;
        end
        10445: begin
            cosine_reg0 <= 36'sb101011001110000011001100001010101001;
            sine_reg0   <= 36'sb100111101010100101100010100110010101;
        end
        10446: begin
            cosine_reg0 <= 36'sb101011001110101001011010111100100011;
            sine_reg0   <= 36'sb100111101010000100111001111111001100;
        end
        10447: begin
            cosine_reg0 <= 36'sb101011001111001111101010100001101101;
            sine_reg0   <= 36'sb100111101001100100010010010100000111;
        end
        10448: begin
            cosine_reg0 <= 36'sb101011001111110101111010111010000110;
            sine_reg0   <= 36'sb100111101001000011101011100101000110;
        end
        10449: begin
            cosine_reg0 <= 36'sb101011010000011100001100000101101011;
            sine_reg0   <= 36'sb100111101000100011000101110010001101;
        end
        10450: begin
            cosine_reg0 <= 36'sb101011010001000010011110000100011101;
            sine_reg0   <= 36'sb100111101000000010100000111011011011;
        end
        10451: begin
            cosine_reg0 <= 36'sb101011010001101000110000110110011000;
            sine_reg0   <= 36'sb100111100111100001111101000000110010;
        end
        10452: begin
            cosine_reg0 <= 36'sb101011010010001111000100011011011101;
            sine_reg0   <= 36'sb100111100111000001011010000010010100;
        end
        10453: begin
            cosine_reg0 <= 36'sb101011010010110101011000110011101000;
            sine_reg0   <= 36'sb100111100110100000111000000000000001;
        end
        10454: begin
            cosine_reg0 <= 36'sb101011010011011011101101111110111001;
            sine_reg0   <= 36'sb100111100110000000010110111001111011;
        end
        10455: begin
            cosine_reg0 <= 36'sb101011010100000010000011111101001111;
            sine_reg0   <= 36'sb100111100101011111110110110000000011;
        end
        10456: begin
            cosine_reg0 <= 36'sb101011010100101000011010101110100111;
            sine_reg0   <= 36'sb100111100100111111010111100010011010;
        end
        10457: begin
            cosine_reg0 <= 36'sb101011010101001110110010010011000000;
            sine_reg0   <= 36'sb100111100100011110111001010001000010;
        end
        10458: begin
            cosine_reg0 <= 36'sb101011010101110101001010101010011010;
            sine_reg0   <= 36'sb100111100011111110011011111011111100;
        end
        10459: begin
            cosine_reg0 <= 36'sb101011010110011011100011110100110001;
            sine_reg0   <= 36'sb100111100011011101111111100011001000;
        end
        10460: begin
            cosine_reg0 <= 36'sb101011010111000001111101110010000101;
            sine_reg0   <= 36'sb100111100010111101100100000110101010;
        end
        10461: begin
            cosine_reg0 <= 36'sb101011010111101000011000100010010101;
            sine_reg0   <= 36'sb100111100010011101001001100110100000;
        end
        10462: begin
            cosine_reg0 <= 36'sb101011011000001110110100000101011111;
            sine_reg0   <= 36'sb100111100001111100110000000010101110;
        end
        10463: begin
            cosine_reg0 <= 36'sb101011011000110101010000011011100001;
            sine_reg0   <= 36'sb100111100001011100010111011011010011;
        end
        10464: begin
            cosine_reg0 <= 36'sb101011011001011011101101100100011010;
            sine_reg0   <= 36'sb100111100000111011111111110000010010;
        end
        10465: begin
            cosine_reg0 <= 36'sb101011011010000010001011100000001000;
            sine_reg0   <= 36'sb100111100000011011101001000001101100;
        end
        10466: begin
            cosine_reg0 <= 36'sb101011011010101000101010001110101011;
            sine_reg0   <= 36'sb100111011111111011010011001111100001;
        end
        10467: begin
            cosine_reg0 <= 36'sb101011011011001111001001101111111111;
            sine_reg0   <= 36'sb100111011111011010111110011001110011;
        end
        10468: begin
            cosine_reg0 <= 36'sb101011011011110101101010000100000101;
            sine_reg0   <= 36'sb100111011110111010101010100000100100;
        end
        10469: begin
            cosine_reg0 <= 36'sb101011011100011100001011001010111010;
            sine_reg0   <= 36'sb100111011110011010010111100011110100;
        end
        10470: begin
            cosine_reg0 <= 36'sb101011011101000010101101000100011110;
            sine_reg0   <= 36'sb100111011101111010000101100011100101;
        end
        10471: begin
            cosine_reg0 <= 36'sb101011011101101001001111110000101110;
            sine_reg0   <= 36'sb100111011101011001110100011111111000;
        end
        10472: begin
            cosine_reg0 <= 36'sb101011011110001111110011001111101000;
            sine_reg0   <= 36'sb100111011100111001100100011000101111;
        end
        10473: begin
            cosine_reg0 <= 36'sb101011011110110110010111100001001101;
            sine_reg0   <= 36'sb100111011100011001010101001110001010;
        end
        10474: begin
            cosine_reg0 <= 36'sb101011011111011100111100100101011001;
            sine_reg0   <= 36'sb100111011011111001000111000000001010;
        end
        10475: begin
            cosine_reg0 <= 36'sb101011100000000011100010011100001101;
            sine_reg0   <= 36'sb100111011011011000111001101110110010;
        end
        10476: begin
            cosine_reg0 <= 36'sb101011100000101010001001000101100101;
            sine_reg0   <= 36'sb100111011010111000101101011010000010;
        end
        10477: begin
            cosine_reg0 <= 36'sb101011100001010000110000100001100000;
            sine_reg0   <= 36'sb100111011010011000100010000001111011;
        end
        10478: begin
            cosine_reg0 <= 36'sb101011100001110111011000101111111110;
            sine_reg0   <= 36'sb100111011001111000010111100110100000;
        end
        10479: begin
            cosine_reg0 <= 36'sb101011100010011110000001110000111101;
            sine_reg0   <= 36'sb100111011001011000001110000111110000;
        end
        10480: begin
            cosine_reg0 <= 36'sb101011100011000100101011100100011011;
            sine_reg0   <= 36'sb100111011000111000000101100101101101;
        end
        10481: begin
            cosine_reg0 <= 36'sb101011100011101011010110001010010110;
            sine_reg0   <= 36'sb100111011000010111111110000000011001;
        end
        10482: begin
            cosine_reg0 <= 36'sb101011100100010010000001100010101101;
            sine_reg0   <= 36'sb100111010111110111110111010111110101;
        end
        10483: begin
            cosine_reg0 <= 36'sb101011100100111000101101101101011111;
            sine_reg0   <= 36'sb100111010111010111110001101100000001;
        end
        10484: begin
            cosine_reg0 <= 36'sb101011100101011111011010101010101011;
            sine_reg0   <= 36'sb100111010110110111101100111101000000;
        end
        10485: begin
            cosine_reg0 <= 36'sb101011100110000110001000011010001110;
            sine_reg0   <= 36'sb100111010110010111101001001010110010;
        end
        10486: begin
            cosine_reg0 <= 36'sb101011100110101100110110111100000111;
            sine_reg0   <= 36'sb100111010101110111100110010101011001;
        end
        10487: begin
            cosine_reg0 <= 36'sb101011100111010011100110010000010101;
            sine_reg0   <= 36'sb100111010101010111100100011100110101;
        end
        10488: begin
            cosine_reg0 <= 36'sb101011100111111010010110010110110110;
            sine_reg0   <= 36'sb100111010100110111100011100001001001;
        end
        10489: begin
            cosine_reg0 <= 36'sb101011101000100001000111001111101001;
            sine_reg0   <= 36'sb100111010100010111100011100010010101;
        end
        10490: begin
            cosine_reg0 <= 36'sb101011101001000111111000111010101100;
            sine_reg0   <= 36'sb100111010011110111100100100000011011;
        end
        10491: begin
            cosine_reg0 <= 36'sb101011101001101110101011010111111101;
            sine_reg0   <= 36'sb100111010011010111100110011011011100;
        end
        10492: begin
            cosine_reg0 <= 36'sb101011101010010101011110100111011100;
            sine_reg0   <= 36'sb100111010010110111101001010011011000;
        end
        10493: begin
            cosine_reg0 <= 36'sb101011101010111100010010101001000111;
            sine_reg0   <= 36'sb100111010010010111101101001000010010;
        end
        10494: begin
            cosine_reg0 <= 36'sb101011101011100011000111011100111100;
            sine_reg0   <= 36'sb100111010001110111110001111010001010;
        end
        10495: begin
            cosine_reg0 <= 36'sb101011101100001001111101000010111001;
            sine_reg0   <= 36'sb100111010001010111110111101001000010;
        end
        10496: begin
            cosine_reg0 <= 36'sb101011101100110000110011011010111110;
            sine_reg0   <= 36'sb100111010000110111111110010100111100;
        end
        10497: begin
            cosine_reg0 <= 36'sb101011101101010111101010100101001001;
            sine_reg0   <= 36'sb100111010000011000000101111101110111;
        end
        10498: begin
            cosine_reg0 <= 36'sb101011101101111110100010100001011000;
            sine_reg0   <= 36'sb100111001111111000001110100011110110;
        end
        10499: begin
            cosine_reg0 <= 36'sb101011101110100101011011001111101001;
            sine_reg0   <= 36'sb100111001111011000011000000110111001;
        end
        10500: begin
            cosine_reg0 <= 36'sb101011101111001100010100101111111100;
            sine_reg0   <= 36'sb100111001110111000100010100111000010;
        end
        10501: begin
            cosine_reg0 <= 36'sb101011101111110011001111000010001111;
            sine_reg0   <= 36'sb100111001110011000101110000100010011;
        end
        10502: begin
            cosine_reg0 <= 36'sb101011110000011010001010000110100000;
            sine_reg0   <= 36'sb100111001101111000111010011110101011;
        end
        10503: begin
            cosine_reg0 <= 36'sb101011110001000001000101111100101101;
            sine_reg0   <= 36'sb100111001101011001000111110110001110;
        end
        10504: begin
            cosine_reg0 <= 36'sb101011110001101000000010100100110110;
            sine_reg0   <= 36'sb100111001100111001010110001010111011;
        end
        10505: begin
            cosine_reg0 <= 36'sb101011110010001110111111111110111001;
            sine_reg0   <= 36'sb100111001100011001100101011100110100;
        end
        10506: begin
            cosine_reg0 <= 36'sb101011110010110101111110001010110011;
            sine_reg0   <= 36'sb100111001011111001110101101011111010;
        end
        10507: begin
            cosine_reg0 <= 36'sb101011110011011100111101001000100101;
            sine_reg0   <= 36'sb100111001011011010000110111000001111;
        end
        10508: begin
            cosine_reg0 <= 36'sb101011110100000011111100111000001100;
            sine_reg0   <= 36'sb100111001010111010011001000001110100;
        end
        10509: begin
            cosine_reg0 <= 36'sb101011110100101010111101011001100110;
            sine_reg0   <= 36'sb100111001010011010101100001000101001;
        end
        10510: begin
            cosine_reg0 <= 36'sb101011110101010001111110101100110011;
            sine_reg0   <= 36'sb100111001001111011000000001100110001;
        end
        10511: begin
            cosine_reg0 <= 36'sb101011110101111001000000110001110000;
            sine_reg0   <= 36'sb100111001001011011010101001110001100;
        end
        10512: begin
            cosine_reg0 <= 36'sb101011110110100000000011101000011101;
            sine_reg0   <= 36'sb100111001000111011101011001100111011;
        end
        10513: begin
            cosine_reg0 <= 36'sb101011110111000111000111010000110111;
            sine_reg0   <= 36'sb100111001000011100000010001001000000;
        end
        10514: begin
            cosine_reg0 <= 36'sb101011110111101110001011101010111110;
            sine_reg0   <= 36'sb100111000111111100011010000010011101;
        end
        10515: begin
            cosine_reg0 <= 36'sb101011111000010101010000110110101111;
            sine_reg0   <= 36'sb100111000111011100110010111001010001;
        end
        10516: begin
            cosine_reg0 <= 36'sb101011111000111100010110110100001010;
            sine_reg0   <= 36'sb100111000110111101001100101101011111;
        end
        10517: begin
            cosine_reg0 <= 36'sb101011111001100011011101100011001100;
            sine_reg0   <= 36'sb100111000110011101100111011111001000;
        end
        10518: begin
            cosine_reg0 <= 36'sb101011111010001010100101000011110100;
            sine_reg0   <= 36'sb100111000101111110000011001110001101;
        end
        10519: begin
            cosine_reg0 <= 36'sb101011111010110001101101010110000001;
            sine_reg0   <= 36'sb100111000101011110011111111010101111;
        end
        10520: begin
            cosine_reg0 <= 36'sb101011111011011000110110011001110001;
            sine_reg0   <= 36'sb100111000100111110111101100100101111;
        end
        10521: begin
            cosine_reg0 <= 36'sb101011111100000000000000001111000011;
            sine_reg0   <= 36'sb100111000100011111011100001100001110;
        end
        10522: begin
            cosine_reg0 <= 36'sb101011111100100111001010110101110101;
            sine_reg0   <= 36'sb100111000011111111111011110001001111;
        end
        10523: begin
            cosine_reg0 <= 36'sb101011111101001110010110001110000110;
            sine_reg0   <= 36'sb100111000011100000011100010011110001;
        end
        10524: begin
            cosine_reg0 <= 36'sb101011111101110101100010010111110011;
            sine_reg0   <= 36'sb100111000011000000111101110011110111;
        end
        10525: begin
            cosine_reg0 <= 36'sb101011111110011100101111010010111101;
            sine_reg0   <= 36'sb100111000010100001100000010001100001;
        end
        10526: begin
            cosine_reg0 <= 36'sb101011111111000011111100111111100000;
            sine_reg0   <= 36'sb100111000010000010000011101100110000;
        end
        10527: begin
            cosine_reg0 <= 36'sb101011111111101011001011011101011100;
            sine_reg0   <= 36'sb100111000001100010101000000101100110;
        end
        10528: begin
            cosine_reg0 <= 36'sb101100000000010010011010101100101111;
            sine_reg0   <= 36'sb100111000001000011001101011100000101;
        end
        10529: begin
            cosine_reg0 <= 36'sb101100000000111001101010101101011000;
            sine_reg0   <= 36'sb100111000000100011110011110000001101;
        end
        10530: begin
            cosine_reg0 <= 36'sb101100000001100000111011011111010101;
            sine_reg0   <= 36'sb100111000000000100011011000001111111;
        end
        10531: begin
            cosine_reg0 <= 36'sb101100000010001000001101000010100100;
            sine_reg0   <= 36'sb100110111111100101000011010001011101;
        end
        10532: begin
            cosine_reg0 <= 36'sb101100000010101111011111010111000100;
            sine_reg0   <= 36'sb100110111111000101101100011110100111;
        end
        10533: begin
            cosine_reg0 <= 36'sb101100000011010110110010011100110100;
            sine_reg0   <= 36'sb100110111110100110010110101001100000;
        end
        10534: begin
            cosine_reg0 <= 36'sb101100000011111110000110010011110010;
            sine_reg0   <= 36'sb100110111110000111000001110010001000;
        end
        10535: begin
            cosine_reg0 <= 36'sb101100000100100101011010111011111100;
            sine_reg0   <= 36'sb100110111101100111101101111000100001;
        end
        10536: begin
            cosine_reg0 <= 36'sb101100000101001100110000010101010001;
            sine_reg0   <= 36'sb100110111101001000011010111100101011;
        end
        10537: begin
            cosine_reg0 <= 36'sb101100000101110100000110011111110000;
            sine_reg0   <= 36'sb100110111100101001001000111110101000;
        end
        10538: begin
            cosine_reg0 <= 36'sb101100000110011011011101011011010110;
            sine_reg0   <= 36'sb100110111100001001110111111110011001;
        end
        10539: begin
            cosine_reg0 <= 36'sb101100000111000010110101001000000011;
            sine_reg0   <= 36'sb100110111011101010100111111100000000;
        end
        10540: begin
            cosine_reg0 <= 36'sb101100000111101010001101100101110101;
            sine_reg0   <= 36'sb100110111011001011011000110111011101;
        end
        10541: begin
            cosine_reg0 <= 36'sb101100001000010001100110110100101010;
            sine_reg0   <= 36'sb100110111010101100001010110000110010;
        end
        10542: begin
            cosine_reg0 <= 36'sb101100001000111001000000110100100010;
            sine_reg0   <= 36'sb100110111010001100111101101000000000;
        end
        10543: begin
            cosine_reg0 <= 36'sb101100001001100000011011100101011001;
            sine_reg0   <= 36'sb100110111001101101110001011101001000;
        end
        10544: begin
            cosine_reg0 <= 36'sb101100001010000111110111000111001111;
            sine_reg0   <= 36'sb100110111001001110100110010000001100;
        end
        10545: begin
            cosine_reg0 <= 36'sb101100001010101111010011011010000011;
            sine_reg0   <= 36'sb100110111000101111011100000001001100;
        end
        10546: begin
            cosine_reg0 <= 36'sb101100001011010110110000011101110010;
            sine_reg0   <= 36'sb100110111000010000010010110000001001;
        end
        10547: begin
            cosine_reg0 <= 36'sb101100001011111110001110010010011100;
            sine_reg0   <= 36'sb100110110111110001001010011101000110;
        end
        10548: begin
            cosine_reg0 <= 36'sb101100001100100101101100110111111110;
            sine_reg0   <= 36'sb100110110111010010000011001000000011;
        end
        10549: begin
            cosine_reg0 <= 36'sb101100001101001101001100001110011000;
            sine_reg0   <= 36'sb100110110110110010111100110001000001;
        end
        10550: begin
            cosine_reg0 <= 36'sb101100001101110100101100010101100111;
            sine_reg0   <= 36'sb100110110110010011110111011000000010;
        end
        10551: begin
            cosine_reg0 <= 36'sb101100001110011100001101001101101010;
            sine_reg0   <= 36'sb100110110101110100110010111101000110;
        end
        10552: begin
            cosine_reg0 <= 36'sb101100001111000011101110110110100000;
            sine_reg0   <= 36'sb100110110101010101101111100000001111;
        end
        10553: begin
            cosine_reg0 <= 36'sb101100001111101011010001010000000111;
            sine_reg0   <= 36'sb100110110100110110101101000001011111;
        end
        10554: begin
            cosine_reg0 <= 36'sb101100010000010010110100011010011110;
            sine_reg0   <= 36'sb100110110100010111101011100000110110;
        end
        10555: begin
            cosine_reg0 <= 36'sb101100010000111010011000010101100011;
            sine_reg0   <= 36'sb100110110011111000101010111110010101;
        end
        10556: begin
            cosine_reg0 <= 36'sb101100010001100001111101000001010100;
            sine_reg0   <= 36'sb100110110011011001101011011001111110;
        end
        10557: begin
            cosine_reg0 <= 36'sb101100010010001001100010011101110001;
            sine_reg0   <= 36'sb100110110010111010101100110011110010;
        end
        10558: begin
            cosine_reg0 <= 36'sb101100010010110001001000101010110110;
            sine_reg0   <= 36'sb100110110010011011101111001011110011;
        end
        10559: begin
            cosine_reg0 <= 36'sb101100010011011000101111101000100100;
            sine_reg0   <= 36'sb100110110001111100110010100010000000;
        end
        10560: begin
            cosine_reg0 <= 36'sb101100010100000000010111010110111001;
            sine_reg0   <= 36'sb100110110001011101110110110110011100;
        end
        10561: begin
            cosine_reg0 <= 36'sb101100010100100111111111110101110010;
            sine_reg0   <= 36'sb100110110000111110111100001001001000;
        end
        10562: begin
            cosine_reg0 <= 36'sb101100010101001111101001000101001110;
            sine_reg0   <= 36'sb100110110000100000000010011010000101;
        end
        10563: begin
            cosine_reg0 <= 36'sb101100010101110111010011000101001101;
            sine_reg0   <= 36'sb100110110000000001001001101001010011;
        end
        10564: begin
            cosine_reg0 <= 36'sb101100010110011110111101110101101011;
            sine_reg0   <= 36'sb100110101111100010010001110110110101;
        end
        10565: begin
            cosine_reg0 <= 36'sb101100010111000110101001010110101001;
            sine_reg0   <= 36'sb100110101111000011011011000010101100;
        end
        10566: begin
            cosine_reg0 <= 36'sb101100010111101110010101101000000100;
            sine_reg0   <= 36'sb100110101110100100100101001100111000;
        end
        10567: begin
            cosine_reg0 <= 36'sb101100011000010110000010101001111010;
            sine_reg0   <= 36'sb100110101110000101110000010101011011;
        end
        10568: begin
            cosine_reg0 <= 36'sb101100011000111101110000011100001011;
            sine_reg0   <= 36'sb100110101101100110111100011100010110;
        end
        10569: begin
            cosine_reg0 <= 36'sb101100011001100101011110111110110100;
            sine_reg0   <= 36'sb100110101101001000001001100001101010;
        end
        10570: begin
            cosine_reg0 <= 36'sb101100011010001101001110010001110101;
            sine_reg0   <= 36'sb100110101100101001010111100101011001;
        end
        10571: begin
            cosine_reg0 <= 36'sb101100011010110100111110010101001011;
            sine_reg0   <= 36'sb100110101100001010100110100111100011;
        end
        10572: begin
            cosine_reg0 <= 36'sb101100011011011100101111001000110101;
            sine_reg0   <= 36'sb100110101011101011110110101000001010;
        end
        10573: begin
            cosine_reg0 <= 36'sb101100011100000100100000101100110010;
            sine_reg0   <= 36'sb100110101011001101000111100111001111;
        end
        10574: begin
            cosine_reg0 <= 36'sb101100011100101100010011000001000000;
            sine_reg0   <= 36'sb100110101010101110011001100100110011;
        end
        10575: begin
            cosine_reg0 <= 36'sb101100011101010100000110000101011101;
            sine_reg0   <= 36'sb100110101010001111101100100000110111;
        end
        10576: begin
            cosine_reg0 <= 36'sb101100011101111011111001111010001001;
            sine_reg0   <= 36'sb100110101001110001000000011011011101;
        end
        10577: begin
            cosine_reg0 <= 36'sb101100011110100011101110011111000000;
            sine_reg0   <= 36'sb100110101001010010010101010100100110;
        end
        10578: begin
            cosine_reg0 <= 36'sb101100011111001011100011110100000011;
            sine_reg0   <= 36'sb100110101000110011101011001100010010;
        end
        10579: begin
            cosine_reg0 <= 36'sb101100011111110011011001111001001111;
            sine_reg0   <= 36'sb100110101000010101000010000010100100;
        end
        10580: begin
            cosine_reg0 <= 36'sb101100100000011011010000101110100010;
            sine_reg0   <= 36'sb100110100111110110011001110111011100;
        end
        10581: begin
            cosine_reg0 <= 36'sb101100100001000011001000010011111100;
            sine_reg0   <= 36'sb100110100111010111110010101010111011;
        end
        10582: begin
            cosine_reg0 <= 36'sb101100100001101011000000101001011011;
            sine_reg0   <= 36'sb100110100110111001001100011101000011;
        end
        10583: begin
            cosine_reg0 <= 36'sb101100100010010010111001101110111101;
            sine_reg0   <= 36'sb100110100110011010100111001101110101;
        end
        10584: begin
            cosine_reg0 <= 36'sb101100100010111010110011100100100000;
            sine_reg0   <= 36'sb100110100101111100000010111101010001;
        end
        10585: begin
            cosine_reg0 <= 36'sb101100100011100010101110001010000100;
            sine_reg0   <= 36'sb100110100101011101011111101011011010;
        end
        10586: begin
            cosine_reg0 <= 36'sb101100100100001010101001011111100110;
            sine_reg0   <= 36'sb100110100100111110111101011000010000;
        end
        10587: begin
            cosine_reg0 <= 36'sb101100100100110010100101100101000101;
            sine_reg0   <= 36'sb100110100100100000011100000011110101;
        end
        10588: begin
            cosine_reg0 <= 36'sb101100100101011010100010011010100000;
            sine_reg0   <= 36'sb100110100100000001111011101110001001;
        end
        10589: begin
            cosine_reg0 <= 36'sb101100100110000010011111111111110101;
            sine_reg0   <= 36'sb100110100011100011011100010111001110;
        end
        10590: begin
            cosine_reg0 <= 36'sb101100100110101010011110010101000010;
            sine_reg0   <= 36'sb100110100011000100111101111111000110;
        end
        10591: begin
            cosine_reg0 <= 36'sb101100100111010010011101011010000110;
            sine_reg0   <= 36'sb100110100010100110100000100101110000;
        end
        10592: begin
            cosine_reg0 <= 36'sb101100100111111010011101001110111111;
            sine_reg0   <= 36'sb100110100010001000000100001011001111;
        end
        10593: begin
            cosine_reg0 <= 36'sb101100101000100010011101110011101100;
            sine_reg0   <= 36'sb100110100001101001101000101111100011;
        end
        10594: begin
            cosine_reg0 <= 36'sb101100101001001010011111001000001011;
            sine_reg0   <= 36'sb100110100001001011001110010010101110;
        end
        10595: begin
            cosine_reg0 <= 36'sb101100101001110010100001001100011011;
            sine_reg0   <= 36'sb100110100000101100110100110100110001;
        end
        10596: begin
            cosine_reg0 <= 36'sb101100101010011010100100000000011011;
            sine_reg0   <= 36'sb100110100000001110011100010101101101;
        end
        10597: begin
            cosine_reg0 <= 36'sb101100101011000010100111100100001000;
            sine_reg0   <= 36'sb100110011111110000000100110101100011;
        end
        10598: begin
            cosine_reg0 <= 36'sb101100101011101010101011110111100000;
            sine_reg0   <= 36'sb100110011111010001101110010100010101;
        end
        10599: begin
            cosine_reg0 <= 36'sb101100101100010010110000111010100100;
            sine_reg0   <= 36'sb100110011110110011011000110010000011;
        end
        10600: begin
            cosine_reg0 <= 36'sb101100101100111010110110101101010000;
            sine_reg0   <= 36'sb100110011110010101000100001110101111;
        end
        10601: begin
            cosine_reg0 <= 36'sb101100101101100010111101001111100100;
            sine_reg0   <= 36'sb100110011101110110110000101010011010;
        end
        10602: begin
            cosine_reg0 <= 36'sb101100101110001011000100100001011110;
            sine_reg0   <= 36'sb100110011101011000011110000101000101;
        end
        10603: begin
            cosine_reg0 <= 36'sb101100101110110011001100100010111100;
            sine_reg0   <= 36'sb100110011100111010001100011110110010;
        end
        10604: begin
            cosine_reg0 <= 36'sb101100101111011011010101010011111101;
            sine_reg0   <= 36'sb100110011100011011111011110111100000;
        end
        10605: begin
            cosine_reg0 <= 36'sb101100110000000011011110110100011111;
            sine_reg0   <= 36'sb100110011011111101101100001111010011;
        end
        10606: begin
            cosine_reg0 <= 36'sb101100110000101011101001000100100001;
            sine_reg0   <= 36'sb100110011011011111011101100110001010;
        end
        10607: begin
            cosine_reg0 <= 36'sb101100110001010011110100000100000001;
            sine_reg0   <= 36'sb100110011011000001001111111100000111;
        end
        10608: begin
            cosine_reg0 <= 36'sb101100110001111011111111110010111101;
            sine_reg0   <= 36'sb100110011010100011000011010001001011;
        end
        10609: begin
            cosine_reg0 <= 36'sb101100110010100100001100010001010101;
            sine_reg0   <= 36'sb100110011010000100110111100101010111;
        end
        10610: begin
            cosine_reg0 <= 36'sb101100110011001100011001011111000110;
            sine_reg0   <= 36'sb100110011001100110101100111000101101;
        end
        10611: begin
            cosine_reg0 <= 36'sb101100110011110100100111011100001111;
            sine_reg0   <= 36'sb100110011001001000100011001011001101;
        end
        10612: begin
            cosine_reg0 <= 36'sb101100110100011100110110001000101111;
            sine_reg0   <= 36'sb100110011000101010011010011100111001;
        end
        10613: begin
            cosine_reg0 <= 36'sb101100110101000101000101100100100011;
            sine_reg0   <= 36'sb100110011000001100010010101101110010;
        end
        10614: begin
            cosine_reg0 <= 36'sb101100110101101101010101101111101011;
            sine_reg0   <= 36'sb100110010111101110001011111101111001;
        end
        10615: begin
            cosine_reg0 <= 36'sb101100110110010101100110101010000101;
            sine_reg0   <= 36'sb100110010111010000000110001101001111;
        end
        10616: begin
            cosine_reg0 <= 36'sb101100110110111101111000010011101110;
            sine_reg0   <= 36'sb100110010110110010000001011011110110;
        end
        10617: begin
            cosine_reg0 <= 36'sb101100110111100110001010101100100110;
            sine_reg0   <= 36'sb100110010110010011111101101001101110;
        end
        10618: begin
            cosine_reg0 <= 36'sb101100111000001110011101110100101100;
            sine_reg0   <= 36'sb100110010101110101111010110110111001;
        end
        10619: begin
            cosine_reg0 <= 36'sb101100111000110110110001101011111101;
            sine_reg0   <= 36'sb100110010101010111111001000011011000;
        end
        10620: begin
            cosine_reg0 <= 36'sb101100111001011111000110010010011000;
            sine_reg0   <= 36'sb100110010100111001111000001111001100;
        end
        10621: begin
            cosine_reg0 <= 36'sb101100111010000111011011100111111011;
            sine_reg0   <= 36'sb100110010100011011111000011010010110;
        end
        10622: begin
            cosine_reg0 <= 36'sb101100111010101111110001101100100101;
            sine_reg0   <= 36'sb100110010011111101111001100100110111;
        end
        10623: begin
            cosine_reg0 <= 36'sb101100111011011000001000100000010101;
            sine_reg0   <= 36'sb100110010011011111111011101110110001;
        end
        10624: begin
            cosine_reg0 <= 36'sb101100111100000000100000000011001000;
            sine_reg0   <= 36'sb100110010011000001111110111000000100;
        end
        10625: begin
            cosine_reg0 <= 36'sb101100111100101000111000010100111110;
            sine_reg0   <= 36'sb100110010010100100000011000000110010;
        end
        10626: begin
            cosine_reg0 <= 36'sb101100111101010001010001010101110100;
            sine_reg0   <= 36'sb100110010010000110001000001000111100;
        end
        10627: begin
            cosine_reg0 <= 36'sb101100111101111001101011000101101001;
            sine_reg0   <= 36'sb100110010001101000001110010000100100;
        end
        10628: begin
            cosine_reg0 <= 36'sb101100111110100010000101100100011100;
            sine_reg0   <= 36'sb100110010001001010010101010111101001;
        end
        10629: begin
            cosine_reg0 <= 36'sb101100111111001010100000110010001011;
            sine_reg0   <= 36'sb100110010000101100011101011110001110;
        end
        10630: begin
            cosine_reg0 <= 36'sb101100111111110010111100101110110100;
            sine_reg0   <= 36'sb100110010000001110100110100100010011;
        end
        10631: begin
            cosine_reg0 <= 36'sb101101000000011011011001011010010110;
            sine_reg0   <= 36'sb100110001111110000110000101001111011;
        end
        10632: begin
            cosine_reg0 <= 36'sb101101000001000011110110110100110000;
            sine_reg0   <= 36'sb100110001111010010111011101111000101;
        end
        10633: begin
            cosine_reg0 <= 36'sb101101000001101100010100111101111111;
            sine_reg0   <= 36'sb100110001110110101000111110011110011;
        end
        10634: begin
            cosine_reg0 <= 36'sb101101000010010100110011110110000010;
            sine_reg0   <= 36'sb100110001110010111010100111000000110;
        end
        10635: begin
            cosine_reg0 <= 36'sb101101000010111101010011011100111000;
            sine_reg0   <= 36'sb100110001101111001100010111100000000;
        end
        10636: begin
            cosine_reg0 <= 36'sb101101000011100101110011110010011111;
            sine_reg0   <= 36'sb100110001101011011110001111111100001;
        end
        10637: begin
            cosine_reg0 <= 36'sb101101000100001110010100110110110101;
            sine_reg0   <= 36'sb100110001100111110000010000010101010;
        end
        10638: begin
            cosine_reg0 <= 36'sb101101000100110110110110101001111010;
            sine_reg0   <= 36'sb100110001100100000010011000101011110;
        end
        10639: begin
            cosine_reg0 <= 36'sb101101000101011111011001001011101011;
            sine_reg0   <= 36'sb100110001100000010100101000111111100;
        end
        10640: begin
            cosine_reg0 <= 36'sb101101000110000111111100011100000110;
            sine_reg0   <= 36'sb100110001011100100111000001010000110;
        end
        10641: begin
            cosine_reg0 <= 36'sb101101000110110000100000011011001011;
            sine_reg0   <= 36'sb100110001011000111001100001011111110;
        end
        10642: begin
            cosine_reg0 <= 36'sb101101000111011001000101001000111000;
            sine_reg0   <= 36'sb100110001010101001100001001101100100;
        end
        10643: begin
            cosine_reg0 <= 36'sb101101001000000001101010100101001010;
            sine_reg0   <= 36'sb100110001010001011110111001110111001;
        end
        10644: begin
            cosine_reg0 <= 36'sb101101001000101010010000110000000010;
            sine_reg0   <= 36'sb100110001001101110001110001111111111;
        end
        10645: begin
            cosine_reg0 <= 36'sb101101001001010010110111101001011100;
            sine_reg0   <= 36'sb100110001001010000100110010000110111;
        end
        10646: begin
            cosine_reg0 <= 36'sb101101001001111011011111010001011000;
            sine_reg0   <= 36'sb100110001000110010111111010001100001;
        end
        10647: begin
            cosine_reg0 <= 36'sb101101001010100100000111100111110011;
            sine_reg0   <= 36'sb100110001000010101011001010010000000;
        end
        10648: begin
            cosine_reg0 <= 36'sb101101001011001100110000101100101101;
            sine_reg0   <= 36'sb100110000111110111110100010010010100;
        end
        10649: begin
            cosine_reg0 <= 36'sb101101001011110101011010100000000011;
            sine_reg0   <= 36'sb100110000111011010010000010010011110;
        end
        10650: begin
            cosine_reg0 <= 36'sb101101001100011110000101000001110101;
            sine_reg0   <= 36'sb100110000110111100101101010010100000;
        end
        10651: begin
            cosine_reg0 <= 36'sb101101001101000110110000010010000000;
            sine_reg0   <= 36'sb100110000110011111001011010010011010;
        end
        10652: begin
            cosine_reg0 <= 36'sb101101001101101111011100010000100100;
            sine_reg0   <= 36'sb100110000110000001101010010010001110;
        end
        10653: begin
            cosine_reg0 <= 36'sb101101001110011000001000111101011110;
            sine_reg0   <= 36'sb100110000101100100001010010001111101;
        end
        10654: begin
            cosine_reg0 <= 36'sb101101001111000000110110011000101100;
            sine_reg0   <= 36'sb100110000101000110101011010001101000;
        end
        10655: begin
            cosine_reg0 <= 36'sb101101001111101001100100100010001110;
            sine_reg0   <= 36'sb100110000100101001001101010001010000;
        end
        10656: begin
            cosine_reg0 <= 36'sb101101010000010010010011011010000010;
            sine_reg0   <= 36'sb100110000100001011110000010000110110;
        end
        10657: begin
            cosine_reg0 <= 36'sb101101010000111011000011000000000110;
            sine_reg0   <= 36'sb100110000011101110010100010000011100;
        end
        10658: begin
            cosine_reg0 <= 36'sb101101010001100011110011010100011000;
            sine_reg0   <= 36'sb100110000011010000111001010000000011;
        end
        10659: begin
            cosine_reg0 <= 36'sb101101010010001100100100010110111000;
            sine_reg0   <= 36'sb100110000010110011011111001111101011;
        end
        10660: begin
            cosine_reg0 <= 36'sb101101010010110101010110000111100011;
            sine_reg0   <= 36'sb100110000010010110000110001111010110;
        end
        10661: begin
            cosine_reg0 <= 36'sb101101010011011110001000100110011000;
            sine_reg0   <= 36'sb100110000001111000101110001111000101;
        end
        10662: begin
            cosine_reg0 <= 36'sb101101010100000110111011110011010101;
            sine_reg0   <= 36'sb100110000001011011010111001110111001;
        end
        10663: begin
            cosine_reg0 <= 36'sb101101010100101111101111101110011001;
            sine_reg0   <= 36'sb100110000000111110000001001110110011;
        end
        10664: begin
            cosine_reg0 <= 36'sb101101010101011000100100010111100010;
            sine_reg0   <= 36'sb100110000000100000101100001110110100;
        end
        10665: begin
            cosine_reg0 <= 36'sb101101010110000001011001101110101111;
            sine_reg0   <= 36'sb100110000000000011011000001110111111;
        end
        10666: begin
            cosine_reg0 <= 36'sb101101010110101010001111110011111101;
            sine_reg0   <= 36'sb100101111111100110000101001111010010;
        end
        10667: begin
            cosine_reg0 <= 36'sb101101010111010011000110100111001100;
            sine_reg0   <= 36'sb100101111111001000110011001111110001;
        end
        10668: begin
            cosine_reg0 <= 36'sb101101010111111011111110001000011011;
            sine_reg0   <= 36'sb100101111110101011100010010000011011;
        end
        10669: begin
            cosine_reg0 <= 36'sb101101011000100100110110010111100110;
            sine_reg0   <= 36'sb100101111110001110010010010001010011;
        end
        10670: begin
            cosine_reg0 <= 36'sb101101011001001101101111010100101101;
            sine_reg0   <= 36'sb100101111101110001000011010010011000;
        end
        10671: begin
            cosine_reg0 <= 36'sb101101011001110110101000111111101110;
            sine_reg0   <= 36'sb100101111101010011110101010011101101;
        end
        10672: begin
            cosine_reg0 <= 36'sb101101011010011111100011011000101000;
            sine_reg0   <= 36'sb100101111100110110101000010101010010;
        end
        10673: begin
            cosine_reg0 <= 36'sb101101011011001000011110011111011001;
            sine_reg0   <= 36'sb100101111100011001011100010111001001;
        end
        10674: begin
            cosine_reg0 <= 36'sb101101011011110001011010010011111111;
            sine_reg0   <= 36'sb100101111011111100010001011001010010;
        end
        10675: begin
            cosine_reg0 <= 36'sb101101011100011010010110110110011001;
            sine_reg0   <= 36'sb100101111011011111000111011011101111;
        end
        10676: begin
            cosine_reg0 <= 36'sb101101011101000011010100000110100101;
            sine_reg0   <= 36'sb100101111011000001111110011110100001;
        end
        10677: begin
            cosine_reg0 <= 36'sb101101011101101100010010000100100010;
            sine_reg0   <= 36'sb100101111010100100110110100001101001;
        end
        10678: begin
            cosine_reg0 <= 36'sb101101011110010101010000110000001110;
            sine_reg0   <= 36'sb100101111010000111101111100101001000;
        end
        10679: begin
            cosine_reg0 <= 36'sb101101011110111110010000001001101000;
            sine_reg0   <= 36'sb100101111001101010101001101001000000;
        end
        10680: begin
            cosine_reg0 <= 36'sb101101011111100111010000010000101101;
            sine_reg0   <= 36'sb100101111001001101100100101101010001;
        end
        10681: begin
            cosine_reg0 <= 36'sb101101100000010000010001000101011101;
            sine_reg0   <= 36'sb100101111000110000100000110001111100;
        end
        10682: begin
            cosine_reg0 <= 36'sb101101100000111001010010100111110110;
            sine_reg0   <= 36'sb100101111000010011011101110111000011;
        end
        10683: begin
            cosine_reg0 <= 36'sb101101100001100010010100110111110110;
            sine_reg0   <= 36'sb100101110111110110011011111100100111;
        end
        10684: begin
            cosine_reg0 <= 36'sb101101100010001011010111110101011011;
            sine_reg0   <= 36'sb100101110111011001011011000010101000;
        end
        10685: begin
            cosine_reg0 <= 36'sb101101100010110100011011100000100101;
            sine_reg0   <= 36'sb100101110110111100011011001001001001;
        end
        10686: begin
            cosine_reg0 <= 36'sb101101100011011101011111111001010000;
            sine_reg0   <= 36'sb100101110110011111011100010000001001;
        end
        10687: begin
            cosine_reg0 <= 36'sb101101100100000110100100111111011101;
            sine_reg0   <= 36'sb100101110110000010011110010111101011;
        end
        10688: begin
            cosine_reg0 <= 36'sb101101100100101111101010110011001001;
            sine_reg0   <= 36'sb100101110101100101100001011111101111;
        end
        10689: begin
            cosine_reg0 <= 36'sb101101100101011000110001010100010011;
            sine_reg0   <= 36'sb100101110101001000100101101000010111;
        end
        10690: begin
            cosine_reg0 <= 36'sb101101100110000001111000100010111001;
            sine_reg0   <= 36'sb100101110100101011101010110001100011;
        end
        10691: begin
            cosine_reg0 <= 36'sb101101100110101011000000011110111001;
            sine_reg0   <= 36'sb100101110100001110110000111011010101;
        end
        10692: begin
            cosine_reg0 <= 36'sb101101100111010100001001001000010011;
            sine_reg0   <= 36'sb100101110011110001111000000101101110;
        end
        10693: begin
            cosine_reg0 <= 36'sb101101100111111101010010011111000011;
            sine_reg0   <= 36'sb100101110011010101000000010000101110;
        end
        10694: begin
            cosine_reg0 <= 36'sb101101101000100110011100100011001010;
            sine_reg0   <= 36'sb100101110010111000001001011100011000;
        end
        10695: begin
            cosine_reg0 <= 36'sb101101101001001111100111010100100100;
            sine_reg0   <= 36'sb100101110010011011010011101000101100;
        end
        10696: begin
            cosine_reg0 <= 36'sb101101101001111000110010110011010010;
            sine_reg0   <= 36'sb100101110001111110011110110101101011;
        end
        10697: begin
            cosine_reg0 <= 36'sb101101101010100001111110111111010000;
            sine_reg0   <= 36'sb100101110001100001101011000011010110;
        end
        10698: begin
            cosine_reg0 <= 36'sb101101101011001011001011111000011110;
            sine_reg0   <= 36'sb100101110001000100111000010001101111;
        end
        10699: begin
            cosine_reg0 <= 36'sb101101101011110100011001011110111001;
            sine_reg0   <= 36'sb100101110000101000000110100000110110;
        end
        10700: begin
            cosine_reg0 <= 36'sb101101101100011101100111110010100001;
            sine_reg0   <= 36'sb100101110000001011010101110000101101;
        end
        10701: begin
            cosine_reg0 <= 36'sb101101101101000110110110110011010011;
            sine_reg0   <= 36'sb100101101111101110100110000001010101;
        end
        10702: begin
            cosine_reg0 <= 36'sb101101101101110000000110100001001111;
            sine_reg0   <= 36'sb100101101111010001110111010010101111;
        end
        10703: begin
            cosine_reg0 <= 36'sb101101101110011001010110111100010010;
            sine_reg0   <= 36'sb100101101110110101001001100100111100;
        end
        10704: begin
            cosine_reg0 <= 36'sb101101101111000010101000000100011010;
            sine_reg0   <= 36'sb100101101110011000011100110111111100;
        end
        10705: begin
            cosine_reg0 <= 36'sb101101101111101011111001111001100111;
            sine_reg0   <= 36'sb100101101101111011110001001011110011;
        end
        10706: begin
            cosine_reg0 <= 36'sb101101110000010101001100011011110111;
            sine_reg0   <= 36'sb100101101101011111000110100000011111;
        end
        10707: begin
            cosine_reg0 <= 36'sb101101110000111110011111101011001000;
            sine_reg0   <= 36'sb100101101101000010011100110110000011;
        end
        10708: begin
            cosine_reg0 <= 36'sb101101110001100111110011100111011001;
            sine_reg0   <= 36'sb100101101100100101110100001100011111;
        end
        10709: begin
            cosine_reg0 <= 36'sb101101110010010001001000010000100111;
            sine_reg0   <= 36'sb100101101100001001001100100011110101;
        end
        10710: begin
            cosine_reg0 <= 36'sb101101110010111010011101100110110010;
            sine_reg0   <= 36'sb100101101011101100100101111100000110;
        end
        10711: begin
            cosine_reg0 <= 36'sb101101110011100011110011101001110111;
            sine_reg0   <= 36'sb100101101011010000000000010101010011;
        end
        10712: begin
            cosine_reg0 <= 36'sb101101110100001101001010011001110110;
            sine_reg0   <= 36'sb100101101010110011011011101111011101;
        end
        10713: begin
            cosine_reg0 <= 36'sb101101110100110110100001110110101100;
            sine_reg0   <= 36'sb100101101010010110111000001010100100;
        end
        10714: begin
            cosine_reg0 <= 36'sb101101110101011111111010000000011000;
            sine_reg0   <= 36'sb100101101001111010010101100110101011;
        end
        10715: begin
            cosine_reg0 <= 36'sb101101110110001001010010110110111000;
            sine_reg0   <= 36'sb100101101001011101110100000011110010;
        end
        10716: begin
            cosine_reg0 <= 36'sb101101110110110010101100011010001011;
            sine_reg0   <= 36'sb100101101001000001010011100001111011;
        end
        10717: begin
            cosine_reg0 <= 36'sb101101110111011100000110101010010000;
            sine_reg0   <= 36'sb100101101000100100110100000001000110;
        end
        10718: begin
            cosine_reg0 <= 36'sb101101111000000101100001100111000011;
            sine_reg0   <= 36'sb100101101000001000010101100001010100;
        end
        10719: begin
            cosine_reg0 <= 36'sb101101111000101110111101010000100101;
            sine_reg0   <= 36'sb100101100111101011111000000010100111;
        end
        10720: begin
            cosine_reg0 <= 36'sb101101111001011000011001100110110100;
            sine_reg0   <= 36'sb100101100111001111011011100101000000;
        end
        10721: begin
            cosine_reg0 <= 36'sb101101111010000001110110101001101101;
            sine_reg0   <= 36'sb100101100110110011000000001000100000;
        end
        10722: begin
            cosine_reg0 <= 36'sb101101111010101011010100011001001111;
            sine_reg0   <= 36'sb100101100110010110100101101101000111;
        end
        10723: begin
            cosine_reg0 <= 36'sb101101111011010100110010110101011001;
            sine_reg0   <= 36'sb100101100101111010001100010010111000;
        end
        10724: begin
            cosine_reg0 <= 36'sb101101111011111110010001111110001000;
            sine_reg0   <= 36'sb100101100101011101110011111001110011;
        end
        10725: begin
            cosine_reg0 <= 36'sb101101111100100111110001110011011100;
            sine_reg0   <= 36'sb100101100101000001011100100001111001;
        end
        10726: begin
            cosine_reg0 <= 36'sb101101111101010001010010010101010011;
            sine_reg0   <= 36'sb100101100100100101000110001011001011;
        end
        10727: begin
            cosine_reg0 <= 36'sb101101111101111010110011100011101100;
            sine_reg0   <= 36'sb100101100100001000110000110101101011;
        end
        10728: begin
            cosine_reg0 <= 36'sb101101111110100100010101011110100011;
            sine_reg0   <= 36'sb100101100011101100011100100001011001;
        end
        10729: begin
            cosine_reg0 <= 36'sb101101111111001101111000000101111001;
            sine_reg0   <= 36'sb100101100011010000001001001110010111;
        end
        10730: begin
            cosine_reg0 <= 36'sb101101111111110111011011011001101011;
            sine_reg0   <= 36'sb100101100010110011110110111100100110;
        end
        10731: begin
            cosine_reg0 <= 36'sb101110000000100000111111011001111000;
            sine_reg0   <= 36'sb100101100010010111100101101100000110;
        end
        10732: begin
            cosine_reg0 <= 36'sb101110000001001010100100000110011110;
            sine_reg0   <= 36'sb100101100001111011010101011100111010;
        end
        10733: begin
            cosine_reg0 <= 36'sb101110000001110100001001011111011011;
            sine_reg0   <= 36'sb100101100001011111000110001111000001;
        end
        10734: begin
            cosine_reg0 <= 36'sb101110000010011101101111100100101111;
            sine_reg0   <= 36'sb100101100001000010111000000010011101;
        end
        10735: begin
            cosine_reg0 <= 36'sb101110000011000111010110010110010111;
            sine_reg0   <= 36'sb100101100000100110101010110111001111;
        end
        10736: begin
            cosine_reg0 <= 36'sb101110000011110000111101110100010001;
            sine_reg0   <= 36'sb100101100000001010011110101101011001;
        end
        10737: begin
            cosine_reg0 <= 36'sb101110000100011010100101111110011101;
            sine_reg0   <= 36'sb100101011111101110010011100100111011;
        end
        10738: begin
            cosine_reg0 <= 36'sb101110000101000100001110110100111001;
            sine_reg0   <= 36'sb100101011111010010001001011101110110;
        end
        10739: begin
            cosine_reg0 <= 36'sb101110000101101101111000010111100010;
            sine_reg0   <= 36'sb100101011110110110000000011000001100;
        end
        10740: begin
            cosine_reg0 <= 36'sb101110000110010111100010100110011000;
            sine_reg0   <= 36'sb100101011110011001111000010011111101;
        end
        10741: begin
            cosine_reg0 <= 36'sb101110000111000001001101100001011000;
            sine_reg0   <= 36'sb100101011101111101110001010001001011;
        end
        10742: begin
            cosine_reg0 <= 36'sb101110000111101010111001001000100001;
            sine_reg0   <= 36'sb100101011101100001101011001111110111;
        end
        10743: begin
            cosine_reg0 <= 36'sb101110001000010100100101011011110011;
            sine_reg0   <= 36'sb100101011101000101100110010000000001;
        end
        10744: begin
            cosine_reg0 <= 36'sb101110001000111110010010011011001001;
            sine_reg0   <= 36'sb100101011100101001100010010001101100;
        end
        10745: begin
            cosine_reg0 <= 36'sb101110001001101000000000000110100101;
            sine_reg0   <= 36'sb100101011100001101011111010100110111;
        end
        10746: begin
            cosine_reg0 <= 36'sb101110001010010001101110011110000011;
            sine_reg0   <= 36'sb100101011011110001011101011001100101;
        end
        10747: begin
            cosine_reg0 <= 36'sb101110001010111011011101100001100010;
            sine_reg0   <= 36'sb100101011011010101011100011111110101;
        end
        10748: begin
            cosine_reg0 <= 36'sb101110001011100101001101010001000000;
            sine_reg0   <= 36'sb100101011010111001011100100111101010;
        end
        10749: begin
            cosine_reg0 <= 36'sb101110001100001110111101101100011101;
            sine_reg0   <= 36'sb100101011010011101011101110001000100;
        end
        10750: begin
            cosine_reg0 <= 36'sb101110001100111000101110110011110101;
            sine_reg0   <= 36'sb100101011010000001011111111100000101;
        end
        10751: begin
            cosine_reg0 <= 36'sb101110001101100010100000100111001001;
            sine_reg0   <= 36'sb100101011001100101100011001000101101;
        end
        10752: begin
            cosine_reg0 <= 36'sb101110001110001100010011000110010101;
            sine_reg0   <= 36'sb100101011001001001100111010110111101;
        end
        10753: begin
            cosine_reg0 <= 36'sb101110001110110110000110010001011001;
            sine_reg0   <= 36'sb100101011000101101101100100110110111;
        end
        10754: begin
            cosine_reg0 <= 36'sb101110001111011111111010001000010010;
            sine_reg0   <= 36'sb100101011000010001110010111000011100;
        end
        10755: begin
            cosine_reg0 <= 36'sb101110010000001001101110101011000000;
            sine_reg0   <= 36'sb100101010111110101111010001011101101;
        end
        10756: begin
            cosine_reg0 <= 36'sb101110010000110011100011111001100000;
            sine_reg0   <= 36'sb100101010111011010000010100000101010;
        end
        10757: begin
            cosine_reg0 <= 36'sb101110010001011101011001110011110010;
            sine_reg0   <= 36'sb100101010110111110001011110111010101;
        end
        10758: begin
            cosine_reg0 <= 36'sb101110010010000111010000011001110011;
            sine_reg0   <= 36'sb100101010110100010010110001111110000;
        end
        10759: begin
            cosine_reg0 <= 36'sb101110010010110001000111101011100001;
            sine_reg0   <= 36'sb100101010110000110100001101001111010;
        end
        10760: begin
            cosine_reg0 <= 36'sb101110010011011010111111101000111100;
            sine_reg0   <= 36'sb100101010101101010101110000101110110;
        end
        10761: begin
            cosine_reg0 <= 36'sb101110010100000100111000010010000001;
            sine_reg0   <= 36'sb100101010101001110111011100011100011;
        end
        10762: begin
            cosine_reg0 <= 36'sb101110010100101110110001100110101111;
            sine_reg0   <= 36'sb100101010100110011001010000011000100;
        end
        10763: begin
            cosine_reg0 <= 36'sb101110010101011000101011100111000100;
            sine_reg0   <= 36'sb100101010100010111011001100100011010;
        end
        10764: begin
            cosine_reg0 <= 36'sb101110010110000010100110010010111111;
            sine_reg0   <= 36'sb100101010011111011101010000111100100;
        end
        10765: begin
            cosine_reg0 <= 36'sb101110010110101100100001101010011110;
            sine_reg0   <= 36'sb100101010011011111111011101100100110;
        end
        10766: begin
            cosine_reg0 <= 36'sb101110010111010110011101101101100000;
            sine_reg0   <= 36'sb100101010011000100001110010011011111;
        end
        10767: begin
            cosine_reg0 <= 36'sb101110011000000000011010011100000010;
            sine_reg0   <= 36'sb100101010010101000100001111100010000;
        end
        10768: begin
            cosine_reg0 <= 36'sb101110011000101010010111110110000100;
            sine_reg0   <= 36'sb100101010010001100110110100110111011;
        end
        10769: begin
            cosine_reg0 <= 36'sb101110011001010100010101111011100011;
            sine_reg0   <= 36'sb100101010001110001001100010011100001;
        end
        10770: begin
            cosine_reg0 <= 36'sb101110011001111110010100101100011110;
            sine_reg0   <= 36'sb100101010001010101100011000010000011;
        end
        10771: begin
            cosine_reg0 <= 36'sb101110011010101000010100001000110100;
            sine_reg0   <= 36'sb100101010000111001111010110010100001;
        end
        10772: begin
            cosine_reg0 <= 36'sb101110011011010010010100010000100010;
            sine_reg0   <= 36'sb100101010000011110010011100100111110;
        end
        10773: begin
            cosine_reg0 <= 36'sb101110011011111100010101000011100111;
            sine_reg0   <= 36'sb100101010000000010101101011001011010;
        end
        10774: begin
            cosine_reg0 <= 36'sb101110011100100110010110100010000010;
            sine_reg0   <= 36'sb100101001111100111001000001111110101;
        end
        10775: begin
            cosine_reg0 <= 36'sb101110011101010000011000101011110001;
            sine_reg0   <= 36'sb100101001111001011100100001000010010;
        end
        10776: begin
            cosine_reg0 <= 36'sb101110011101111010011011100000110010;
            sine_reg0   <= 36'sb100101001110110000000001000010110001;
        end
        10777: begin
            cosine_reg0 <= 36'sb101110011110100100011111000001000100;
            sine_reg0   <= 36'sb100101001110010100011110111111010011;
        end
        10778: begin
            cosine_reg0 <= 36'sb101110011111001110100011001100100100;
            sine_reg0   <= 36'sb100101001101111000111101111101111010;
        end
        10779: begin
            cosine_reg0 <= 36'sb101110011111111000101000000011010010;
            sine_reg0   <= 36'sb100101001101011101011101111110100110;
        end
        10780: begin
            cosine_reg0 <= 36'sb101110100000100010101101100101001100;
            sine_reg0   <= 36'sb100101001101000001111111000001011001;
        end
        10781: begin
            cosine_reg0 <= 36'sb101110100001001100110011110010010000;
            sine_reg0   <= 36'sb100101001100100110100001000110010011;
        end
        10782: begin
            cosine_reg0 <= 36'sb101110100001110110111010101010011101;
            sine_reg0   <= 36'sb100101001100001011000100001101010101;
        end
        10783: begin
            cosine_reg0 <= 36'sb101110100010100001000010001101110000;
            sine_reg0   <= 36'sb100101001011101111101000010110100001;
        end
        10784: begin
            cosine_reg0 <= 36'sb101110100011001011001010011100001001;
            sine_reg0   <= 36'sb100101001011010100001101100001111000;
        end
        10785: begin
            cosine_reg0 <= 36'sb101110100011110101010011010101100101;
            sine_reg0   <= 36'sb100101001010111000110011101111011011;
        end
        10786: begin
            cosine_reg0 <= 36'sb101110100100011111011100111010000100;
            sine_reg0   <= 36'sb100101001010011101011010111111001011;
        end
        10787: begin
            cosine_reg0 <= 36'sb101110100101001001100111001001100010;
            sine_reg0   <= 36'sb100101001010000010000011010001001000;
        end
        10788: begin
            cosine_reg0 <= 36'sb101110100101110011110010000100000000;
            sine_reg0   <= 36'sb100101001001100110101100100101010100;
        end
        10789: begin
            cosine_reg0 <= 36'sb101110100110011101111101101001011011;
            sine_reg0   <= 36'sb100101001001001011010110111011110000;
        end
        10790: begin
            cosine_reg0 <= 36'sb101110100111001000001001111001110001;
            sine_reg0   <= 36'sb100101001000110000000010010100011110;
        end
        10791: begin
            cosine_reg0 <= 36'sb101110100111110010010110110101000001;
            sine_reg0   <= 36'sb100101001000010100101110101111011101;
        end
        10792: begin
            cosine_reg0 <= 36'sb101110101000011100100100011011001010;
            sine_reg0   <= 36'sb100101000111111001011100001100101111;
        end
        10793: begin
            cosine_reg0 <= 36'sb101110101001000110110010101100001001;
            sine_reg0   <= 36'sb100101000111011110001010101100010110;
        end
        10794: begin
            cosine_reg0 <= 36'sb101110101001110001000001100111111101;
            sine_reg0   <= 36'sb100101000111000010111010001110010010;
        end
        10795: begin
            cosine_reg0 <= 36'sb101110101010011011010001001110100100;
            sine_reg0   <= 36'sb100101000110100111101010110010100100;
        end
        10796: begin
            cosine_reg0 <= 36'sb101110101011000101100001011111111110;
            sine_reg0   <= 36'sb100101000110001100011100011001001110;
        end
        10797: begin
            cosine_reg0 <= 36'sb101110101011101111110010011100000111;
            sine_reg0   <= 36'sb100101000101110001001111000010001111;
        end
        10798: begin
            cosine_reg0 <= 36'sb101110101100011010000100000010111111;
            sine_reg0   <= 36'sb100101000101010110000010101101101011;
        end
        10799: begin
            cosine_reg0 <= 36'sb101110101101000100010110010100100100;
            sine_reg0   <= 36'sb100101000100111010110111011011100000;
        end
        10800: begin
            cosine_reg0 <= 36'sb101110101101101110101001010000110100;
            sine_reg0   <= 36'sb100101000100011111101101001011110010;
        end
        10801: begin
            cosine_reg0 <= 36'sb101110101110011000111100110111101101;
            sine_reg0   <= 36'sb100101000100000100100011111110100000;
        end
        10802: begin
            cosine_reg0 <= 36'sb101110101111000011010001001001001111;
            sine_reg0   <= 36'sb100101000011101001011011110011101011;
        end
        10803: begin
            cosine_reg0 <= 36'sb101110101111101101100110000101010111;
            sine_reg0   <= 36'sb100101000011001110010100101011010101;
        end
        10804: begin
            cosine_reg0 <= 36'sb101110110000010111111011101100000100;
            sine_reg0   <= 36'sb100101000010110011001110100101011111;
        end
        10805: begin
            cosine_reg0 <= 36'sb101110110001000010010001111101010011;
            sine_reg0   <= 36'sb100101000010011000001001100010001010;
        end
        10806: begin
            cosine_reg0 <= 36'sb101110110001101100101000111001000101;
            sine_reg0   <= 36'sb100101000001111101000101100001010110;
        end
        10807: begin
            cosine_reg0 <= 36'sb101110110010010111000000011111010110;
            sine_reg0   <= 36'sb100101000001100010000010100011000110;
        end
        10808: begin
            cosine_reg0 <= 36'sb101110110011000001011000110000000101;
            sine_reg0   <= 36'sb100101000001000111000000100111011001;
        end
        10809: begin
            cosine_reg0 <= 36'sb101110110011101011110001101011010001;
            sine_reg0   <= 36'sb100101000000101011111111101110010001;
        end
        10810: begin
            cosine_reg0 <= 36'sb101110110100010110001011010000111000;
            sine_reg0   <= 36'sb100101000000010000111111110111101111;
        end
        10811: begin
            cosine_reg0 <= 36'sb101110110101000000100101100000111000;
            sine_reg0   <= 36'sb100100111111110110000001000011110100;
        end
        10812: begin
            cosine_reg0 <= 36'sb101110110101101011000000011011001111;
            sine_reg0   <= 36'sb100100111111011011000011010010100010;
        end
        10813: begin
            cosine_reg0 <= 36'sb101110110110010101011011111111111101;
            sine_reg0   <= 36'sb100100111111000000000110100011111000;
        end
        10814: begin
            cosine_reg0 <= 36'sb101110110110111111111000001110111111;
            sine_reg0   <= 36'sb100100111110100101001010110111111000;
        end
        10815: begin
            cosine_reg0 <= 36'sb101110110111101010010101001000010100;
            sine_reg0   <= 36'sb100100111110001010010000001110100100;
        end
        10816: begin
            cosine_reg0 <= 36'sb101110111000010100110010101011111010;
            sine_reg0   <= 36'sb100100111101101111010110100111111100;
        end
        10817: begin
            cosine_reg0 <= 36'sb101110111000111111010000111001101111;
            sine_reg0   <= 36'sb100100111101010100011110000100000001;
        end
        10818: begin
            cosine_reg0 <= 36'sb101110111001101001101111110001110010;
            sine_reg0   <= 36'sb100100111100111001100110100010110100;
        end
        10819: begin
            cosine_reg0 <= 36'sb101110111010010100001111010100000010;
            sine_reg0   <= 36'sb100100111100011110110000000100010111;
        end
        10820: begin
            cosine_reg0 <= 36'sb101110111010111110101111100000011100;
            sine_reg0   <= 36'sb100100111100000011111010101000101010;
        end
        10821: begin
            cosine_reg0 <= 36'sb101110111011101001010000010110111111;
            sine_reg0   <= 36'sb100100111011101001000110001111101110;
        end
        10822: begin
            cosine_reg0 <= 36'sb101110111100010011110001110111101001;
            sine_reg0   <= 36'sb100100111011001110010010111001100101;
        end
        10823: begin
            cosine_reg0 <= 36'sb101110111100111110010100000010011001;
            sine_reg0   <= 36'sb100100111010110011100000100110001111;
        end
        10824: begin
            cosine_reg0 <= 36'sb101110111101101000110110110111001100;
            sine_reg0   <= 36'sb100100111010011000101111010101101110;
        end
        10825: begin
            cosine_reg0 <= 36'sb101110111110010011011010010110000011;
            sine_reg0   <= 36'sb100100111001111101111111001000000010;
        end
        10826: begin
            cosine_reg0 <= 36'sb101110111110111101111110011110111001;
            sine_reg0   <= 36'sb100100111001100011001111111101001101;
        end
        10827: begin
            cosine_reg0 <= 36'sb101110111111101000100011010001101111;
            sine_reg0   <= 36'sb100100111001001000100001110101001111;
        end
        10828: begin
            cosine_reg0 <= 36'sb101111000000010011001000101110100011;
            sine_reg0   <= 36'sb100100111000101101110100110000001010;
        end
        10829: begin
            cosine_reg0 <= 36'sb101111000000111101101110110101010010;
            sine_reg0   <= 36'sb100100111000010011001000101101111111;
        end
        10830: begin
            cosine_reg0 <= 36'sb101111000001101000010101100101111011;
            sine_reg0   <= 36'sb100100110111111000011101101110101110;
        end
        10831: begin
            cosine_reg0 <= 36'sb101111000010010010111101000000011101;
            sine_reg0   <= 36'sb100100110111011101110011110010011001;
        end
        10832: begin
            cosine_reg0 <= 36'sb101111000010111101100101000100110110;
            sine_reg0   <= 36'sb100100110111000011001010111001000001;
        end
        10833: begin
            cosine_reg0 <= 36'sb101111000011101000001101110011000100;
            sine_reg0   <= 36'sb100100110110101000100011000010100110;
        end
        10834: begin
            cosine_reg0 <= 36'sb101111000100010010110111001011000101;
            sine_reg0   <= 36'sb100100110110001101111100001111001011;
        end
        10835: begin
            cosine_reg0 <= 36'sb101111000100111101100001001100111001;
            sine_reg0   <= 36'sb100100110101110011010110011110101111;
        end
        10836: begin
            cosine_reg0 <= 36'sb101111000101101000001011111000011101;
            sine_reg0   <= 36'sb100100110101011000110001110001010100;
        end
        10837: begin
            cosine_reg0 <= 36'sb101111000110010010110111001101101111;
            sine_reg0   <= 36'sb100100110100111110001110000110111010;
        end
        10838: begin
            cosine_reg0 <= 36'sb101111000110111101100011001100101110;
            sine_reg0   <= 36'sb100100110100100011101011011111100100;
        end
        10839: begin
            cosine_reg0 <= 36'sb101111000111101000001111110101011001;
            sine_reg0   <= 36'sb100100110100001001001001111011010010;
        end
        10840: begin
            cosine_reg0 <= 36'sb101111001000010010111101000111101110;
            sine_reg0   <= 36'sb100100110011101110101001011010000100;
        end
        10841: begin
            cosine_reg0 <= 36'sb101111001000111101101011000011101010;
            sine_reg0   <= 36'sb100100110011010100001001111011111100;
        end
        10842: begin
            cosine_reg0 <= 36'sb101111001001101000011001101001001101;
            sine_reg0   <= 36'sb100100110010111001101011100000111100;
        end
        10843: begin
            cosine_reg0 <= 36'sb101111001010010011001000111000010101;
            sine_reg0   <= 36'sb100100110010011111001110001001000011;
        end
        10844: begin
            cosine_reg0 <= 36'sb101111001010111101111000110001000000;
            sine_reg0   <= 36'sb100100110010000100110001110100010100;
        end
        10845: begin
            cosine_reg0 <= 36'sb101111001011101000101001010011001100;
            sine_reg0   <= 36'sb100100110001101010010110100010101110;
        end
        10846: begin
            cosine_reg0 <= 36'sb101111001100010011011010011110111000;
            sine_reg0   <= 36'sb100100110001001111111100010100010011;
        end
        10847: begin
            cosine_reg0 <= 36'sb101111001100111110001100010100000010;
            sine_reg0   <= 36'sb100100110000110101100011001001000101;
        end
        10848: begin
            cosine_reg0 <= 36'sb101111001101101000111110110010101001;
            sine_reg0   <= 36'sb100100110000011011001011000001000100;
        end
        10849: begin
            cosine_reg0 <= 36'sb101111001110010011110001111010101011;
            sine_reg0   <= 36'sb100100110000000000110011111100010000;
        end
        10850: begin
            cosine_reg0 <= 36'sb101111001110111110100101101100000110;
            sine_reg0   <= 36'sb100100101111100110011101111010101100;
        end
        10851: begin
            cosine_reg0 <= 36'sb101111001111101001011010000110111000;
            sine_reg0   <= 36'sb100100101111001100001000111100011000;
        end
        10852: begin
            cosine_reg0 <= 36'sb101111010000010100001111001011000001;
            sine_reg0   <= 36'sb100100101110110001110101000001010101;
        end
        10853: begin
            cosine_reg0 <= 36'sb101111010000111111000100111000011101;
            sine_reg0   <= 36'sb100100101110010111100010001001100100;
        end
        10854: begin
            cosine_reg0 <= 36'sb101111010001101001111011001111001101;
            sine_reg0   <= 36'sb100100101101111101010000010101000111;
        end
        10855: begin
            cosine_reg0 <= 36'sb101111010010010100110010001111001101;
            sine_reg0   <= 36'sb100100101101100010111111100011111101;
        end
        10856: begin
            cosine_reg0 <= 36'sb101111010010111111101001111000011101;
            sine_reg0   <= 36'sb100100101101001000101111110110001001;
        end
        10857: begin
            cosine_reg0 <= 36'sb101111010011101010100010001010111010;
            sine_reg0   <= 36'sb100100101100101110100001001011101011;
        end
        10858: begin
            cosine_reg0 <= 36'sb101111010100010101011011000110100011;
            sine_reg0   <= 36'sb100100101100010100010011100100100101;
        end
        10859: begin
            cosine_reg0 <= 36'sb101111010101000000010100101011010111;
            sine_reg0   <= 36'sb100100101011111010000111000000110110;
        end
        10860: begin
            cosine_reg0 <= 36'sb101111010101101011001110111001010011;
            sine_reg0   <= 36'sb100100101011011111111011100000100001;
        end
        10861: begin
            cosine_reg0 <= 36'sb101111010110010110001001110000010111;
            sine_reg0   <= 36'sb100100101011000101110001000011100110;
        end
        10862: begin
            cosine_reg0 <= 36'sb101111010111000001000101010000011111;
            sine_reg0   <= 36'sb100100101010101011100111101010000110;
        end
        10863: begin
            cosine_reg0 <= 36'sb101111010111101100000001011001101100;
            sine_reg0   <= 36'sb100100101010010001011111010100000011;
        end
        10864: begin
            cosine_reg0 <= 36'sb101111011000010110111110001011111011;
            sine_reg0   <= 36'sb100100101001110111011000000001011100;
        end
        10865: begin
            cosine_reg0 <= 36'sb101111011001000001111011100111001010;
            sine_reg0   <= 36'sb100100101001011101010001110010010100;
        end
        10866: begin
            cosine_reg0 <= 36'sb101111011001101100111001101011010111;
            sine_reg0   <= 36'sb100100101001000011001100100110101100;
        end
        10867: begin
            cosine_reg0 <= 36'sb101111011010010111111000011000100010;
            sine_reg0   <= 36'sb100100101000101001001000011110100011;
        end
        10868: begin
            cosine_reg0 <= 36'sb101111011011000010110111101110101001;
            sine_reg0   <= 36'sb100100101000001111000101011001111100;
        end
        10869: begin
            cosine_reg0 <= 36'sb101111011011101101110111101101101001;
            sine_reg0   <= 36'sb100100100111110101000011011000111000;
        end
        10870: begin
            cosine_reg0 <= 36'sb101111011100011000111000010101100001;
            sine_reg0   <= 36'sb100100100111011011000010011011010110;
        end
        10871: begin
            cosine_reg0 <= 36'sb101111011101000011111001100110010000;
            sine_reg0   <= 36'sb100100100111000001000010100001011001;
        end
        10872: begin
            cosine_reg0 <= 36'sb101111011101101110111011011111110100;
            sine_reg0   <= 36'sb100100100110100111000011101011000001;
        end
        10873: begin
            cosine_reg0 <= 36'sb101111011110011001111110000010001011;
            sine_reg0   <= 36'sb100100100110001101000101111000010000;
        end
        10874: begin
            cosine_reg0 <= 36'sb101111011111000101000001001101010011;
            sine_reg0   <= 36'sb100100100101110011001001001001000110;
        end
        10875: begin
            cosine_reg0 <= 36'sb101111011111110000000101000001001011;
            sine_reg0   <= 36'sb100100100101011001001101011101100100;
        end
        10876: begin
            cosine_reg0 <= 36'sb101111100000011011001001011101110010;
            sine_reg0   <= 36'sb100100100100111111010010110101101011;
        end
        10877: begin
            cosine_reg0 <= 36'sb101111100001000110001110100011000100;
            sine_reg0   <= 36'sb100100100100100101011001010001011101;
        end
        10878: begin
            cosine_reg0 <= 36'sb101111100001110001010100010001000010;
            sine_reg0   <= 36'sb100100100100001011100000110000111010;
        end
        10879: begin
            cosine_reg0 <= 36'sb101111100010011100011010100111101001;
            sine_reg0   <= 36'sb100100100011110001101001010100000100;
        end
        10880: begin
            cosine_reg0 <= 36'sb101111100011000111100001100110111000;
            sine_reg0   <= 36'sb100100100011010111110010111010111011;
        end
        10881: begin
            cosine_reg0 <= 36'sb101111100011110010101001001110101100;
            sine_reg0   <= 36'sb100100100010111101111101100101100000;
        end
        10882: begin
            cosine_reg0 <= 36'sb101111100100011101110001011111000101;
            sine_reg0   <= 36'sb100100100010100100001001010011110100;
        end
        10883: begin
            cosine_reg0 <= 36'sb101111100101001000111010011000000000;
            sine_reg0   <= 36'sb100100100010001010010110000101111001;
        end
        10884: begin
            cosine_reg0 <= 36'sb101111100101110100000011111001011100;
            sine_reg0   <= 36'sb100100100001110000100011111011101110;
        end
        10885: begin
            cosine_reg0 <= 36'sb101111100110011111001110000011010111;
            sine_reg0   <= 36'sb100100100001010110110010110101010111;
        end
        10886: begin
            cosine_reg0 <= 36'sb101111100111001010011000110101110000;
            sine_reg0   <= 36'sb100100100000111101000010110010110010;
        end
        10887: begin
            cosine_reg0 <= 36'sb101111100111110101100100010000100101;
            sine_reg0   <= 36'sb100100100000100011010011110100000010;
        end
        10888: begin
            cosine_reg0 <= 36'sb101111101000100000110000010011110100;
            sine_reg0   <= 36'sb100100100000001001100101111001000111;
        end
        10889: begin
            cosine_reg0 <= 36'sb101111101001001011111100111111011100;
            sine_reg0   <= 36'sb100100011111101111111001000010000010;
        end
        10890: begin
            cosine_reg0 <= 36'sb101111101001110111001010010011011010;
            sine_reg0   <= 36'sb100100011111010110001101001110110101;
        end
        10891: begin
            cosine_reg0 <= 36'sb101111101010100010011000001111101110;
            sine_reg0   <= 36'sb100100011110111100100010011111100000;
        end
        10892: begin
            cosine_reg0 <= 36'sb101111101011001101100110110100010101;
            sine_reg0   <= 36'sb100100011110100010111000110100000100;
        end
        10893: begin
            cosine_reg0 <= 36'sb101111101011111000110110000001001110;
            sine_reg0   <= 36'sb100100011110001001010000001100100010;
        end
        10894: begin
            cosine_reg0 <= 36'sb101111101100100100000101110110011000;
            sine_reg0   <= 36'sb100100011101101111101000101000111011;
        end
        10895: begin
            cosine_reg0 <= 36'sb101111101101001111010110010011110000;
            sine_reg0   <= 36'sb100100011101010110000010001001010001;
        end
        10896: begin
            cosine_reg0 <= 36'sb101111101101111010100111011001010101;
            sine_reg0   <= 36'sb100100011100111100011100101101100100;
        end
        10897: begin
            cosine_reg0 <= 36'sb101111101110100101111001000111000101;
            sine_reg0   <= 36'sb100100011100100010111000010101110101;
        end
        10898: begin
            cosine_reg0 <= 36'sb101111101111010001001011011100111111;
            sine_reg0   <= 36'sb100100011100001001010101000010000101;
        end
        10899: begin
            cosine_reg0 <= 36'sb101111101111111100011110011011000001;
            sine_reg0   <= 36'sb100100011011101111110010110010010101;
        end
        10900: begin
            cosine_reg0 <= 36'sb101111110000100111110010000001001001;
            sine_reg0   <= 36'sb100100011011010110010001100110100110;
        end
        10901: begin
            cosine_reg0 <= 36'sb101111110001010011000110001111010101;
            sine_reg0   <= 36'sb100100011010111100110001011110111010;
        end
        10902: begin
            cosine_reg0 <= 36'sb101111110001111110011011000101100100;
            sine_reg0   <= 36'sb100100011010100011010010011011010000;
        end
        10903: begin
            cosine_reg0 <= 36'sb101111110010101001110000100011110101;
            sine_reg0   <= 36'sb100100011010001001110100011011101011;
        end
        10904: begin
            cosine_reg0 <= 36'sb101111110011010101000110101010000101;
            sine_reg0   <= 36'sb100100011001110000010111100000001011;
        end
        10905: begin
            cosine_reg0 <= 36'sb101111110100000000011101011000010011;
            sine_reg0   <= 36'sb100100011001010110111011101000110000;
        end
        10906: begin
            cosine_reg0 <= 36'sb101111110100101011110100101110011101;
            sine_reg0   <= 36'sb100100011000111101100000110101011101;
        end
        10907: begin
            cosine_reg0 <= 36'sb101111110101010111001100101100100010;
            sine_reg0   <= 36'sb100100011000100100000111000110010010;
        end
        10908: begin
            cosine_reg0 <= 36'sb101111110110000010100101010010100000;
            sine_reg0   <= 36'sb100100011000001010101110011011001111;
        end
        10909: begin
            cosine_reg0 <= 36'sb101111110110101101111110100000010101;
            sine_reg0   <= 36'sb100100010111110001010110110100010111;
        end
        10910: begin
            cosine_reg0 <= 36'sb101111110111011001011000010101111111;
            sine_reg0   <= 36'sb100100010111011000000000010001101010;
        end
        10911: begin
            cosine_reg0 <= 36'sb101111111000000100110010110011011101;
            sine_reg0   <= 36'sb100100010110111110101010110011001000;
        end
        10912: begin
            cosine_reg0 <= 36'sb101111111000110000001101111000101101;
            sine_reg0   <= 36'sb100100010110100101010110011000110011;
        end
        10913: begin
            cosine_reg0 <= 36'sb101111111001011011101001100101101110;
            sine_reg0   <= 36'sb100100010110001100000011000010101101;
        end
        10914: begin
            cosine_reg0 <= 36'sb101111111010000111000101111010011110;
            sine_reg0   <= 36'sb100100010101110010110000110000110101;
        end
        10915: begin
            cosine_reg0 <= 36'sb101111111010110010100010110110111011;
            sine_reg0   <= 36'sb100100010101011001011111100011001101;
        end
        10916: begin
            cosine_reg0 <= 36'sb101111111011011110000000011011000011;
            sine_reg0   <= 36'sb100100010101000000001111011001110101;
        end
        10917: begin
            cosine_reg0 <= 36'sb101111111100001001011110100110110101;
            sine_reg0   <= 36'sb100100010100100111000000010100110000;
        end
        10918: begin
            cosine_reg0 <= 36'sb101111111100110100111101011010001111;
            sine_reg0   <= 36'sb100100010100001101110010010011111101;
        end
        10919: begin
            cosine_reg0 <= 36'sb101111111101100000011100110101010000;
            sine_reg0   <= 36'sb100100010011110100100101010111011110;
        end
        10920: begin
            cosine_reg0 <= 36'sb101111111110001011111100110111110110;
            sine_reg0   <= 36'sb100100010011011011011001011111010011;
        end
        10921: begin
            cosine_reg0 <= 36'sb101111111110110111011101100001111110;
            sine_reg0   <= 36'sb100100010011000010001110101011011110;
        end
        10922: begin
            cosine_reg0 <= 36'sb101111111111100010111110110011101000;
            sine_reg0   <= 36'sb100100010010101001000100111100000000;
        end
        10923: begin
            cosine_reg0 <= 36'sb110000000000001110100000101100110010;
            sine_reg0   <= 36'sb100100010010001111111100010000111001;
        end
        10924: begin
            cosine_reg0 <= 36'sb110000000000111010000011001101011010;
            sine_reg0   <= 36'sb100100010001110110110100101010001011;
        end
        10925: begin
            cosine_reg0 <= 36'sb110000000001100101100110010101011110;
            sine_reg0   <= 36'sb100100010001011101101110000111110111;
        end
        10926: begin
            cosine_reg0 <= 36'sb110000000010010001001010000100111101;
            sine_reg0   <= 36'sb100100010001000100101000101001111101;
        end
        10927: begin
            cosine_reg0 <= 36'sb110000000010111100101110011011110100;
            sine_reg0   <= 36'sb100100010000101011100100010000011110;
        end
        10928: begin
            cosine_reg0 <= 36'sb110000000011101000010011011010000100;
            sine_reg0   <= 36'sb100100010000010010100000111011011100;
        end
        10929: begin
            cosine_reg0 <= 36'sb110000000100010011111000111111101000;
            sine_reg0   <= 36'sb100100001111111001011110101010110111;
        end
        10930: begin
            cosine_reg0 <= 36'sb110000000100111111011111001100100001;
            sine_reg0   <= 36'sb100100001111100000011101011110110001;
        end
        10931: begin
            cosine_reg0 <= 36'sb110000000101101011000110000000101100;
            sine_reg0   <= 36'sb100100001111000111011101010111001010;
        end
        10932: begin
            cosine_reg0 <= 36'sb110000000110010110101101011100001000;
            sine_reg0   <= 36'sb100100001110101110011110010100000011;
        end
        10933: begin
            cosine_reg0 <= 36'sb110000000111000010010101011110110011;
            sine_reg0   <= 36'sb100100001110010101100000010101011101;
        end
        10934: begin
            cosine_reg0 <= 36'sb110000000111101101111110001000101011;
            sine_reg0   <= 36'sb100100001101111100100011011011011010;
        end
        10935: begin
            cosine_reg0 <= 36'sb110000001000011001100111011001101110;
            sine_reg0   <= 36'sb100100001101100011100111100101111010;
        end
        10936: begin
            cosine_reg0 <= 36'sb110000001001000101010001010001111100;
            sine_reg0   <= 36'sb100100001101001010101100110100111110;
        end
        10937: begin
            cosine_reg0 <= 36'sb110000001001110000111011110001010010;
            sine_reg0   <= 36'sb100100001100110001110011001000100111;
        end
        10938: begin
            cosine_reg0 <= 36'sb110000001010011100100110110111101110;
            sine_reg0   <= 36'sb100100001100011000111010100000110110;
        end
        10939: begin
            cosine_reg0 <= 36'sb110000001011001000010010100101001111;
            sine_reg0   <= 36'sb100100001100000000000010111101101100;
        end
        10940: begin
            cosine_reg0 <= 36'sb110000001011110011111110111001110011;
            sine_reg0   <= 36'sb100100001011100111001100011111001010;
        end
        10941: begin
            cosine_reg0 <= 36'sb110000001100011111101011110101011001;
            sine_reg0   <= 36'sb100100001011001110010111000101010001;
        end
        10942: begin
            cosine_reg0 <= 36'sb110000001101001011011001010111111110;
            sine_reg0   <= 36'sb100100001010110101100010110000000010;
        end
        10943: begin
            cosine_reg0 <= 36'sb110000001101110111000111100001100001;
            sine_reg0   <= 36'sb100100001010011100101111011111011101;
        end
        10944: begin
            cosine_reg0 <= 36'sb110000001110100010110110010010000001;
            sine_reg0   <= 36'sb100100001010000011111101010011100101;
        end
        10945: begin
            cosine_reg0 <= 36'sb110000001111001110100101101001011100;
            sine_reg0   <= 36'sb100100001001101011001100001100011001;
        end
        10946: begin
            cosine_reg0 <= 36'sb110000001111111010010101100111110000;
            sine_reg0   <= 36'sb100100001001010010011100001001111011;
        end
        10947: begin
            cosine_reg0 <= 36'sb110000010000100110000110001100111011;
            sine_reg0   <= 36'sb100100001000111001101101001100001100;
        end
        10948: begin
            cosine_reg0 <= 36'sb110000010001010001110111011000111100;
            sine_reg0   <= 36'sb100100001000100000111111010011001100;
        end
        10949: begin
            cosine_reg0 <= 36'sb110000010001111101101001001011110000;
            sine_reg0   <= 36'sb100100001000001000010010011110111101;
        end
        10950: begin
            cosine_reg0 <= 36'sb110000010010101001011011100101010111;
            sine_reg0   <= 36'sb100100000111101111100110101111011111;
        end
        10951: begin
            cosine_reg0 <= 36'sb110000010011010101001110100101101111;
            sine_reg0   <= 36'sb100100000111010110111100000100110100;
        end
        10952: begin
            cosine_reg0 <= 36'sb110000010100000001000010001100110110;
            sine_reg0   <= 36'sb100100000110111110010010011110111101;
        end
        10953: begin
            cosine_reg0 <= 36'sb110000010100101100110110011010101001;
            sine_reg0   <= 36'sb100100000110100101101001111101111001;
        end
        10954: begin
            cosine_reg0 <= 36'sb110000010101011000101011001111001001;
            sine_reg0   <= 36'sb100100000110001101000010100001101011;
        end
        10955: begin
            cosine_reg0 <= 36'sb110000010110000100100000101010010010;
            sine_reg0   <= 36'sb100100000101110100011100001010010011;
        end
        10956: begin
            cosine_reg0 <= 36'sb110000010110110000010110101100000011;
            sine_reg0   <= 36'sb100100000101011011110110110111110011;
        end
        10957: begin
            cosine_reg0 <= 36'sb110000010111011100001101010100011011;
            sine_reg0   <= 36'sb100100000101000011010010101010001011;
        end
        10958: begin
            cosine_reg0 <= 36'sb110000011000001000000100100011011000;
            sine_reg0   <= 36'sb100100000100101010101111100001011011;
        end
        10959: begin
            cosine_reg0 <= 36'sb110000011000110011111100011000110111;
            sine_reg0   <= 36'sb100100000100010010001101011101100110;
        end
        10960: begin
            cosine_reg0 <= 36'sb110000011001011111110100110100111001;
            sine_reg0   <= 36'sb100100000011111001101100011110101100;
        end
        10961: begin
            cosine_reg0 <= 36'sb110000011010001011101101110111011001;
            sine_reg0   <= 36'sb100100000011100001001100100100101110;
        end
        10962: begin
            cosine_reg0 <= 36'sb110000011010110111100111100000011000;
            sine_reg0   <= 36'sb100100000011001000101101101111101101;
        end
        10963: begin
            cosine_reg0 <= 36'sb110000011011100011100001101111110011;
            sine_reg0   <= 36'sb100100000010110000001111111111101001;
        end
        10964: begin
            cosine_reg0 <= 36'sb110000011100001111011100100101101001;
            sine_reg0   <= 36'sb100100000010010111110011010100100100;
        end
        10965: begin
            cosine_reg0 <= 36'sb110000011100111011011000000001111000;
            sine_reg0   <= 36'sb100100000001111111010111101110011111;
        end
        10966: begin
            cosine_reg0 <= 36'sb110000011101100111010100000100011110;
            sine_reg0   <= 36'sb100100000001100110111101001101011011;
        end
        10967: begin
            cosine_reg0 <= 36'sb110000011110010011010000101101011001;
            sine_reg0   <= 36'sb100100000001001110100011110001011001;
        end
        10968: begin
            cosine_reg0 <= 36'sb110000011110111111001101111100101000;
            sine_reg0   <= 36'sb100100000000110110001011011010011000;
        end
        10969: begin
            cosine_reg0 <= 36'sb110000011111101011001011110010001010;
            sine_reg0   <= 36'sb100100000000011101110100001000011100;
        end
        10970: begin
            cosine_reg0 <= 36'sb110000100000010111001010001101111100;
            sine_reg0   <= 36'sb100100000000000101011101111011100100;
        end
        10971: begin
            cosine_reg0 <= 36'sb110000100001000011001001001111111101;
            sine_reg0   <= 36'sb100011111111101101001000110011110001;
        end
        10972: begin
            cosine_reg0 <= 36'sb110000100001101111001000111000001011;
            sine_reg0   <= 36'sb100011111111010100110100110001000100;
        end
        10973: begin
            cosine_reg0 <= 36'sb110000100010011011001001000110100100;
            sine_reg0   <= 36'sb100011111110111100100001110011011111;
        end
        10974: begin
            cosine_reg0 <= 36'sb110000100011000111001001111011000111;
            sine_reg0   <= 36'sb100011111110100100001111111011000010;
        end
        10975: begin
            cosine_reg0 <= 36'sb110000100011110011001011010101110001;
            sine_reg0   <= 36'sb100011111110001011111111000111101110;
        end
        10976: begin
            cosine_reg0 <= 36'sb110000100100011111001101010110100011;
            sine_reg0   <= 36'sb100011111101110011101111011001100100;
        end
        10977: begin
            cosine_reg0 <= 36'sb110000100101001011001111111101011000;
            sine_reg0   <= 36'sb100011111101011011100000110000100101;
        end
        10978: begin
            cosine_reg0 <= 36'sb110000100101110111010011001010010001;
            sine_reg0   <= 36'sb100011111101000011010011001100110010;
        end
        10979: begin
            cosine_reg0 <= 36'sb110000100110100011010110111101001011;
            sine_reg0   <= 36'sb100011111100101011000110101110001100;
        end
        10980: begin
            cosine_reg0 <= 36'sb110000100111001111011011010110000100;
            sine_reg0   <= 36'sb100011111100010010111011010100110100;
        end
        10981: begin
            cosine_reg0 <= 36'sb110000100111111011100000010100111011;
            sine_reg0   <= 36'sb100011111011111010110001000000101010;
        end
        10982: begin
            cosine_reg0 <= 36'sb110000101000100111100101111001101110;
            sine_reg0   <= 36'sb100011111011100010100111110001110000;
        end
        10983: begin
            cosine_reg0 <= 36'sb110000101001010011101100000100011100;
            sine_reg0   <= 36'sb100011111011001010011111101000000111;
        end
        10984: begin
            cosine_reg0 <= 36'sb110000101001111111110010110101000010;
            sine_reg0   <= 36'sb100011111010110010011000100011101111;
        end
        10985: begin
            cosine_reg0 <= 36'sb110000101010101011111010001011011111;
            sine_reg0   <= 36'sb100011111010011010010010100100101010;
        end
        10986: begin
            cosine_reg0 <= 36'sb110000101011011000000010000111110010;
            sine_reg0   <= 36'sb100011111010000010001101101010111000;
        end
        10987: begin
            cosine_reg0 <= 36'sb110000101100000100001010101001111000;
            sine_reg0   <= 36'sb100011111001101010001001110110011010;
        end
        10988: begin
            cosine_reg0 <= 36'sb110000101100110000010011110001110000;
            sine_reg0   <= 36'sb100011111001010010000111000111010010;
        end
        10989: begin
            cosine_reg0 <= 36'sb110000101101011100011101011111011001;
            sine_reg0   <= 36'sb100011111000111010000101011101011111;
        end
        10990: begin
            cosine_reg0 <= 36'sb110000101110001000100111110010101111;
            sine_reg0   <= 36'sb100011111000100010000100111001000100;
        end
        10991: begin
            cosine_reg0 <= 36'sb110000101110110100110010101011110011;
            sine_reg0   <= 36'sb100011111000001010000101011010000001;
        end
        10992: begin
            cosine_reg0 <= 36'sb110000101111100000111110001010100001;
            sine_reg0   <= 36'sb100011110111110010000111000000010111;
        end
        10993: begin
            cosine_reg0 <= 36'sb110000110000001101001010001110111001;
            sine_reg0   <= 36'sb100011110111011010001001101100000110;
        end
        10994: begin
            cosine_reg0 <= 36'sb110000110000111001010110111000111001;
            sine_reg0   <= 36'sb100011110111000010001101011101010000;
        end
        10995: begin
            cosine_reg0 <= 36'sb110000110001100101100100001000011111;
            sine_reg0   <= 36'sb100011110110101010010010010011110110;
        end
        10996: begin
            cosine_reg0 <= 36'sb110000110010010001110001111101101001;
            sine_reg0   <= 36'sb100011110110010010011000001111111001;
        end
        10997: begin
            cosine_reg0 <= 36'sb110000110010111110000000011000010101;
            sine_reg0   <= 36'sb100011110101111010011111010001011001;
        end
        10998: begin
            cosine_reg0 <= 36'sb110000110011101010001111011000100010;
            sine_reg0   <= 36'sb100011110101100010100111011000011000;
        end
        10999: begin
            cosine_reg0 <= 36'sb110000110100010110011110111110001111;
            sine_reg0   <= 36'sb100011110101001010110000100100110110;
        end
        11000: begin
            cosine_reg0 <= 36'sb110000110101000010101111001001011001;
            sine_reg0   <= 36'sb100011110100110010111010110110110100;
        end
        11001: begin
            cosine_reg0 <= 36'sb110000110101101110111111111001111111;
            sine_reg0   <= 36'sb100011110100011011000110001110010100;
        end
        11002: begin
            cosine_reg0 <= 36'sb110000110110011011010001001111111110;
            sine_reg0   <= 36'sb100011110100000011010010101011010110;
        end
        11003: begin
            cosine_reg0 <= 36'sb110000110111000111100011001011010110;
            sine_reg0   <= 36'sb100011110011101011100000001101111011;
        end
        11004: begin
            cosine_reg0 <= 36'sb110000110111110011110101101100000101;
            sine_reg0   <= 36'sb100011110011010011101110110110000011;
        end
        11005: begin
            cosine_reg0 <= 36'sb110000111000100000001000110010001001;
            sine_reg0   <= 36'sb100011110010111011111110100011110001;
        end
        11006: begin
            cosine_reg0 <= 36'sb110000111001001100011100011101011111;
            sine_reg0   <= 36'sb100011110010100100001111010111000101;
        end
        11007: begin
            cosine_reg0 <= 36'sb110000111001111000110000101110001000;
            sine_reg0   <= 36'sb100011110010001100100001001111111111;
        end
        11008: begin
            cosine_reg0 <= 36'sb110000111010100101000101100100000000;
            sine_reg0   <= 36'sb100011110001110100110100001110100001;
        end
        11009: begin
            cosine_reg0 <= 36'sb110000111011010001011010111111000110;
            sine_reg0   <= 36'sb100011110001011101001000010010101011;
        end
        11010: begin
            cosine_reg0 <= 36'sb110000111011111101110000111111011000;
            sine_reg0   <= 36'sb100011110001000101011101011100011111;
        end
        11011: begin
            cosine_reg0 <= 36'sb110000111100101010000111100100110101;
            sine_reg0   <= 36'sb100011110000101101110011101011111101;
        end
        11012: begin
            cosine_reg0 <= 36'sb110000111101010110011110101111011100;
            sine_reg0   <= 36'sb100011110000010110001011000001000111;
        end
        11013: begin
            cosine_reg0 <= 36'sb110000111110000010110110011111001001;
            sine_reg0   <= 36'sb100011101111111110100011011011111101;
        end
        11014: begin
            cosine_reg0 <= 36'sb110000111110101111001110110011111100;
            sine_reg0   <= 36'sb100011101111100110111100111100100000;
        end
        11015: begin
            cosine_reg0 <= 36'sb110000111111011011100111101101110010;
            sine_reg0   <= 36'sb100011101111001111010111100010110001;
        end
        11016: begin
            cosine_reg0 <= 36'sb110001000000001000000001001100101011;
            sine_reg0   <= 36'sb100011101110110111110011001110110000;
        end
        11017: begin
            cosine_reg0 <= 36'sb110001000000110100011011010000100101;
            sine_reg0   <= 36'sb100011101110100000010000000000100000;
        end
        11018: begin
            cosine_reg0 <= 36'sb110001000001100000110101111001011100;
            sine_reg0   <= 36'sb100011101110001000101101111000000001;
        end
        11019: begin
            cosine_reg0 <= 36'sb110001000010001101010001000111010001;
            sine_reg0   <= 36'sb100011101101110001001100110101010011;
        end
        11020: begin
            cosine_reg0 <= 36'sb110001000010111001101100111010000001;
            sine_reg0   <= 36'sb100011101101011001101100111000010111;
        end
        11021: begin
            cosine_reg0 <= 36'sb110001000011100110001001010001101011;
            sine_reg0   <= 36'sb100011101101000010001110000001010000;
        end
        11022: begin
            cosine_reg0 <= 36'sb110001000100010010100110001110001101;
            sine_reg0   <= 36'sb100011101100101010110000001111111100;
        end
        11023: begin
            cosine_reg0 <= 36'sb110001000100111111000011101111100100;
            sine_reg0   <= 36'sb100011101100010011010011100100011110;
        end
        11024: begin
            cosine_reg0 <= 36'sb110001000101101011100001110101110000;
            sine_reg0   <= 36'sb100011101011111011110111111110110110;
        end
        11025: begin
            cosine_reg0 <= 36'sb110001000110011000000000100000101111;
            sine_reg0   <= 36'sb100011101011100100011101011111000101;
        end
        11026: begin
            cosine_reg0 <= 36'sb110001000111000100011111110000011111;
            sine_reg0   <= 36'sb100011101011001101000100000101001100;
        end
        11027: begin
            cosine_reg0 <= 36'sb110001000111110000111111100100111110;
            sine_reg0   <= 36'sb100011101010110101101011110001001100;
        end
        11028: begin
            cosine_reg0 <= 36'sb110001001000011101011111111110001010;
            sine_reg0   <= 36'sb100011101010011110010100100011000110;
        end
        11029: begin
            cosine_reg0 <= 36'sb110001001001001010000000111100000010;
            sine_reg0   <= 36'sb100011101010000110111110011010111011;
        end
        11030: begin
            cosine_reg0 <= 36'sb110001001001110110100010011110100101;
            sine_reg0   <= 36'sb100011101001101111101001011000101011;
        end
        11031: begin
            cosine_reg0 <= 36'sb110001001010100011000100100101110000;
            sine_reg0   <= 36'sb100011101001011000010101011100010111;
        end
        11032: begin
            cosine_reg0 <= 36'sb110001001011001111100111010001100001;
            sine_reg0   <= 36'sb100011101001000001000010100110000001;
        end
        11033: begin
            cosine_reg0 <= 36'sb110001001011111100001010100001111000;
            sine_reg0   <= 36'sb100011101000101001110000110101101001;
        end
        11034: begin
            cosine_reg0 <= 36'sb110001001100101000101110010110110001;
            sine_reg0   <= 36'sb100011101000010010100000001011010001;
        end
        11035: begin
            cosine_reg0 <= 36'sb110001001101010101010010110000001101;
            sine_reg0   <= 36'sb100011100111111011010000100110111000;
        end
        11036: begin
            cosine_reg0 <= 36'sb110001001110000001110111101110001000;
            sine_reg0   <= 36'sb100011100111100100000010001000100001;
        end
        11037: begin
            cosine_reg0 <= 36'sb110001001110101110011101010000100001;
            sine_reg0   <= 36'sb100011100111001100110100110000001011;
        end
        11038: begin
            cosine_reg0 <= 36'sb110001001111011011000011010111010110;
            sine_reg0   <= 36'sb100011100110110101101000011101111001;
        end
        11039: begin
            cosine_reg0 <= 36'sb110001010000000111101010000010100111;
            sine_reg0   <= 36'sb100011100110011110011101010001101001;
        end
        11040: begin
            cosine_reg0 <= 36'sb110001010000110100010001010010010000;
            sine_reg0   <= 36'sb100011100110000111010011001011011111;
        end
        11041: begin
            cosine_reg0 <= 36'sb110001010001100000111001000110010000;
            sine_reg0   <= 36'sb100011100101110000001010001011011010;
        end
        11042: begin
            cosine_reg0 <= 36'sb110001010010001101100001011110100110;
            sine_reg0   <= 36'sb100011100101011001000010010001011011;
        end
        11043: begin
            cosine_reg0 <= 36'sb110001010010111010001010011011001111;
            sine_reg0   <= 36'sb100011100101000001111011011101100011;
        end
        11044: begin
            cosine_reg0 <= 36'sb110001010011100110110011111100001011;
            sine_reg0   <= 36'sb100011100100101010110101101111110100;
        end
        11045: begin
            cosine_reg0 <= 36'sb110001010100010011011110000001010111;
            sine_reg0   <= 36'sb100011100100010011110001001000001101;
        end
        11046: begin
            cosine_reg0 <= 36'sb110001010101000000001000101010110001;
            sine_reg0   <= 36'sb100011100011111100101101100110110001;
        end
        11047: begin
            cosine_reg0 <= 36'sb110001010101101100110011111000011001;
            sine_reg0   <= 36'sb100011100011100101101011001011011111;
        end
        11048: begin
            cosine_reg0 <= 36'sb110001010110011001011111101010001011;
            sine_reg0   <= 36'sb100011100011001110101001110110011001;
        end
        11049: begin
            cosine_reg0 <= 36'sb110001010111000110001100000000000111;
            sine_reg0   <= 36'sb100011100010110111101001100111100000;
        end
        11050: begin
            cosine_reg0 <= 36'sb110001010111110010111000111010001011;
            sine_reg0   <= 36'sb100011100010100000101010011110110100;
        end
        11051: begin
            cosine_reg0 <= 36'sb110001011000011111100110011000010101;
            sine_reg0   <= 36'sb100011100010001001101100011100010110;
        end
        11052: begin
            cosine_reg0 <= 36'sb110001011001001100010100011010100011;
            sine_reg0   <= 36'sb100011100001110010101111100000001000;
        end
        11053: begin
            cosine_reg0 <= 36'sb110001011001111001000011000000110100;
            sine_reg0   <= 36'sb100011100001011011110011101010001001;
        end
        11054: begin
            cosine_reg0 <= 36'sb110001011010100101110010001011000101;
            sine_reg0   <= 36'sb100011100001000100111000111010011100;
        end
        11055: begin
            cosine_reg0 <= 36'sb110001011011010010100001111001010101;
            sine_reg0   <= 36'sb100011100000101101111111010001000001;
        end
        11056: begin
            cosine_reg0 <= 36'sb110001011011111111010010001011100011;
            sine_reg0   <= 36'sb100011100000010111000110101101111000;
        end
        11057: begin
            cosine_reg0 <= 36'sb110001011100101100000011000001101101;
            sine_reg0   <= 36'sb100011100000000000001111010001000011;
        end
        11058: begin
            cosine_reg0 <= 36'sb110001011101011000110100011011110000;
            sine_reg0   <= 36'sb100011011111101001011000111010100011;
        end
        11059: begin
            cosine_reg0 <= 36'sb110001011110000101100110011001101100;
            sine_reg0   <= 36'sb100011011111010010100011101010011000;
        end
        11060: begin
            cosine_reg0 <= 36'sb110001011110110010011000111011011110;
            sine_reg0   <= 36'sb100011011110111011101111100000100011;
        end
        11061: begin
            cosine_reg0 <= 36'sb110001011111011111001100000001000101;
            sine_reg0   <= 36'sb100011011110100100111100011101000101;
        end
        11062: begin
            cosine_reg0 <= 36'sb110001100000001011111111101010011110;
            sine_reg0   <= 36'sb100011011110001110001010100000000000;
        end
        11063: begin
            cosine_reg0 <= 36'sb110001100000111000110011110111101010;
            sine_reg0   <= 36'sb100011011101110111011001101001010011;
        end
        11064: begin
            cosine_reg0 <= 36'sb110001100001100101101000101000100100;
            sine_reg0   <= 36'sb100011011101100000101001111001000000;
        end
        11065: begin
            cosine_reg0 <= 36'sb110001100010010010011101111101001101;
            sine_reg0   <= 36'sb100011011101001001111011001111001000;
        end
        11066: begin
            cosine_reg0 <= 36'sb110001100010111111010011110101100001;
            sine_reg0   <= 36'sb100011011100110011001101101011101100;
        end
        11067: begin
            cosine_reg0 <= 36'sb110001100011101100001010010001100000;
            sine_reg0   <= 36'sb100011011100011100100001001110101011;
        end
        11068: begin
            cosine_reg0 <= 36'sb110001100100011001000001010001001000;
            sine_reg0   <= 36'sb100011011100000101110101111000001001;
        end
        11069: begin
            cosine_reg0 <= 36'sb110001100101000101111000110100010110;
            sine_reg0   <= 36'sb100011011011101111001011101000000100;
        end
        11070: begin
            cosine_reg0 <= 36'sb110001100101110010110000111011001010;
            sine_reg0   <= 36'sb100011011011011000100010011110011110;
        end
        11071: begin
            cosine_reg0 <= 36'sb110001100110011111101001100101100001;
            sine_reg0   <= 36'sb100011011011000001111010011011011001;
        end
        11072: begin
            cosine_reg0 <= 36'sb110001100111001100100010110011011010;
            sine_reg0   <= 36'sb100011011010101011010011011110110100;
        end
        11073: begin
            cosine_reg0 <= 36'sb110001100111111001011100100100110011;
            sine_reg0   <= 36'sb100011011010010100101101101000110001;
        end
        11074: begin
            cosine_reg0 <= 36'sb110001101000100110010110111001101010;
            sine_reg0   <= 36'sb100011011001111110001000111001010000;
        end
        11075: begin
            cosine_reg0 <= 36'sb110001101001010011010001110001111110;
            sine_reg0   <= 36'sb100011011001100111100101010000010011;
        end
        11076: begin
            cosine_reg0 <= 36'sb110001101010000000001101001101101100;
            sine_reg0   <= 36'sb100011011001010001000010101101111010;
        end
        11077: begin
            cosine_reg0 <= 36'sb110001101010101101001001001100110100;
            sine_reg0   <= 36'sb100011011000111010100001010010000110;
        end
        11078: begin
            cosine_reg0 <= 36'sb110001101011011010000101101111010011;
            sine_reg0   <= 36'sb100011011000100100000000111100111000;
        end
        11079: begin
            cosine_reg0 <= 36'sb110001101100000111000010110101000111;
            sine_reg0   <= 36'sb100011011000001101100001101110010010;
        end
        11080: begin
            cosine_reg0 <= 36'sb110001101100110100000000011110010000;
            sine_reg0   <= 36'sb100011010111110111000011100110010010;
        end
        11081: begin
            cosine_reg0 <= 36'sb110001101101100000111110101010101010;
            sine_reg0   <= 36'sb100011010111100000100110100100111100;
        end
        11082: begin
            cosine_reg0 <= 36'sb110001101110001101111101011010010101;
            sine_reg0   <= 36'sb100011010111001010001010101010001111;
        end
        11083: begin
            cosine_reg0 <= 36'sb110001101110111010111100101101001111;
            sine_reg0   <= 36'sb100011010110110011101111110110001100;
        end
        11084: begin
            cosine_reg0 <= 36'sb110001101111100111111100100011010101;
            sine_reg0   <= 36'sb100011010110011101010110001000110101;
        end
        11085: begin
            cosine_reg0 <= 36'sb110001110000010100111100111100100111;
            sine_reg0   <= 36'sb100011010110000110111101100010001010;
        end
        11086: begin
            cosine_reg0 <= 36'sb110001110001000001111101111001000010;
            sine_reg0   <= 36'sb100011010101110000100110000010001011;
        end
        11087: begin
            cosine_reg0 <= 36'sb110001110001101110111111011000100101;
            sine_reg0   <= 36'sb100011010101011010001111101000111011;
        end
        11088: begin
            cosine_reg0 <= 36'sb110001110010011100000001011011001110;
            sine_reg0   <= 36'sb100011010101000011111010010110011001;
        end
        11089: begin
            cosine_reg0 <= 36'sb110001110011001001000100000000111011;
            sine_reg0   <= 36'sb100011010100101101100110001010100110;
        end
        11090: begin
            cosine_reg0 <= 36'sb110001110011110110000111001001101010;
            sine_reg0   <= 36'sb100011010100010111010011000101100100;
        end
        11091: begin
            cosine_reg0 <= 36'sb110001110100100011001010110101011011;
            sine_reg0   <= 36'sb100011010100000001000001000111010100;
        end
        11092: begin
            cosine_reg0 <= 36'sb110001110101010000001111000100001010;
            sine_reg0   <= 36'sb100011010011101010110000001111110101;
        end
        11093: begin
            cosine_reg0 <= 36'sb110001110101111101010011110101110111;
            sine_reg0   <= 36'sb100011010011010100100000011111001001;
        end
        11094: begin
            cosine_reg0 <= 36'sb110001110110101010011001001010011111;
            sine_reg0   <= 36'sb100011010010111110010001110101010001;
        end
        11095: begin
            cosine_reg0 <= 36'sb110001110111010111011111000010000001;
            sine_reg0   <= 36'sb100011010010101000000100010010001110;
        end
        11096: begin
            cosine_reg0 <= 36'sb110001111000000100100101011100011100;
            sine_reg0   <= 36'sb100011010010010001110111110110000001;
        end
        11097: begin
            cosine_reg0 <= 36'sb110001111000110001101100011001101100;
            sine_reg0   <= 36'sb100011010001111011101100100000101001;
        end
        11098: begin
            cosine_reg0 <= 36'sb110001111001011110110011111001110001;
            sine_reg0   <= 36'sb100011010001100101100010010010001001;
        end
        11099: begin
            cosine_reg0 <= 36'sb110001111010001011111011111100101010;
            sine_reg0   <= 36'sb100011010001001111011001001010100010;
        end
        11100: begin
            cosine_reg0 <= 36'sb110001111010111001000100100010010011;
            sine_reg0   <= 36'sb100011010000111001010001001001110011;
        end
        11101: begin
            cosine_reg0 <= 36'sb110001111011100110001101101010101011;
            sine_reg0   <= 36'sb100011010000100011001010001111111110;
        end
        11102: begin
            cosine_reg0 <= 36'sb110001111100010011010111010101110010;
            sine_reg0   <= 36'sb100011010000001101000100011101000011;
        end
        11103: begin
            cosine_reg0 <= 36'sb110001111101000000100001100011100100;
            sine_reg0   <= 36'sb100011001111110110111111110001000100;
        end
        11104: begin
            cosine_reg0 <= 36'sb110001111101101101101100010100000000;
            sine_reg0   <= 36'sb100011001111100000111100001100000010;
        end
        11105: begin
            cosine_reg0 <= 36'sb110001111110011010110111100111000101;
            sine_reg0   <= 36'sb100011001111001010111001101101111100;
        end
        11106: begin
            cosine_reg0 <= 36'sb110001111111001000000011011100110001;
            sine_reg0   <= 36'sb100011001110110100111000010110110101;
        end
        11107: begin
            cosine_reg0 <= 36'sb110001111111110101001111110101000001;
            sine_reg0   <= 36'sb100011001110011110111000000110101101;
        end
        11108: begin
            cosine_reg0 <= 36'sb110010000000100010011100101111110101;
            sine_reg0   <= 36'sb100011001110001000111000111101100100;
        end
        11109: begin
            cosine_reg0 <= 36'sb110010000001001111101010001101001010;
            sine_reg0   <= 36'sb100011001101110010111010111011011100;
        end
        11110: begin
            cosine_reg0 <= 36'sb110010000001111100111000001100111111;
            sine_reg0   <= 36'sb100011001101011100111110000000010110;
        end
        11111: begin
            cosine_reg0 <= 36'sb110010000010101010000110101111010001;
            sine_reg0   <= 36'sb100011001101000111000010001100010001;
        end
        11112: begin
            cosine_reg0 <= 36'sb110010000011010111010101110100000000;
            sine_reg0   <= 36'sb100011001100110001000111011111010000;
        end
        11113: begin
            cosine_reg0 <= 36'sb110010000100000100100101011011001010;
            sine_reg0   <= 36'sb100011001100011011001101111001010011;
        end
        11114: begin
            cosine_reg0 <= 36'sb110010000100110001110101100100101100;
            sine_reg0   <= 36'sb100011001100000101010101011010011011;
        end
        11115: begin
            cosine_reg0 <= 36'sb110010000101011111000110010000100110;
            sine_reg0   <= 36'sb100011001011101111011110000010101000;
        end
        11116: begin
            cosine_reg0 <= 36'sb110010000110001100010111011110110100;
            sine_reg0   <= 36'sb100011001011011001100111110001111100;
        end
        11117: begin
            cosine_reg0 <= 36'sb110010000110111001101001001111010110;
            sine_reg0   <= 36'sb100011001011000011110010101000011000;
        end
        11118: begin
            cosine_reg0 <= 36'sb110010000111100110111011100010001010;
            sine_reg0   <= 36'sb100011001010101101111110100101111011;
        end
        11119: begin
            cosine_reg0 <= 36'sb110010001000010100001110010111001110;
            sine_reg0   <= 36'sb100011001010011000001011101010101000;
        end
        11120: begin
            cosine_reg0 <= 36'sb110010001001000001100001101110100000;
            sine_reg0   <= 36'sb100011001010000010011001110110011110;
        end
        11121: begin
            cosine_reg0 <= 36'sb110010001001101110110101100111111110;
            sine_reg0   <= 36'sb100011001001101100101001001001011111;
        end
        11122: begin
            cosine_reg0 <= 36'sb110010001010011100001010000011101000;
            sine_reg0   <= 36'sb100011001001010110111001100011101100;
        end
        11123: begin
            cosine_reg0 <= 36'sb110010001011001001011111000001011010;
            sine_reg0   <= 36'sb100011001001000001001011000101000101;
        end
        11124: begin
            cosine_reg0 <= 36'sb110010001011110110110100100001010100;
            sine_reg0   <= 36'sb100011001000101011011101101101101100;
        end
        11125: begin
            cosine_reg0 <= 36'sb110010001100100100001010100011010011;
            sine_reg0   <= 36'sb100011001000010101110001011101100000;
        end
        11126: begin
            cosine_reg0 <= 36'sb110010001101010001100001000111010110;
            sine_reg0   <= 36'sb100011001000000000000110010100100100;
        end
        11127: begin
            cosine_reg0 <= 36'sb110010001101111110111000001101011011;
            sine_reg0   <= 36'sb100011000111101010011100010010110111;
        end
        11128: begin
            cosine_reg0 <= 36'sb110010001110101100001111110101100001;
            sine_reg0   <= 36'sb100011000111010100110011011000011010;
        end
        11129: begin
            cosine_reg0 <= 36'sb110010001111011001100111111111100101;
            sine_reg0   <= 36'sb100011000110111111001011100101010000;
        end
        11130: begin
            cosine_reg0 <= 36'sb110010010000000111000000101011100101;
            sine_reg0   <= 36'sb100011000110101001100100111001010111;
        end
        11131: begin
            cosine_reg0 <= 36'sb110010010000110100011001111001100001;
            sine_reg0   <= 36'sb100011000110010011111111010100110010;
        end
        11132: begin
            cosine_reg0 <= 36'sb110010010001100001110011101001010110;
            sine_reg0   <= 36'sb100011000101111110011010110111100000;
        end
        11133: begin
            cosine_reg0 <= 36'sb110010010010001111001101111011000011;
            sine_reg0   <= 36'sb100011000101101000110111100001100011;
        end
        11134: begin
            cosine_reg0 <= 36'sb110010010010111100101000101110100101;
            sine_reg0   <= 36'sb100011000101010011010101010010111100;
        end
        11135: begin
            cosine_reg0 <= 36'sb110010010011101010000100000011111100;
            sine_reg0   <= 36'sb100011000100111101110100001011101011;
        end
        11136: begin
            cosine_reg0 <= 36'sb110010010100010111011111111011000100;
            sine_reg0   <= 36'sb100011000100101000010100001011110010;
        end
        11137: begin
            cosine_reg0 <= 36'sb110010010101000100111100010011111101;
            sine_reg0   <= 36'sb100011000100010010110101010011010000;
        end
        11138: begin
            cosine_reg0 <= 36'sb110010010101110010011001001110100110;
            sine_reg0   <= 36'sb100011000011111101010111100010001000;
        end
        11139: begin
            cosine_reg0 <= 36'sb110010010110011111110110101010111011;
            sine_reg0   <= 36'sb100011000011100111111010111000011001;
        end
        11140: begin
            cosine_reg0 <= 36'sb110010010111001101010100101000111011;
            sine_reg0   <= 36'sb100011000011010010011111010110000100;
        end
        11141: begin
            cosine_reg0 <= 36'sb110010010111111010110011001000100101;
            sine_reg0   <= 36'sb100011000010111101000100111011001100;
        end
        11142: begin
            cosine_reg0 <= 36'sb110010011000101000010010001001110110;
            sine_reg0   <= 36'sb100011000010100111101011100111101111;
        end
        11143: begin
            cosine_reg0 <= 36'sb110010011001010101110001101100101110;
            sine_reg0   <= 36'sb100011000010010010010011011011101111;
        end
        11144: begin
            cosine_reg0 <= 36'sb110010011010000011010001110001001010;
            sine_reg0   <= 36'sb100011000001111100111100010111001101;
        end
        11145: begin
            cosine_reg0 <= 36'sb110010011010110000110010010111001000;
            sine_reg0   <= 36'sb100011000001100111100110011010001010;
        end
        11146: begin
            cosine_reg0 <= 36'sb110010011011011110010011011110101000;
            sine_reg0   <= 36'sb100011000001010010010001100100100111;
        end
        11147: begin
            cosine_reg0 <= 36'sb110010011100001011110101000111100110;
            sine_reg0   <= 36'sb100011000000111100111101110110100011;
        end
        11148: begin
            cosine_reg0 <= 36'sb110010011100111001010111010010000001;
            sine_reg0   <= 36'sb100011000000100111101011010000000001;
        end
        11149: begin
            cosine_reg0 <= 36'sb110010011101100110111001111101111000;
            sine_reg0   <= 36'sb100011000000010010011001110001000001;
        end
        11150: begin
            cosine_reg0 <= 36'sb110010011110010100011101001011001001;
            sine_reg0   <= 36'sb100010111111111101001001011001100011;
        end
        11151: begin
            cosine_reg0 <= 36'sb110010011111000010000000111001110010;
            sine_reg0   <= 36'sb100010111111100111111010001001101010;
        end
        11152: begin
            cosine_reg0 <= 36'sb110010011111101111100101001001110001;
            sine_reg0   <= 36'sb100010111111010010101100000001010100;
        end
        11153: begin
            cosine_reg0 <= 36'sb110010100000011101001001111011000100;
            sine_reg0   <= 36'sb100010111110111101011111000000100100;
        end
        11154: begin
            cosine_reg0 <= 36'sb110010100001001010101111001101101010;
            sine_reg0   <= 36'sb100010111110101000010011000111011010;
        end
        11155: begin
            cosine_reg0 <= 36'sb110010100001111000010101000001100001;
            sine_reg0   <= 36'sb100010111110010011001000010101110111;
        end
        11156: begin
            cosine_reg0 <= 36'sb110010100010100101111011010110100111;
            sine_reg0   <= 36'sb100010111101111101111110101011111011;
        end
        11157: begin
            cosine_reg0 <= 36'sb110010100011010011100010001100111011;
            sine_reg0   <= 36'sb100010111101101000110110001001101000;
        end
        11158: begin
            cosine_reg0 <= 36'sb110010100100000001001001100100011010;
            sine_reg0   <= 36'sb100010111101010011101110101110111111;
        end
        11159: begin
            cosine_reg0 <= 36'sb110010100100101110110001011101000011;
            sine_reg0   <= 36'sb100010111100111110101000011011111111;
        end
        11160: begin
            cosine_reg0 <= 36'sb110010100101011100011001110110110101;
            sine_reg0   <= 36'sb100010111100101001100011010000101010;
        end
        11161: begin
            cosine_reg0 <= 36'sb110010100110001010000010110001101101;
            sine_reg0   <= 36'sb100010111100010100011111001101000010;
        end
        11162: begin
            cosine_reg0 <= 36'sb110010100110110111101100001101101001;
            sine_reg0   <= 36'sb100010111011111111011100010001000101;
        end
        11163: begin
            cosine_reg0 <= 36'sb110010100111100101010110001010101000;
            sine_reg0   <= 36'sb100010111011101010011010011100110111;
        end
        11164: begin
            cosine_reg0 <= 36'sb110010101000010011000000101000101001;
            sine_reg0   <= 36'sb100010111011010101011001110000010110;
        end
        11165: begin
            cosine_reg0 <= 36'sb110010101001000000101011100111101001;
            sine_reg0   <= 36'sb100010111011000000011010001011100100;
        end
        11166: begin
            cosine_reg0 <= 36'sb110010101001101110010111000111100110;
            sine_reg0   <= 36'sb100010111010101011011011101110100010;
        end
        11167: begin
            cosine_reg0 <= 36'sb110010101010011100000011001000011111;
            sine_reg0   <= 36'sb100010111010010110011110011001010001;
        end
        11168: begin
            cosine_reg0 <= 36'sb110010101011001001101111101010010011;
            sine_reg0   <= 36'sb100010111010000001100010001011110001;
        end
        11169: begin
            cosine_reg0 <= 36'sb110010101011110111011100101100111110;
            sine_reg0   <= 36'sb100010111001101100100111000110000100;
        end
        11170: begin
            cosine_reg0 <= 36'sb110010101100100101001010010000100001;
            sine_reg0   <= 36'sb100010111001010111101101001000001001;
        end
        11171: begin
            cosine_reg0 <= 36'sb110010101101010010111000010100111000;
            sine_reg0   <= 36'sb100010111001000010110100010010000011;
        end
        11172: begin
            cosine_reg0 <= 36'sb110010101110000000100110111010000010;
            sine_reg0   <= 36'sb100010111000101101111100100011110001;
        end
        11173: begin
            cosine_reg0 <= 36'sb110010101110101110010101111111111101;
            sine_reg0   <= 36'sb100010111000011001000101111101010100;
        end
        11174: begin
            cosine_reg0 <= 36'sb110010101111011100000101100110101000;
            sine_reg0   <= 36'sb100010111000000100010000011110101110;
        end
        11175: begin
            cosine_reg0 <= 36'sb110010110000001001110101101110000000;
            sine_reg0   <= 36'sb100010110111101111011100000111111111;
        end
        11176: begin
            cosine_reg0 <= 36'sb110010110000110111100110010110000101;
            sine_reg0   <= 36'sb100010110111011010101000111001000111;
        end
        11177: begin
            cosine_reg0 <= 36'sb110010110001100101010111011110110100;
            sine_reg0   <= 36'sb100010110111000101110110110010001001;
        end
        11178: begin
            cosine_reg0 <= 36'sb110010110010010011001001001000001011;
            sine_reg0   <= 36'sb100010110110110001000101110011000100;
        end
        11179: begin
            cosine_reg0 <= 36'sb110010110011000000111011010010001001;
            sine_reg0   <= 36'sb100010110110011100010101111011111001;
        end
        11180: begin
            cosine_reg0 <= 36'sb110010110011101110101101111100101100;
            sine_reg0   <= 36'sb100010110110000111100111001100101001;
        end
        11181: begin
            cosine_reg0 <= 36'sb110010110100011100100001000111110001;
            sine_reg0   <= 36'sb100010110101110010111001100101010101;
        end
        11182: begin
            cosine_reg0 <= 36'sb110010110101001010010100110011011001;
            sine_reg0   <= 36'sb100010110101011110001101000101111110;
        end
        11183: begin
            cosine_reg0 <= 36'sb110010110101111000001000111111100000;
            sine_reg0   <= 36'sb100010110101001001100001101110100100;
        end
        11184: begin
            cosine_reg0 <= 36'sb110010110110100101111101101100000101;
            sine_reg0   <= 36'sb100010110100110100110111011111001001;
        end
        11185: begin
            cosine_reg0 <= 36'sb110010110111010011110010111001000101;
            sine_reg0   <= 36'sb100010110100100000001110010111101100;
        end
        11186: begin
            cosine_reg0 <= 36'sb110010111000000001101000100110100001;
            sine_reg0   <= 36'sb100010110100001011100110011000010000;
        end
        11187: begin
            cosine_reg0 <= 36'sb110010111000101111011110110100010100;
            sine_reg0   <= 36'sb100010110011110110111111100000110100;
        end
        11188: begin
            cosine_reg0 <= 36'sb110010111001011101010101100010011111;
            sine_reg0   <= 36'sb100010110011100010011001110001011001;
        end
        11189: begin
            cosine_reg0 <= 36'sb110010111010001011001100110000111111;
            sine_reg0   <= 36'sb100010110011001101110101001010000001;
        end
        11190: begin
            cosine_reg0 <= 36'sb110010111010111001000100011111110001;
            sine_reg0   <= 36'sb100010110010111001010001101010101100;
        end
        11191: begin
            cosine_reg0 <= 36'sb110010111011100110111100101110110110;
            sine_reg0   <= 36'sb100010110010100100101111010011011011;
        end
        11192: begin
            cosine_reg0 <= 36'sb110010111100010100110101011110001010;
            sine_reg0   <= 36'sb100010110010010000001110000100001110;
        end
        11193: begin
            cosine_reg0 <= 36'sb110010111101000010101110101101101100;
            sine_reg0   <= 36'sb100010110001111011101101111101000111;
        end
        11194: begin
            cosine_reg0 <= 36'sb110010111101110000101000011101011010;
            sine_reg0   <= 36'sb100010110001100111001110111110000110;
        end
        11195: begin
            cosine_reg0 <= 36'sb110010111110011110100010101101010010;
            sine_reg0   <= 36'sb100010110001010010110001000111001011;
        end
        11196: begin
            cosine_reg0 <= 36'sb110010111111001100011101011101010100;
            sine_reg0   <= 36'sb100010110000111110010100011000011001;
        end
        11197: begin
            cosine_reg0 <= 36'sb110010111111111010011000101101011100;
            sine_reg0   <= 36'sb100010110000101001111000110001101111;
        end
        11198: begin
            cosine_reg0 <= 36'sb110011000000101000010100011101101001;
            sine_reg0   <= 36'sb100010110000010101011110010011001111;
        end
        11199: begin
            cosine_reg0 <= 36'sb110011000001010110010000101101111001;
            sine_reg0   <= 36'sb100010110000000001000100111100111001;
        end
        11200: begin
            cosine_reg0 <= 36'sb110011000010000100001101011110001011;
            sine_reg0   <= 36'sb100010101111101100101100101110101101;
        end
        11201: begin
            cosine_reg0 <= 36'sb110011000010110010001010101110011101;
            sine_reg0   <= 36'sb100010101111011000010101101000101110;
        end
        11202: begin
            cosine_reg0 <= 36'sb110011000011100000001000011110101101;
            sine_reg0   <= 36'sb100010101111000011111111101010111011;
        end
        11203: begin
            cosine_reg0 <= 36'sb110011000100001110000110101110111001;
            sine_reg0   <= 36'sb100010101110101111101010110101010101;
        end
        11204: begin
            cosine_reg0 <= 36'sb110011000100111100000101011110111111;
            sine_reg0   <= 36'sb100010101110011011010111000111111101;
        end
        11205: begin
            cosine_reg0 <= 36'sb110011000101101010000100101110111111;
            sine_reg0   <= 36'sb100010101110000111000100100010110100;
        end
        11206: begin
            cosine_reg0 <= 36'sb110011000110011000000100011110110101;
            sine_reg0   <= 36'sb100010101101110010110011000101111011;
        end
        11207: begin
            cosine_reg0 <= 36'sb110011000111000110000100101110100000;
            sine_reg0   <= 36'sb100010101101011110100010110001010010;
        end
        11208: begin
            cosine_reg0 <= 36'sb110011000111110100000101011101111111;
            sine_reg0   <= 36'sb100010101101001010010011100100111011;
        end
        11209: begin
            cosine_reg0 <= 36'sb110011001000100010000110101101001111;
            sine_reg0   <= 36'sb100010101100110110000101100000110101;
        end
        11210: begin
            cosine_reg0 <= 36'sb110011001001010000001000011100001111;
            sine_reg0   <= 36'sb100010101100100001111000100101000010;
        end
        11211: begin
            cosine_reg0 <= 36'sb110011001001111110001010101010111101;
            sine_reg0   <= 36'sb100010101100001101101100110001100011;
        end
        11212: begin
            cosine_reg0 <= 36'sb110011001010101100001101011001010111;
            sine_reg0   <= 36'sb100010101011111001100010000110011000;
        end
        11213: begin
            cosine_reg0 <= 36'sb110011001011011010010000100111011100;
            sine_reg0   <= 36'sb100010101011100101011000100011100010;
        end
        11214: begin
            cosine_reg0 <= 36'sb110011001100001000010100010101001010;
            sine_reg0   <= 36'sb100010101011010001010000001001000010;
        end
        11215: begin
            cosine_reg0 <= 36'sb110011001100110110011000100010011110;
            sine_reg0   <= 36'sb100010101010111101001000110110111001;
        end
        11216: begin
            cosine_reg0 <= 36'sb110011001101100100011101001111011000;
            sine_reg0   <= 36'sb100010101010101001000010101101000111;
        end
        11217: begin
            cosine_reg0 <= 36'sb110011001110010010100010011011110101;
            sine_reg0   <= 36'sb100010101010010100111101101011101101;
        end
        11218: begin
            cosine_reg0 <= 36'sb110011001111000000101000000111110100;
            sine_reg0   <= 36'sb100010101010000000111001110010101100;
        end
        11219: begin
            cosine_reg0 <= 36'sb110011001111101110101110010011010011;
            sine_reg0   <= 36'sb100010101001101100110111000010000101;
        end
        11220: begin
            cosine_reg0 <= 36'sb110011010000011100110100111110001111;
            sine_reg0   <= 36'sb100010101001011000110101011001111000;
        end
        11221: begin
            cosine_reg0 <= 36'sb110011010001001010111100001000101000;
            sine_reg0   <= 36'sb100010101001000100110100111010000111;
        end
        11222: begin
            cosine_reg0 <= 36'sb110011010001111001000011110010011100;
            sine_reg0   <= 36'sb100010101000110000110101100010110010;
        end
        11223: begin
            cosine_reg0 <= 36'sb110011010010100111001011111011101000;
            sine_reg0   <= 36'sb100010101000011100110111010011111010;
        end
        11224: begin
            cosine_reg0 <= 36'sb110011010011010101010100100100001011;
            sine_reg0   <= 36'sb100010101000001000111010001101011111;
        end
        11225: begin
            cosine_reg0 <= 36'sb110011010100000011011101101100000011;
            sine_reg0   <= 36'sb100010100111110100111110001111100010;
        end
        11226: begin
            cosine_reg0 <= 36'sb110011010100110001100111010011001111;
            sine_reg0   <= 36'sb100010100111100001000011011010000101;
        end
        11227: begin
            cosine_reg0 <= 36'sb110011010101011111110001011001101100;
            sine_reg0   <= 36'sb100010100111001101001001101101001000;
        end
        11228: begin
            cosine_reg0 <= 36'sb110011010110001101111011111111011001;
            sine_reg0   <= 36'sb100010100110111001010001001000101011;
        end
        11229: begin
            cosine_reg0 <= 36'sb110011010110111100000111000100010101;
            sine_reg0   <= 36'sb100010100110100101011001101100110000;
        end
        11230: begin
            cosine_reg0 <= 36'sb110011010111101010010010101000011100;
            sine_reg0   <= 36'sb100010100110010001100011011001010111;
        end
        11231: begin
            cosine_reg0 <= 36'sb110011011000011000011110101011101110;
            sine_reg0   <= 36'sb100010100101111101101110001110100001;
        end
        11232: begin
            cosine_reg0 <= 36'sb110011011001000110101011001110001001;
            sine_reg0   <= 36'sb100010100101101001111010001100001110;
        end
        11233: begin
            cosine_reg0 <= 36'sb110011011001110100111000001111101010;
            sine_reg0   <= 36'sb100010100101010110000111010010100001;
        end
        11234: begin
            cosine_reg0 <= 36'sb110011011010100011000101110000010001;
            sine_reg0   <= 36'sb100010100101000010010101100001011000;
        end
        11235: begin
            cosine_reg0 <= 36'sb110011011011010001010011101111111011;
            sine_reg0   <= 36'sb100010100100101110100100111000110110;
        end
        11236: begin
            cosine_reg0 <= 36'sb110011011011111111100010001110100111;
            sine_reg0   <= 36'sb100010100100011010110101011000111010;
        end
        11237: begin
            cosine_reg0 <= 36'sb110011011100101101110001001100010011;
            sine_reg0   <= 36'sb100010100100000111000111000001100110;
        end
        11238: begin
            cosine_reg0 <= 36'sb110011011101011100000000101000111100;
            sine_reg0   <= 36'sb100010100011110011011001110010111010;
        end
        11239: begin
            cosine_reg0 <= 36'sb110011011110001010010000100100100010;
            sine_reg0   <= 36'sb100010100011011111101101101100110111;
        end
        11240: begin
            cosine_reg0 <= 36'sb110011011110111000100000111111000010;
            sine_reg0   <= 36'sb100010100011001100000010101111011110;
        end
        11241: begin
            cosine_reg0 <= 36'sb110011011111100110110001111000011011;
            sine_reg0   <= 36'sb100010100010111000011000111010110000;
        end
        11242: begin
            cosine_reg0 <= 36'sb110011100000010101000011010000101011;
            sine_reg0   <= 36'sb100010100010100100110000001110101100;
        end
        11243: begin
            cosine_reg0 <= 36'sb110011100001000011010101000111110000;
            sine_reg0   <= 36'sb100010100010010001001000101011010101;
        end
        11244: begin
            cosine_reg0 <= 36'sb110011100001110001100111011101101001;
            sine_reg0   <= 36'sb100010100001111101100010010000101011;
        end
        11245: begin
            cosine_reg0 <= 36'sb110011100010011111111010010010010010;
            sine_reg0   <= 36'sb100010100001101001111100111110101111;
        end
        11246: begin
            cosine_reg0 <= 36'sb110011100011001110001101100101101100;
            sine_reg0   <= 36'sb100010100001010110011000110101100001;
        end
        11247: begin
            cosine_reg0 <= 36'sb110011100011111100100001010111110100;
            sine_reg0   <= 36'sb100010100001000010110101110101000010;
        end
        11248: begin
            cosine_reg0 <= 36'sb110011100100101010110101101000100111;
            sine_reg0   <= 36'sb100010100000101111010011111101010011;
        end
        11249: begin
            cosine_reg0 <= 36'sb110011100101011001001010011000000101;
            sine_reg0   <= 36'sb100010100000011011110011001110010100;
        end
        11250: begin
            cosine_reg0 <= 36'sb110011100110000111011111100110001100;
            sine_reg0   <= 36'sb100010100000001000010011101000000111;
        end
        11251: begin
            cosine_reg0 <= 36'sb110011100110110101110101010010111010;
            sine_reg0   <= 36'sb100010011111110100110101001010101100;
        end
        11252: begin
            cosine_reg0 <= 36'sb110011100111100100001011011110001100;
            sine_reg0   <= 36'sb100010011111100001010111110110000100;
        end
        11253: begin
            cosine_reg0 <= 36'sb110011101000010010100010001000000010;
            sine_reg0   <= 36'sb100010011111001101111011101010010000;
        end
        11254: begin
            cosine_reg0 <= 36'sb110011101001000000111001010000011010;
            sine_reg0   <= 36'sb100010011110111010100000100111010000;
        end
        11255: begin
            cosine_reg0 <= 36'sb110011101001101111010000110111010001;
            sine_reg0   <= 36'sb100010011110100111000110101101000101;
        end
        11256: begin
            cosine_reg0 <= 36'sb110011101010011101101000111100100110;
            sine_reg0   <= 36'sb100010011110010011101101111011110000;
        end
        11257: begin
            cosine_reg0 <= 36'sb110011101011001100000001100000010111;
            sine_reg0   <= 36'sb100010011110000000010110010011010001;
        end
        11258: begin
            cosine_reg0 <= 36'sb110011101011111010011010100010100010;
            sine_reg0   <= 36'sb100010011101101100111111110011101010;
        end
        11259: begin
            cosine_reg0 <= 36'sb110011101100101000110100000011000110;
            sine_reg0   <= 36'sb100010011101011001101010011100111011;
        end
        11260: begin
            cosine_reg0 <= 36'sb110011101101010111001110000010000001;
            sine_reg0   <= 36'sb100010011101000110010110001111000101;
        end
        11261: begin
            cosine_reg0 <= 36'sb110011101110000101101000011111010000;
            sine_reg0   <= 36'sb100010011100110011000011001010001001;
        end
        11262: begin
            cosine_reg0 <= 36'sb110011101110110100000011011010110011;
            sine_reg0   <= 36'sb100010011100011111110001001110000110;
        end
        11263: begin
            cosine_reg0 <= 36'sb110011101111100010011110110100100111;
            sine_reg0   <= 36'sb100010011100001100100000011010111111;
        end
        11264: begin
            cosine_reg0 <= 36'sb110011110000010000111010101100101011;
            sine_reg0   <= 36'sb100010011011111001010000110000110100;
        end
        11265: begin
            cosine_reg0 <= 36'sb110011110000111111010111000010111100;
            sine_reg0   <= 36'sb100010011011100110000010001111100110;
        end
        11266: begin
            cosine_reg0 <= 36'sb110011110001101101110011110111011001;
            sine_reg0   <= 36'sb100010011011010010110100110111010100;
        end
        11267: begin
            cosine_reg0 <= 36'sb110011110010011100010001001010000001;
            sine_reg0   <= 36'sb100010011010111111101000101000000001;
        end
        11268: begin
            cosine_reg0 <= 36'sb110011110011001010101110111010110001;
            sine_reg0   <= 36'sb100010011010101100011101100001101101;
        end
        11269: begin
            cosine_reg0 <= 36'sb110011110011111001001101001001101000;
            sine_reg0   <= 36'sb100010011010011001010011100100011000;
        end
        11270: begin
            cosine_reg0 <= 36'sb110011110100100111101011110110100011;
            sine_reg0   <= 36'sb100010011010000110001010110000000011;
        end
        11271: begin
            cosine_reg0 <= 36'sb110011110101010110001011000001100010;
            sine_reg0   <= 36'sb100010011001110011000011000100110000;
        end
        11272: begin
            cosine_reg0 <= 36'sb110011110110000100101010101010100010;
            sine_reg0   <= 36'sb100010011001011111111100100010011110;
        end
        11273: begin
            cosine_reg0 <= 36'sb110011110110110011001010110001100001;
            sine_reg0   <= 36'sb100010011001001100110111001001001111;
        end
        11274: begin
            cosine_reg0 <= 36'sb110011110111100001101011010110011110;
            sine_reg0   <= 36'sb100010011000111001110010111001000011;
        end
        11275: begin
            cosine_reg0 <= 36'sb110011111000010000001100011001010111;
            sine_reg0   <= 36'sb100010011000100110101111110001111011;
        end
        11276: begin
            cosine_reg0 <= 36'sb110011111000111110101101111010001010;
            sine_reg0   <= 36'sb100010011000010011101101110011110111;
        end
        11277: begin
            cosine_reg0 <= 36'sb110011111001101101001111111000110101;
            sine_reg0   <= 36'sb100010011000000000101100111110111001;
        end
        11278: begin
            cosine_reg0 <= 36'sb110011111010011011110010010101010111;
            sine_reg0   <= 36'sb100010010111101101101101010011000001;
        end
        11279: begin
            cosine_reg0 <= 36'sb110011111011001010010101001111101101;
            sine_reg0   <= 36'sb100010010111011010101110110000010001;
        end
        11280: begin
            cosine_reg0 <= 36'sb110011111011111000111000100111110111;
            sine_reg0   <= 36'sb100010010111000111110001010110100111;
        end
        11281: begin
            cosine_reg0 <= 36'sb110011111100100111011100011101110001;
            sine_reg0   <= 36'sb100010010110110100110101000110000110;
        end
        11282: begin
            cosine_reg0 <= 36'sb110011111101010110000000110001011011;
            sine_reg0   <= 36'sb100010010110100001111001111110101111;
        end
        11283: begin
            cosine_reg0 <= 36'sb110011111110000100100101100010110010;
            sine_reg0   <= 36'sb100010010110001111000000000000100001;
        end
        11284: begin
            cosine_reg0 <= 36'sb110011111110110011001010110001110101;
            sine_reg0   <= 36'sb100010010101111100000111001011011101;
        end
        11285: begin
            cosine_reg0 <= 36'sb110011111111100001110000011110100010;
            sine_reg0   <= 36'sb100010010101101001001111011111100101;
        end
        11286: begin
            cosine_reg0 <= 36'sb110100000000010000010110101000110111;
            sine_reg0   <= 36'sb100010010101010110011000111100111001;
        end
        11287: begin
            cosine_reg0 <= 36'sb110100000000111110111101010000110010;
            sine_reg0   <= 36'sb100010010101000011100011100011011001;
        end
        11288: begin
            cosine_reg0 <= 36'sb110100000001101101100100010110010010;
            sine_reg0   <= 36'sb100010010100110000101111010011000111;
        end
        11289: begin
            cosine_reg0 <= 36'sb110100000010011100001011111001010101;
            sine_reg0   <= 36'sb100010010100011101111100001100000011;
        end
        11290: begin
            cosine_reg0 <= 36'sb110100000011001010110011111001111000;
            sine_reg0   <= 36'sb100010010100001011001010001110001111;
        end
        11291: begin
            cosine_reg0 <= 36'sb110100000011111001011100010111111011;
            sine_reg0   <= 36'sb100010010011111000011001011001101001;
        end
        11292: begin
            cosine_reg0 <= 36'sb110100000100101000000101010011011011;
            sine_reg0   <= 36'sb100010010011100101101001101110010100;
        end
        11293: begin
            cosine_reg0 <= 36'sb110100000101010110101110101100010111;
            sine_reg0   <= 36'sb100010010011010010111011001100010001;
        end
        11294: begin
            cosine_reg0 <= 36'sb110100000110000101011000100010101100;
            sine_reg0   <= 36'sb100010010011000000001101110011011111;
        end
        11295: begin
            cosine_reg0 <= 36'sb110100000110110100000010110110011001;
            sine_reg0   <= 36'sb100010010010101101100001100011111111;
        end
        11296: begin
            cosine_reg0 <= 36'sb110100000111100010101101100111011101;
            sine_reg0   <= 36'sb100010010010011010110110011101110011;
        end
        11297: begin
            cosine_reg0 <= 36'sb110100001000010001011000110101110100;
            sine_reg0   <= 36'sb100010010010001000001100100000111010;
        end
        11298: begin
            cosine_reg0 <= 36'sb110100001001000000000100100001011111;
            sine_reg0   <= 36'sb100010010001110101100011101101010111;
        end
        11299: begin
            cosine_reg0 <= 36'sb110100001001101110110000101010011010;
            sine_reg0   <= 36'sb100010010001100010111100000011001001;
        end
        11300: begin
            cosine_reg0 <= 36'sb110100001010011101011101010000100100;
            sine_reg0   <= 36'sb100010010001010000010101100010010000;
        end
        11301: begin
            cosine_reg0 <= 36'sb110100001011001100001010010011111011;
            sine_reg0   <= 36'sb100010010000111101110000001010101111;
        end
        11302: begin
            cosine_reg0 <= 36'sb110100001011111010110111110100011110;
            sine_reg0   <= 36'sb100010010000101011001011111100100101;
        end
        11303: begin
            cosine_reg0 <= 36'sb110100001100101001100101110010001010;
            sine_reg0   <= 36'sb100010010000011000101000110111110100;
        end
        11304: begin
            cosine_reg0 <= 36'sb110100001101011000010100001100111110;
            sine_reg0   <= 36'sb100010010000000110000110111100011100;
        end
        11305: begin
            cosine_reg0 <= 36'sb110100001110000111000011000100111000;
            sine_reg0   <= 36'sb100010001111110011100110001010011101;
        end
        11306: begin
            cosine_reg0 <= 36'sb110100001110110101110010011001110110;
            sine_reg0   <= 36'sb100010001111100001000110100001111000;
        end
        11307: begin
            cosine_reg0 <= 36'sb110100001111100100100010001011110110;
            sine_reg0   <= 36'sb100010001111001110101000000010101111;
        end
        11308: begin
            cosine_reg0 <= 36'sb110100010000010011010010011010110111;
            sine_reg0   <= 36'sb100010001110111100001010101101000010;
        end
        11309: begin
            cosine_reg0 <= 36'sb110100010001000010000011000110110111;
            sine_reg0   <= 36'sb100010001110101001101110100000110001;
        end
        11310: begin
            cosine_reg0 <= 36'sb110100010001110000110100001111110011;
            sine_reg0   <= 36'sb100010001110010111010011011101111101;
        end
        11311: begin
            cosine_reg0 <= 36'sb110100010010011111100101110101101011;
            sine_reg0   <= 36'sb100010001110000100111001100100101000;
        end
        11312: begin
            cosine_reg0 <= 36'sb110100010011001110010111111000011100;
            sine_reg0   <= 36'sb100010001101110010100000110100110001;
        end
        11313: begin
            cosine_reg0 <= 36'sb110100010011111101001010011000000100;
            sine_reg0   <= 36'sb100010001101100000001001001110011001;
        end
        11314: begin
            cosine_reg0 <= 36'sb110100010100101011111101010100100011;
            sine_reg0   <= 36'sb100010001101001101110010110001100010;
        end
        11315: begin
            cosine_reg0 <= 36'sb110100010101011010110000101101110101;
            sine_reg0   <= 36'sb100010001100111011011101011110001011;
        end
        11316: begin
            cosine_reg0 <= 36'sb110100010110001001100100100011111001;
            sine_reg0   <= 36'sb100010001100101001001001010100010110;
        end
        11317: begin
            cosine_reg0 <= 36'sb110100010110111000011000110110101110;
            sine_reg0   <= 36'sb100010001100010110110110010100000011;
        end
        11318: begin
            cosine_reg0 <= 36'sb110100010111100111001101100110010001;
            sine_reg0   <= 36'sb100010001100000100100100011101010011;
        end
        11319: begin
            cosine_reg0 <= 36'sb110100011000010110000010110010100001;
            sine_reg0   <= 36'sb100010001011110010010011110000000110;
        end
        11320: begin
            cosine_reg0 <= 36'sb110100011001000100111000011011011100;
            sine_reg0   <= 36'sb100010001011100000000100001100011110;
        end
        11321: begin
            cosine_reg0 <= 36'sb110100011001110011101110100000111111;
            sine_reg0   <= 36'sb100010001011001101110101110010011011;
        end
        11322: begin
            cosine_reg0 <= 36'sb110100011010100010100101000011001011;
            sine_reg0   <= 36'sb100010001010111011101000100001111110;
        end
        11323: begin
            cosine_reg0 <= 36'sb110100011011010001011100000001111011;
            sine_reg0   <= 36'sb100010001010101001011100011011000111;
        end
        11324: begin
            cosine_reg0 <= 36'sb110100011100000000010011011101001111;
            sine_reg0   <= 36'sb100010001010010111010001011101110111;
        end
        11325: begin
            cosine_reg0 <= 36'sb110100011100101111001011010101000110;
            sine_reg0   <= 36'sb100010001010000101000111101010001111;
        end
        11326: begin
            cosine_reg0 <= 36'sb110100011101011110000011101001011100;
            sine_reg0   <= 36'sb100010001001110010111111000000010000;
        end
        11327: begin
            cosine_reg0 <= 36'sb110100011110001100111100011010010000;
            sine_reg0   <= 36'sb100010001001100000110111011111111010;
        end
        11328: begin
            cosine_reg0 <= 36'sb110100011110111011110101100111100001;
            sine_reg0   <= 36'sb100010001001001110110001001001001110;
        end
        11329: begin
            cosine_reg0 <= 36'sb110100011111101010101111010001001101;
            sine_reg0   <= 36'sb100010001000111100101011111100001100;
        end
        11330: begin
            cosine_reg0 <= 36'sb110100100000011001101001010111010001;
            sine_reg0   <= 36'sb100010001000101010100111111000110110;
        end
        11331: begin
            cosine_reg0 <= 36'sb110100100001001000100011111001101100;
            sine_reg0   <= 36'sb100010001000011000100100111111001100;
        end
        11332: begin
            cosine_reg0 <= 36'sb110100100001110111011110111000011101;
            sine_reg0   <= 36'sb100010001000000110100011001111001110;
        end
        11333: begin
            cosine_reg0 <= 36'sb110100100010100110011010010011100001;
            sine_reg0   <= 36'sb100010000111110100100010101000111110;
        end
        11334: begin
            cosine_reg0 <= 36'sb110100100011010101010110001010110110;
            sine_reg0   <= 36'sb100010000111100010100011001100011100;
        end
        11335: begin
            cosine_reg0 <= 36'sb110100100100000100010010011110011100;
            sine_reg0   <= 36'sb100010000111010000100100111001101001;
        end
        11336: begin
            cosine_reg0 <= 36'sb110100100100110011001111001110001111;
            sine_reg0   <= 36'sb100010000110111110100111110000100110;
        end
        11337: begin
            cosine_reg0 <= 36'sb110100100101100010001100011010001111;
            sine_reg0   <= 36'sb100010000110101100101011110001010010;
        end
        11338: begin
            cosine_reg0 <= 36'sb110100100110010001001010000010011000;
            sine_reg0   <= 36'sb100010000110011010110000111011110000;
        end
        11339: begin
            cosine_reg0 <= 36'sb110100100111000000001000000110101011;
            sine_reg0   <= 36'sb100010000110001000110111001111111111;
        end
        11340: begin
            cosine_reg0 <= 36'sb110100100111101111000110100111000100;
            sine_reg0   <= 36'sb100010000101110110111110101110000000;
        end
        11341: begin
            cosine_reg0 <= 36'sb110100101000011110000101100011100010;
            sine_reg0   <= 36'sb100010000101100101000111010101110100;
        end
        11342: begin
            cosine_reg0 <= 36'sb110100101001001101000100111100000011;
            sine_reg0   <= 36'sb100010000101010011010001000111011100;
        end
        11343: begin
            cosine_reg0 <= 36'sb110100101001111100000100110000100110;
            sine_reg0   <= 36'sb100010000101000001011100000010111000;
        end
        11344: begin
            cosine_reg0 <= 36'sb110100101010101011000101000001000111;
            sine_reg0   <= 36'sb100010000100101111101000001000001001;
        end
        11345: begin
            cosine_reg0 <= 36'sb110100101011011010000101101101100111;
            sine_reg0   <= 36'sb100010000100011101110101010111010000;
        end
        11346: begin
            cosine_reg0 <= 36'sb110100101100001001000110110110000010;
            sine_reg0   <= 36'sb100010000100001100000011110000001110;
        end
        11347: begin
            cosine_reg0 <= 36'sb110100101100111000001000011010011000;
            sine_reg0   <= 36'sb100010000011111010010011010011000010;
        end
        11348: begin
            cosine_reg0 <= 36'sb110100101101100111001010011010100110;
            sine_reg0   <= 36'sb100010000011101000100011111111101110;
        end
        11349: begin
            cosine_reg0 <= 36'sb110100101110010110001100110110101010;
            sine_reg0   <= 36'sb100010000011010110110101110110010011;
        end
        11350: begin
            cosine_reg0 <= 36'sb110100101111000101001111101110100011;
            sine_reg0   <= 36'sb100010000011000101001000110110110000;
        end
        11351: begin
            cosine_reg0 <= 36'sb110100101111110100010011000010001110;
            sine_reg0   <= 36'sb100010000010110011011101000001001000;
        end
        11352: begin
            cosine_reg0 <= 36'sb110100110000100011010110110001101011;
            sine_reg0   <= 36'sb100010000010100001110010010101011010;
        end
        11353: begin
            cosine_reg0 <= 36'sb110100110001010010011010111100110110;
            sine_reg0   <= 36'sb100010000010010000001000110011100111;
        end
        11354: begin
            cosine_reg0 <= 36'sb110100110010000001011111100011101111;
            sine_reg0   <= 36'sb100010000001111110100000011011110000;
        end
        11355: begin
            cosine_reg0 <= 36'sb110100110010110000100100100110010100;
            sine_reg0   <= 36'sb100010000001101100111001001101110110;
        end
        11356: begin
            cosine_reg0 <= 36'sb110100110011011111101010000100100010;
            sine_reg0   <= 36'sb100010000001011011010011001001111001;
        end
        11357: begin
            cosine_reg0 <= 36'sb110100110100001110101111111110011001;
            sine_reg0   <= 36'sb100010000001001001101110001111111001;
        end
        11358: begin
            cosine_reg0 <= 36'sb110100110100111101110110010011110101;
            sine_reg0   <= 36'sb100010000000111000001010011111111001;
        end
        11359: begin
            cosine_reg0 <= 36'sb110100110101101100111101000100110101;
            sine_reg0   <= 36'sb100010000000100110100111111001110111;
        end
        11360: begin
            cosine_reg0 <= 36'sb110100110110011100000100010001011000;
            sine_reg0   <= 36'sb100010000000010101000110011101110110;
        end
        11361: begin
            cosine_reg0 <= 36'sb110100110111001011001011111001011100;
            sine_reg0   <= 36'sb100010000000000011100110001011110101;
        end
        11362: begin
            cosine_reg0 <= 36'sb110100110111111010010011111100111111;
            sine_reg0   <= 36'sb100001111111110010000111000011110101;
        end
        11363: begin
            cosine_reg0 <= 36'sb110100111000101001011100011011111110;
            sine_reg0   <= 36'sb100001111111100000101001000101110111;
        end
        11364: begin
            cosine_reg0 <= 36'sb110100111001011000100101010110011001;
            sine_reg0   <= 36'sb100001111111001111001100010001111100;
        end
        11365: begin
            cosine_reg0 <= 36'sb110100111010000111101110101100001101;
            sine_reg0   <= 36'sb100001111110111101110000101000000100;
        end
        11366: begin
            cosine_reg0 <= 36'sb110100111010110110111000011101011001;
            sine_reg0   <= 36'sb100001111110101100010110001000010000;
        end
        11367: begin
            cosine_reg0 <= 36'sb110100111011100110000010101001111010;
            sine_reg0   <= 36'sb100001111110011010111100110010100001;
        end
        11368: begin
            cosine_reg0 <= 36'sb110100111100010101001101010001101111;
            sine_reg0   <= 36'sb100001111110001001100100100110110111;
        end
        11369: begin
            cosine_reg0 <= 36'sb110100111101000100011000010100110111;
            sine_reg0   <= 36'sb100001111101111000001101100101010011;
        end
        11370: begin
            cosine_reg0 <= 36'sb110100111101110011100011110011001110;
            sine_reg0   <= 36'sb100001111101100110110111101101110110;
        end
        11371: begin
            cosine_reg0 <= 36'sb110100111110100010101111101100110100;
            sine_reg0   <= 36'sb100001111101010101100011000000100000;
        end
        11372: begin
            cosine_reg0 <= 36'sb110100111111010001111100000001100111;
            sine_reg0   <= 36'sb100001111101000100001111011101010010;
        end
        11373: begin
            cosine_reg0 <= 36'sb110101000000000001001000110001100101;
            sine_reg0   <= 36'sb100001111100110010111101000100001100;
        end
        11374: begin
            cosine_reg0 <= 36'sb110101000000110000010101111100101100;
            sine_reg0   <= 36'sb100001111100100001101011110101010000;
        end
        11375: begin
            cosine_reg0 <= 36'sb110101000001011111100011100010111001;
            sine_reg0   <= 36'sb100001111100010000011011110000011110;
        end
        11376: begin
            cosine_reg0 <= 36'sb110101000010001110110001100100001101;
            sine_reg0   <= 36'sb100001111011111111001100110101110111;
        end
        11377: begin
            cosine_reg0 <= 36'sb110101000010111110000000000000100011;
            sine_reg0   <= 36'sb100001111011101101111111000101011010;
        end
        11378: begin
            cosine_reg0 <= 36'sb110101000011101101001110110111111100;
            sine_reg0   <= 36'sb100001111011011100110010011111001010;
        end
        11379: begin
            cosine_reg0 <= 36'sb110101000100011100011110001010010100;
            sine_reg0   <= 36'sb100001111011001011100111000011000111;
        end
        11380: begin
            cosine_reg0 <= 36'sb110101000101001011101101110111101010;
            sine_reg0   <= 36'sb100001111010111010011100110001010001;
        end
        11381: begin
            cosine_reg0 <= 36'sb110101000101111010111101111111111101;
            sine_reg0   <= 36'sb100001111010101001010011101001101000;
        end
        11382: begin
            cosine_reg0 <= 36'sb110101000110101010001110100011001010;
            sine_reg0   <= 36'sb100001111010011000001011101100001111;
        end
        11383: begin
            cosine_reg0 <= 36'sb110101000111011001011111100001010000;
            sine_reg0   <= 36'sb100001111010000111000100111001000100;
        end
        11384: begin
            cosine_reg0 <= 36'sb110101001000001000110000111010001101;
            sine_reg0   <= 36'sb100001111001110101111111010000001010;
        end
        11385: begin
            cosine_reg0 <= 36'sb110101001000111000000010101101111110;
            sine_reg0   <= 36'sb100001111001100100111010110001100000;
        end
        11386: begin
            cosine_reg0 <= 36'sb110101001001100111010100111100100011;
            sine_reg0   <= 36'sb100001111001010011110111011101000111;
        end
        11387: begin
            cosine_reg0 <= 36'sb110101001010010110100111100101111001;
            sine_reg0   <= 36'sb100001111001000010110101010011000001;
        end
        11388: begin
            cosine_reg0 <= 36'sb110101001011000101111010101001111110;
            sine_reg0   <= 36'sb100001111000110001110100010011001101;
        end
        11389: begin
            cosine_reg0 <= 36'sb110101001011110101001110001000110010;
            sine_reg0   <= 36'sb100001111000100000110100011101101100;
        end
        11390: begin
            cosine_reg0 <= 36'sb110101001100100100100010000010010001;
            sine_reg0   <= 36'sb100001111000001111110101110010011111;
        end
        11391: begin
            cosine_reg0 <= 36'sb110101001101010011110110010110011010;
            sine_reg0   <= 36'sb100001110111111110111000010001100111;
        end
        11392: begin
            cosine_reg0 <= 36'sb110101001110000011001011000101001011;
            sine_reg0   <= 36'sb100001110111101101111011111011000011;
        end
        11393: begin
            cosine_reg0 <= 36'sb110101001110110010100000001110100011;
            sine_reg0   <= 36'sb100001110111011101000000101110110110;
        end
        11394: begin
            cosine_reg0 <= 36'sb110101001111100001110101110010011111;
            sine_reg0   <= 36'sb100001110111001100000110101100111111;
        end
        11395: begin
            cosine_reg0 <= 36'sb110101010000010001001011110000111110;
            sine_reg0   <= 36'sb100001110110111011001101110101011111;
        end
        11396: begin
            cosine_reg0 <= 36'sb110101010001000000100010001001111110;
            sine_reg0   <= 36'sb100001110110101010010110001000010111;
        end
        11397: begin
            cosine_reg0 <= 36'sb110101010001101111111000111101011101;
            sine_reg0   <= 36'sb100001110110011001011111100101101000;
        end
        11398: begin
            cosine_reg0 <= 36'sb110101010010011111010000001011011001;
            sine_reg0   <= 36'sb100001110110001000101010001101010010;
        end
        11399: begin
            cosine_reg0 <= 36'sb110101010011001110100111110011110001;
            sine_reg0   <= 36'sb100001110101110111110101111111010101;
        end
        11400: begin
            cosine_reg0 <= 36'sb110101010011111101111111110110100010;
            sine_reg0   <= 36'sb100001110101100111000010111011110011;
        end
        11401: begin
            cosine_reg0 <= 36'sb110101010100101101011000010011101011;
            sine_reg0   <= 36'sb100001110101010110010001000010101011;
        end
        11402: begin
            cosine_reg0 <= 36'sb110101010101011100110001001011001010;
            sine_reg0   <= 36'sb100001110101000101100000010100000000;
        end
        11403: begin
            cosine_reg0 <= 36'sb110101010110001100001010011100111101;
            sine_reg0   <= 36'sb100001110100110100110000101111110001;
        end
        11404: begin
            cosine_reg0 <= 36'sb110101010110111011100100001001000010;
            sine_reg0   <= 36'sb100001110100100100000010010101111111;
        end
        11405: begin
            cosine_reg0 <= 36'sb110101010111101010111110001111011000;
            sine_reg0   <= 36'sb100001110100010011010101000110101010;
        end
        11406: begin
            cosine_reg0 <= 36'sb110101011000011010011000101111111101;
            sine_reg0   <= 36'sb100001110100000010101001000001110100;
        end
        11407: begin
            cosine_reg0 <= 36'sb110101011001001001110011101010101110;
            sine_reg0   <= 36'sb100001110011110001111110000111011101;
        end
        11408: begin
            cosine_reg0 <= 36'sb110101011001111001001110111111101010;
            sine_reg0   <= 36'sb100001110011100001010100010111100101;
        end
        11409: begin
            cosine_reg0 <= 36'sb110101011010101000101010101110110000;
            sine_reg0   <= 36'sb100001110011010000101011110010001101;
        end
        11410: begin
            cosine_reg0 <= 36'sb110101011011011000000110110111111101;
            sine_reg0   <= 36'sb100001110011000000000100010111010110;
        end
        11411: begin
            cosine_reg0 <= 36'sb110101011100000111100011011011001111;
            sine_reg0   <= 36'sb100001110010101111011110000111000001;
        end
        11412: begin
            cosine_reg0 <= 36'sb110101011100110111000000011000100101;
            sine_reg0   <= 36'sb100001110010011110111001000001001110;
        end
        11413: begin
            cosine_reg0 <= 36'sb110101011101100110011101101111111101;
            sine_reg0   <= 36'sb100001110010001110010101000101111110;
        end
        11414: begin
            cosine_reg0 <= 36'sb110101011110010101111011100001010101;
            sine_reg0   <= 36'sb100001110001111101110010010101010001;
        end
        11415: begin
            cosine_reg0 <= 36'sb110101011111000101011001101100101011;
            sine_reg0   <= 36'sb100001110001101101010000101111001000;
        end
        11416: begin
            cosine_reg0 <= 36'sb110101011111110100111000010001111101;
            sine_reg0   <= 36'sb100001110001011100110000010011100011;
        end
        11417: begin
            cosine_reg0 <= 36'sb110101100000100100010111010001001010;
            sine_reg0   <= 36'sb100001110001001100010001000010100101;
        end
        11418: begin
            cosine_reg0 <= 36'sb110101100001010011110110101010010000;
            sine_reg0   <= 36'sb100001110000111011110010111100001100;
        end
        11419: begin
            cosine_reg0 <= 36'sb110101100010000011010110011101001100;
            sine_reg0   <= 36'sb100001110000101011010110000000011001;
        end
        11420: begin
            cosine_reg0 <= 36'sb110101100010110010110110101001111110;
            sine_reg0   <= 36'sb100001110000011010111010001111001110;
        end
        11421: begin
            cosine_reg0 <= 36'sb110101100011100010010111010000100010;
            sine_reg0   <= 36'sb100001110000001010011111101000101011;
        end
        11422: begin
            cosine_reg0 <= 36'sb110101100100010001111000010000111000;
            sine_reg0   <= 36'sb100001101111111010000110001100110000;
        end
        11423: begin
            cosine_reg0 <= 36'sb110101100101000001011001101010111110;
            sine_reg0   <= 36'sb100001101111101001101101111011011110;
        end
        11424: begin
            cosine_reg0 <= 36'sb110101100101110000111011011110110001;
            sine_reg0   <= 36'sb100001101111011001010110110100110110;
        end
        11425: begin
            cosine_reg0 <= 36'sb110101100110100000011101101100010000;
            sine_reg0   <= 36'sb100001101111001001000000111000111000;
        end
        11426: begin
            cosine_reg0 <= 36'sb110101100111010000000000010011011010;
            sine_reg0   <= 36'sb100001101110111000101100000111100110;
        end
        11427: begin
            cosine_reg0 <= 36'sb110101100111111111100011010100001011;
            sine_reg0   <= 36'sb100001101110101000011000100000111111;
        end
        11428: begin
            cosine_reg0 <= 36'sb110101101000101111000110101110100011;
            sine_reg0   <= 36'sb100001101110011000000110000101000100;
        end
        11429: begin
            cosine_reg0 <= 36'sb110101101001011110101010100010011111;
            sine_reg0   <= 36'sb100001101110000111110100110011110110;
        end
        11430: begin
            cosine_reg0 <= 36'sb110101101010001110001110101111111110;
            sine_reg0   <= 36'sb100001101101110111100100101101010110;
        end
        11431: begin
            cosine_reg0 <= 36'sb110101101010111101110011010110111110;
            sine_reg0   <= 36'sb100001101101100111010101110001100100;
        end
        11432: begin
            cosine_reg0 <= 36'sb110101101011101101011000010111011101;
            sine_reg0   <= 36'sb100001101101010111001000000000100000;
        end
        11433: begin
            cosine_reg0 <= 36'sb110101101100011100111101110001011001;
            sine_reg0   <= 36'sb100001101101000110111011011010001101;
        end
        11434: begin
            cosine_reg0 <= 36'sb110101101101001100100011100100110001;
            sine_reg0   <= 36'sb100001101100110110101111111110101001;
        end
        11435: begin
            cosine_reg0 <= 36'sb110101101101111100001001110001100010;
            sine_reg0   <= 36'sb100001101100100110100101101101110101;
        end
        11436: begin
            cosine_reg0 <= 36'sb110101101110101011110000010111101010;
            sine_reg0   <= 36'sb100001101100010110011100100111110011;
        end
        11437: begin
            cosine_reg0 <= 36'sb110101101111011011010111010111001001;
            sine_reg0   <= 36'sb100001101100000110010100101100100011;
        end
        11438: begin
            cosine_reg0 <= 36'sb110101110000001010111110101111111011;
            sine_reg0   <= 36'sb100001101011110110001101111100000110;
        end
        11439: begin
            cosine_reg0 <= 36'sb110101110000111010100110100010000000;
            sine_reg0   <= 36'sb100001101011100110001000010110011011;
        end
        11440: begin
            cosine_reg0 <= 36'sb110101110001101010001110101101010101;
            sine_reg0   <= 36'sb100001101011010110000011111011100100;
        end
        11441: begin
            cosine_reg0 <= 36'sb110101110010011001110111010001111001;
            sine_reg0   <= 36'sb100001101011000110000000101011100010;
        end
        11442: begin
            cosine_reg0 <= 36'sb110101110011001001100000001111101001;
            sine_reg0   <= 36'sb100001101010110101111110100110010101;
        end
        11443: begin
            cosine_reg0 <= 36'sb110101110011111001001001100110100101;
            sine_reg0   <= 36'sb100001101010100101111101101011111101;
        end
        11444: begin
            cosine_reg0 <= 36'sb110101110100101000110011010110101001;
            sine_reg0   <= 36'sb100001101010010101111101111100011011;
        end
        11445: begin
            cosine_reg0 <= 36'sb110101110101011000011101011111110100;
            sine_reg0   <= 36'sb100001101010000101111111010111110001;
        end
        11446: begin
            cosine_reg0 <= 36'sb110101110110001000001000000010000101;
            sine_reg0   <= 36'sb100001101001110110000001111101111101;
        end
        11447: begin
            cosine_reg0 <= 36'sb110101110110110111110010111101011001;
            sine_reg0   <= 36'sb100001101001100110000101101111000010;
        end
        11448: begin
            cosine_reg0 <= 36'sb110101110111100111011110010001101111;
            sine_reg0   <= 36'sb100001101001010110001010101011000000;
        end
        11449: begin
            cosine_reg0 <= 36'sb110101111000010111001001111111000101;
            sine_reg0   <= 36'sb100001101001000110010000110001110111;
        end
        11450: begin
            cosine_reg0 <= 36'sb110101111001000110110110000101011001;
            sine_reg0   <= 36'sb100001101000110110011000000011100111;
        end
        11451: begin
            cosine_reg0 <= 36'sb110101111001110110100010100100101000;
            sine_reg0   <= 36'sb100001101000100110100000100000010011;
        end
        11452: begin
            cosine_reg0 <= 36'sb110101111010100110001111011100110011;
            sine_reg0   <= 36'sb100001101000010110101010000111111001;
        end
        11453: begin
            cosine_reg0 <= 36'sb110101111011010101111100101101110101;
            sine_reg0   <= 36'sb100001101000000110110100111010011011;
        end
        11454: begin
            cosine_reg0 <= 36'sb110101111100000101101010010111101110;
            sine_reg0   <= 36'sb100001100111110111000000110111111010;
        end
        11455: begin
            cosine_reg0 <= 36'sb110101111100110101011000011010011100;
            sine_reg0   <= 36'sb100001100111100111001110000000010110;
        end
        11456: begin
            cosine_reg0 <= 36'sb110101111101100101000110110101111101;
            sine_reg0   <= 36'sb100001100111010111011100010011101111;
        end
        11457: begin
            cosine_reg0 <= 36'sb110101111110010100110101101010001111;
            sine_reg0   <= 36'sb100001100111000111101011110010000110;
        end
        11458: begin
            cosine_reg0 <= 36'sb110101111111000100100100110111010001;
            sine_reg0   <= 36'sb100001100110110111111100011011011100;
        end
        11459: begin
            cosine_reg0 <= 36'sb110101111111110100010100011101000000;
            sine_reg0   <= 36'sb100001100110101000001110001111110010;
        end
        11460: begin
            cosine_reg0 <= 36'sb110110000000100100000100011011011010;
            sine_reg0   <= 36'sb100001100110011000100001001111000111;
        end
        11461: begin
            cosine_reg0 <= 36'sb110110000001010011110100110010011110;
            sine_reg0   <= 36'sb100001100110001000110101011001011101;
        end
        11462: begin
            cosine_reg0 <= 36'sb110110000010000011100101100010001010;
            sine_reg0   <= 36'sb100001100101111001001010101110110101;
        end
        11463: begin
            cosine_reg0 <= 36'sb110110000010110011010110101010011100;
            sine_reg0   <= 36'sb100001100101101001100001001111001110;
        end
        11464: begin
            cosine_reg0 <= 36'sb110110000011100011001000001011010010;
            sine_reg0   <= 36'sb100001100101011001111000111010101010;
        end
        11465: begin
            cosine_reg0 <= 36'sb110110000100010010111010000100101011;
            sine_reg0   <= 36'sb100001100101001010010001110001001000;
        end
        11466: begin
            cosine_reg0 <= 36'sb110110000101000010101100010110100100;
            sine_reg0   <= 36'sb100001100100111010101011110010101011;
        end
        11467: begin
            cosine_reg0 <= 36'sb110110000101110010011111000000111100;
            sine_reg0   <= 36'sb100001100100101011000110111111010001;
        end
        11468: begin
            cosine_reg0 <= 36'sb110110000110100010010010000011110001;
            sine_reg0   <= 36'sb100001100100011011100011010110111100;
        end
        11469: begin
            cosine_reg0 <= 36'sb110110000111010010000101011111000001;
            sine_reg0   <= 36'sb100001100100001100000000111001101101;
        end
        11470: begin
            cosine_reg0 <= 36'sb110110001000000001111001010010101010;
            sine_reg0   <= 36'sb100001100011111100011111100111100100;
        end
        11471: begin
            cosine_reg0 <= 36'sb110110001000110001101101011110101010;
            sine_reg0   <= 36'sb100001100011101100111111100000100010;
        end
        11472: begin
            cosine_reg0 <= 36'sb110110001001100001100010000011000000;
            sine_reg0   <= 36'sb100001100011011101100000100100100110;
        end
        11473: begin
            cosine_reg0 <= 36'sb110110001010010001010110111111101001;
            sine_reg0   <= 36'sb100001100011001110000010110011110011;
        end
        11474: begin
            cosine_reg0 <= 36'sb110110001011000001001100010100100100;
            sine_reg0   <= 36'sb100001100010111110100110001110001000;
        end
        11475: begin
            cosine_reg0 <= 36'sb110110001011110001000010000001110000;
            sine_reg0   <= 36'sb100001100010101111001010110011100110;
        end
        11476: begin
            cosine_reg0 <= 36'sb110110001100100000111000000111001001;
            sine_reg0   <= 36'sb100001100010011111110000100100001101;
        end
        11477: begin
            cosine_reg0 <= 36'sb110110001101010000101110100100101110;
            sine_reg0   <= 36'sb100001100010010000010111011111111111;
        end
        11478: begin
            cosine_reg0 <= 36'sb110110001110000000100101011010011110;
            sine_reg0   <= 36'sb100001100010000000111111100110111100;
        end
        11479: begin
            cosine_reg0 <= 36'sb110110001110110000011100101000010111;
            sine_reg0   <= 36'sb100001100001110001101000111001000100;
        end
        11480: begin
            cosine_reg0 <= 36'sb110110001111100000010100001110010110;
            sine_reg0   <= 36'sb100001100001100010010011010110011000;
        end
        11481: begin
            cosine_reg0 <= 36'sb110110010000010000001100001100011010;
            sine_reg0   <= 36'sb100001100001010010111110111110111000;
        end
        11482: begin
            cosine_reg0 <= 36'sb110110010001000000000100100010100001;
            sine_reg0   <= 36'sb100001100001000011101011110010100110;
        end
        11483: begin
            cosine_reg0 <= 36'sb110110010001101111111101010000101001;
            sine_reg0   <= 36'sb100001100000110100011001110001100001;
        end
        11484: begin
            cosine_reg0 <= 36'sb110110010010011111110110010110110001;
            sine_reg0   <= 36'sb100001100000100101001000111011101011;
        end
        11485: begin
            cosine_reg0 <= 36'sb110110010011001111101111110100110110;
            sine_reg0   <= 36'sb100001100000010101111001010001000100;
        end
        11486: begin
            cosine_reg0 <= 36'sb110110010011111111101001101010110111;
            sine_reg0   <= 36'sb100001100000000110101010110001101100;
        end
        11487: begin
            cosine_reg0 <= 36'sb110110010100101111100011111000110010;
            sine_reg0   <= 36'sb100001011111110111011101011101100101;
        end
        11488: begin
            cosine_reg0 <= 36'sb110110010101011111011110011110100100;
            sine_reg0   <= 36'sb100001011111101000010001010100101110;
        end
        11489: begin
            cosine_reg0 <= 36'sb110110010110001111011001011100001101;
            sine_reg0   <= 36'sb100001011111011001000110010111001000;
        end
        11490: begin
            cosine_reg0 <= 36'sb110110010110111111010100110001101010;
            sine_reg0   <= 36'sb100001011111001001111100100100110100;
        end
        11491: begin
            cosine_reg0 <= 36'sb110110010111101111010000011110111001;
            sine_reg0   <= 36'sb100001011110111010110011111101110011;
        end
        11492: begin
            cosine_reg0 <= 36'sb110110011000011111001100100011111001;
            sine_reg0   <= 36'sb100001011110101011101100100010000101;
        end
        11493: begin
            cosine_reg0 <= 36'sb110110011001001111001001000000101000;
            sine_reg0   <= 36'sb100001011110011100100110010001101010;
        end
        11494: begin
            cosine_reg0 <= 36'sb110110011001111111000101110101000011;
            sine_reg0   <= 36'sb100001011110001101100001001100100100;
        end
        11495: begin
            cosine_reg0 <= 36'sb110110011010101111000011000001001010;
            sine_reg0   <= 36'sb100001011101111110011101010010110010;
        end
        11496: begin
            cosine_reg0 <= 36'sb110110011011011111000000100100111001;
            sine_reg0   <= 36'sb100001011101101111011010100100010110;
        end
        11497: begin
            cosine_reg0 <= 36'sb110110011100001110111110100000010000;
            sine_reg0   <= 36'sb100001011101100000011001000001001111;
        end
        11498: begin
            cosine_reg0 <= 36'sb110110011100111110111100110011001101;
            sine_reg0   <= 36'sb100001011101010001011000101001011111;
        end
        11499: begin
            cosine_reg0 <= 36'sb110110011101101110111011011101101101;
            sine_reg0   <= 36'sb100001011101000010011001011101000111;
        end
        11500: begin
            cosine_reg0 <= 36'sb110110011110011110111010011111101111;
            sine_reg0   <= 36'sb100001011100110011011011011100000110;
        end
        11501: begin
            cosine_reg0 <= 36'sb110110011111001110111001111001010000;
            sine_reg0   <= 36'sb100001011100100100011110100110011101;
        end
        11502: begin
            cosine_reg0 <= 36'sb110110011111111110111001101010010000;
            sine_reg0   <= 36'sb100001011100010101100010111100001101;
        end
        11503: begin
            cosine_reg0 <= 36'sb110110100000101110111001110010101100;
            sine_reg0   <= 36'sb100001011100000110101000011101010110;
        end
        11504: begin
            cosine_reg0 <= 36'sb110110100001011110111010010010100011;
            sine_reg0   <= 36'sb100001011011110111101111001001111001;
        end
        11505: begin
            cosine_reg0 <= 36'sb110110100010001110111011001001110010;
            sine_reg0   <= 36'sb100001011011101000110111000001110111;
        end
        11506: begin
            cosine_reg0 <= 36'sb110110100010111110111100011000010111;
            sine_reg0   <= 36'sb100001011011011010000000000101010000;
        end
        11507: begin
            cosine_reg0 <= 36'sb110110100011101110111101111110010010;
            sine_reg0   <= 36'sb100001011011001011001010010100000101;
        end
        11508: begin
            cosine_reg0 <= 36'sb110110100100011110111111111011011111;
            sine_reg0   <= 36'sb100001011010111100010101101110010110;
        end
        11509: begin
            cosine_reg0 <= 36'sb110110100101001111000010001111111110;
            sine_reg0   <= 36'sb100001011010101101100010010100000100;
        end
        11510: begin
            cosine_reg0 <= 36'sb110110100101111111000100111011101100;
            sine_reg0   <= 36'sb100001011010011110110000000101001111;
        end
        11511: begin
            cosine_reg0 <= 36'sb110110100110101111000111111110100111;
            sine_reg0   <= 36'sb100001011010001111111111000001111001;
        end
        11512: begin
            cosine_reg0 <= 36'sb110110100111011111001011011000101110;
            sine_reg0   <= 36'sb100001011010000001001111001010000001;
        end
        11513: begin
            cosine_reg0 <= 36'sb110110101000001111001111001001111110;
            sine_reg0   <= 36'sb100001011001110010100000011101101000;
        end
        11514: begin
            cosine_reg0 <= 36'sb110110101000111111010011010010010110;
            sine_reg0   <= 36'sb100001011001100011110010111100101110;
        end
        11515: begin
            cosine_reg0 <= 36'sb110110101001101111010111110001110101;
            sine_reg0   <= 36'sb100001011001010101000110100111010101;
        end
        11516: begin
            cosine_reg0 <= 36'sb110110101010011111011100101000010111;
            sine_reg0   <= 36'sb100001011001000110011011011101011101;
        end
        11517: begin
            cosine_reg0 <= 36'sb110110101011001111100001110101111100;
            sine_reg0   <= 36'sb100001011000110111110001011111000110;
        end
        11518: begin
            cosine_reg0 <= 36'sb110110101011111111100111011010100001;
            sine_reg0   <= 36'sb100001011000101001001000101100010001;
        end
        11519: begin
            cosine_reg0 <= 36'sb110110101100101111101101010110000101;
            sine_reg0   <= 36'sb100001011000011010100001000100111111;
        end
        11520: begin
            cosine_reg0 <= 36'sb110110101101011111110011101000100110;
            sine_reg0   <= 36'sb100001011000001011111010101001001111;
        end
        11521: begin
            cosine_reg0 <= 36'sb110110101110001111111010010010000001;
            sine_reg0   <= 36'sb100001010111111101010101011001000100;
        end
        11522: begin
            cosine_reg0 <= 36'sb110110101111000000000001010010010101;
            sine_reg0   <= 36'sb100001010111101110110001010100011100;
        end
        11523: begin
            cosine_reg0 <= 36'sb110110101111110000001000101001100001;
            sine_reg0   <= 36'sb100001010111100000001110011011011010;
        end
        11524: begin
            cosine_reg0 <= 36'sb110110110000100000010000010111100010;
            sine_reg0   <= 36'sb100001010111010001101100101101111100;
        end
        11525: begin
            cosine_reg0 <= 36'sb110110110001010000011000011100010110;
            sine_reg0   <= 36'sb100001010111000011001100001100000101;
        end
        11526: begin
            cosine_reg0 <= 36'sb110110110010000000100000110111111100;
            sine_reg0   <= 36'sb100001010110110100101100110101110100;
        end
        11527: begin
            cosine_reg0 <= 36'sb110110110010110000101001101010010010;
            sine_reg0   <= 36'sb100001010110100110001110101011001010;
        end
        11528: begin
            cosine_reg0 <= 36'sb110110110011100000110010110011010110;
            sine_reg0   <= 36'sb100001010110010111110001101100000111;
        end
        11529: begin
            cosine_reg0 <= 36'sb110110110100010000111100010011000101;
            sine_reg0   <= 36'sb100001010110001001010101111000101101;
        end
        11530: begin
            cosine_reg0 <= 36'sb110110110101000001000110001001011111;
            sine_reg0   <= 36'sb100001010101111010111011010000111011;
        end
        11531: begin
            cosine_reg0 <= 36'sb110110110101110001010000010110100001;
            sine_reg0   <= 36'sb100001010101101100100001110100110011;
        end
        11532: begin
            cosine_reg0 <= 36'sb110110110110100001011010111010001010;
            sine_reg0   <= 36'sb100001010101011110001001100100010100;
        end
        11533: begin
            cosine_reg0 <= 36'sb110110110111010001100101110100010111;
            sine_reg0   <= 36'sb100001010101001111110010011111100000;
        end
        11534: begin
            cosine_reg0 <= 36'sb110110111000000001110001000101000111;
            sine_reg0   <= 36'sb100001010101000001011100100110010111;
        end
        11535: begin
            cosine_reg0 <= 36'sb110110111000110001111100101100011000;
            sine_reg0   <= 36'sb100001010100110011000111111000111001;
        end
        11536: begin
            cosine_reg0 <= 36'sb110110111001100010001000101010001000;
            sine_reg0   <= 36'sb100001010100100100110100010111000111;
        end
        11537: begin
            cosine_reg0 <= 36'sb110110111010010010010100111110010101;
            sine_reg0   <= 36'sb100001010100010110100010000001000010;
        end
        11538: begin
            cosine_reg0 <= 36'sb110110111011000010100001101000111101;
            sine_reg0   <= 36'sb100001010100001000010000110110101001;
        end
        11539: begin
            cosine_reg0 <= 36'sb110110111011110010101110101001111111;
            sine_reg0   <= 36'sb100001010011111010000000110111111111;
        end
        11540: begin
            cosine_reg0 <= 36'sb110110111100100010111100000001011001;
            sine_reg0   <= 36'sb100001010011101011110010000101000011;
        end
        11541: begin
            cosine_reg0 <= 36'sb110110111101010011001001101111001000;
            sine_reg0   <= 36'sb100001010011011101100100011101110101;
        end
        11542: begin
            cosine_reg0 <= 36'sb110110111110000011010111110011001011;
            sine_reg0   <= 36'sb100001010011001111011000000010010111;
        end
        11543: begin
            cosine_reg0 <= 36'sb110110111110110011100110001101100000;
            sine_reg0   <= 36'sb100001010011000001001100110010101000;
        end
        11544: begin
            cosine_reg0 <= 36'sb110110111111100011110100111110000101;
            sine_reg0   <= 36'sb100001010010110011000010101110101010;
        end
        11545: begin
            cosine_reg0 <= 36'sb110111000000010100000100000100111001;
            sine_reg0   <= 36'sb100001010010100100111001110110011101;
        end
        11546: begin
            cosine_reg0 <= 36'sb110111000001000100010011100001111001;
            sine_reg0   <= 36'sb100001010010010110110010001010000001;
        end
        11547: begin
            cosine_reg0 <= 36'sb110111000001110100100011010101000100;
            sine_reg0   <= 36'sb100001010010001000101011101001011000;
        end
        11548: begin
            cosine_reg0 <= 36'sb110111000010100100110011011110010111;
            sine_reg0   <= 36'sb100001010001111010100110010100100001;
        end
        11549: begin
            cosine_reg0 <= 36'sb110111000011010101000011111101110001;
            sine_reg0   <= 36'sb100001010001101100100010001011011101;
        end
        11550: begin
            cosine_reg0 <= 36'sb110111000100000101010100110011010001;
            sine_reg0   <= 36'sb100001010001011110011111001110001101;
        end
        11551: begin
            cosine_reg0 <= 36'sb110111000100110101100101111110110011;
            sine_reg0   <= 36'sb100001010001010000011101011100110000;
        end
        11552: begin
            cosine_reg0 <= 36'sb110111000101100101110111100000010111;
            sine_reg0   <= 36'sb100001010001000010011100110111001001;
        end
        11553: begin
            cosine_reg0 <= 36'sb110111000110010110001001010111111010;
            sine_reg0   <= 36'sb100001010000110100011101011101010111;
        end
        11554: begin
            cosine_reg0 <= 36'sb110111000111000110011011100101011010;
            sine_reg0   <= 36'sb100001010000100110011111001111011011;
        end
        11555: begin
            cosine_reg0 <= 36'sb110111000111110110101110001000110111;
            sine_reg0   <= 36'sb100001010000011000100010001101010101;
        end
        11556: begin
            cosine_reg0 <= 36'sb110111001000100111000001000010001101;
            sine_reg0   <= 36'sb100001010000001010100110010111000110;
        end
        11557: begin
            cosine_reg0 <= 36'sb110111001001010111010100010001011011;
            sine_reg0   <= 36'sb100001001111111100101011101100101111;
        end
        11558: begin
            cosine_reg0 <= 36'sb110111001010000111100111110110100000;
            sine_reg0   <= 36'sb100001001111101110110010001110001111;
        end
        11559: begin
            cosine_reg0 <= 36'sb110111001010110111111011110001011000;
            sine_reg0   <= 36'sb100001001111100000111001111011101000;
        end
        11560: begin
            cosine_reg0 <= 36'sb110111001011101000010000000010000011;
            sine_reg0   <= 36'sb100001001111010011000010110100111010;
        end
        11561: begin
            cosine_reg0 <= 36'sb110111001100011000100100101000011111;
            sine_reg0   <= 36'sb100001001111000101001100111010000110;
        end
        11562: begin
            cosine_reg0 <= 36'sb110111001101001000111001100100101001;
            sine_reg0   <= 36'sb100001001110110111011000001011001100;
        end
        11563: begin
            cosine_reg0 <= 36'sb110111001101111001001110110110100000;
            sine_reg0   <= 36'sb100001001110101001100100101000001100;
        end
        11564: begin
            cosine_reg0 <= 36'sb110111001110101001100100011110000010;
            sine_reg0   <= 36'sb100001001110011011110010010001000111;
        end
        11565: begin
            cosine_reg0 <= 36'sb110111001111011001111010011011001101;
            sine_reg0   <= 36'sb100001001110001110000001000101111111;
        end
        11566: begin
            cosine_reg0 <= 36'sb110111010000001010010000101101111111;
            sine_reg0   <= 36'sb100001001110000000010001000110110010;
        end
        11567: begin
            cosine_reg0 <= 36'sb110111010000111010100111010110010110;
            sine_reg0   <= 36'sb100001001101110010100010010011100010;
        end
        11568: begin
            cosine_reg0 <= 36'sb110111010001101010111110010100010001;
            sine_reg0   <= 36'sb100001001101100100110100101100010000;
        end
        11569: begin
            cosine_reg0 <= 36'sb110111010010011011010101100111101110;
            sine_reg0   <= 36'sb100001001101010111001000010000111011;
        end
        11570: begin
            cosine_reg0 <= 36'sb110111010011001011101101010000101011;
            sine_reg0   <= 36'sb100001001101001001011101000001100101;
        end
        11571: begin
            cosine_reg0 <= 36'sb110111010011111100000101001111000101;
            sine_reg0   <= 36'sb100001001100111011110010111110001110;
        end
        11572: begin
            cosine_reg0 <= 36'sb110111010100101100011101100010111011;
            sine_reg0   <= 36'sb100001001100101110001010000110110110;
        end
        11573: begin
            cosine_reg0 <= 36'sb110111010101011100110110001100001100;
            sine_reg0   <= 36'sb100001001100100000100010011011011110;
        end
        11574: begin
            cosine_reg0 <= 36'sb110111010110001101001111001010110100;
            sine_reg0   <= 36'sb100001001100010010111011111100000110;
        end
        11575: begin
            cosine_reg0 <= 36'sb110111010110111101101000011110110100;
            sine_reg0   <= 36'sb100001001100000101010110101000110000;
        end
        11576: begin
            cosine_reg0 <= 36'sb110111010111101110000010001000000111;
            sine_reg0   <= 36'sb100001001011110111110010100001011011;
        end
        11577: begin
            cosine_reg0 <= 36'sb110111011000011110011100000110101110;
            sine_reg0   <= 36'sb100001001011101010001111100110001000;
        end
        11578: begin
            cosine_reg0 <= 36'sb110111011001001110110110011010100101;
            sine_reg0   <= 36'sb100001001011011100101101110110110111;
        end
        11579: begin
            cosine_reg0 <= 36'sb110111011001111111010001000011101100;
            sine_reg0   <= 36'sb100001001011001111001101010011101010;
        end
        11580: begin
            cosine_reg0 <= 36'sb110111011010101111101100000001111111;
            sine_reg0   <= 36'sb100001001011000001101101111100100000;
        end
        11581: begin
            cosine_reg0 <= 36'sb110111011011100000000111010101011101;
            sine_reg0   <= 36'sb100001001010110100001111110001011010;
        end
        11582: begin
            cosine_reg0 <= 36'sb110111011100010000100010111110000101;
            sine_reg0   <= 36'sb100001001010100110110010110010011001;
        end
        11583: begin
            cosine_reg0 <= 36'sb110111011101000000111110111011110101;
            sine_reg0   <= 36'sb100001001010011001010110111111011101;
        end
        11584: begin
            cosine_reg0 <= 36'sb110111011101110001011011001110101010;
            sine_reg0   <= 36'sb100001001010001011111100011000100111;
        end
        11585: begin
            cosine_reg0 <= 36'sb110111011110100001110111110110100011;
            sine_reg0   <= 36'sb100001001001111110100010111101110111;
        end
        11586: begin
            cosine_reg0 <= 36'sb110111011111010010010100110011011110;
            sine_reg0   <= 36'sb100001001001110001001010101111001101;
        end
        11587: begin
            cosine_reg0 <= 36'sb110111100000000010110010000101011000;
            sine_reg0   <= 36'sb100001001001100011110011101100101011;
        end
        11588: begin
            cosine_reg0 <= 36'sb110111100000110011001111101100010001;
            sine_reg0   <= 36'sb100001001001010110011101110110010001;
        end
        11589: begin
            cosine_reg0 <= 36'sb110111100001100011101101101000000111;
            sine_reg0   <= 36'sb100001001001001001001001001011111111;
        end
        11590: begin
            cosine_reg0 <= 36'sb110111100010010100001011111000110110;
            sine_reg0   <= 36'sb100001001000111011110101101101110101;
        end
        11591: begin
            cosine_reg0 <= 36'sb110111100011000100101010011110011110;
            sine_reg0   <= 36'sb100001001000101110100011011011110101;
        end
        11592: begin
            cosine_reg0 <= 36'sb110111100011110101001001011000111101;
            sine_reg0   <= 36'sb100001001000100001010010010101111111;
        end
        11593: begin
            cosine_reg0 <= 36'sb110111100100100101101000101000010001;
            sine_reg0   <= 36'sb100001001000010100000010011100010011;
        end
        11594: begin
            cosine_reg0 <= 36'sb110111100101010110001000001100011000;
            sine_reg0   <= 36'sb100001001000000110110011101110110010;
        end
        11595: begin
            cosine_reg0 <= 36'sb110111100110000110101000000101001111;
            sine_reg0   <= 36'sb100001000111111001100110001101011100;
        end
        11596: begin
            cosine_reg0 <= 36'sb110111100110110111001000010010110110;
            sine_reg0   <= 36'sb100001000111101100011001111000010010;
        end
        11597: begin
            cosine_reg0 <= 36'sb110111100111100111101000110101001011;
            sine_reg0   <= 36'sb100001000111011111001110101111010100;
        end
        11598: begin
            cosine_reg0 <= 36'sb110111101000011000001001101100001010;
            sine_reg0   <= 36'sb100001000111010010000100110010100011;
        end
        11599: begin
            cosine_reg0 <= 36'sb110111101001001000101010110111110100;
            sine_reg0   <= 36'sb100001000111000100111100000010000000;
        end
        11600: begin
            cosine_reg0 <= 36'sb110111101001111001001100011000000101;
            sine_reg0   <= 36'sb100001000110110111110100011101101010;
        end
        11601: begin
            cosine_reg0 <= 36'sb110111101010101001101110001100111100;
            sine_reg0   <= 36'sb100001000110101010101110000101100011;
        end
        11602: begin
            cosine_reg0 <= 36'sb110111101011011010010000010110010111;
            sine_reg0   <= 36'sb100001000110011101101000111001101011;
        end
        11603: begin
            cosine_reg0 <= 36'sb110111101100001010110010110100010100;
            sine_reg0   <= 36'sb100001000110010000100100111010000010;
        end
        11604: begin
            cosine_reg0 <= 36'sb110111101100111011010101100110110001;
            sine_reg0   <= 36'sb100001000110000011100010000110101001;
        end
        11605: begin
            cosine_reg0 <= 36'sb110111101101101011111000101101101100;
            sine_reg0   <= 36'sb100001000101110110100000011111100000;
        end
        11606: begin
            cosine_reg0 <= 36'sb110111101110011100011100001001000101;
            sine_reg0   <= 36'sb100001000101101001100000000100101000;
        end
        11607: begin
            cosine_reg0 <= 36'sb110111101111001100111111111000110111;
            sine_reg0   <= 36'sb100001000101011100100000110110000001;
        end
        11608: begin
            cosine_reg0 <= 36'sb110111101111111101100011111101000011;
            sine_reg0   <= 36'sb100001000101001111100010110011101101;
        end
        11609: begin
            cosine_reg0 <= 36'sb110111110000101110001000010101100101;
            sine_reg0   <= 36'sb100001000101000010100101111101101011;
        end
        11610: begin
            cosine_reg0 <= 36'sb110111110001011110101101000010011101;
            sine_reg0   <= 36'sb100001000100110101101010010011111011;
        end
        11611: begin
            cosine_reg0 <= 36'sb110111110010001111010010000011100111;
            sine_reg0   <= 36'sb100001000100101000101111110110011111;
        end
        11612: begin
            cosine_reg0 <= 36'sb110111110010111111110111011001000011;
            sine_reg0   <= 36'sb100001000100011011110110100101010111;
        end
        11613: begin
            cosine_reg0 <= 36'sb110111110011110000011101000010101110;
            sine_reg0   <= 36'sb100001000100001110111110100000100100;
        end
        11614: begin
            cosine_reg0 <= 36'sb110111110100100001000011000000100111;
            sine_reg0   <= 36'sb100001000100000010000111101000000101;
        end
        11615: begin
            cosine_reg0 <= 36'sb110111110101010001101001010010101011;
            sine_reg0   <= 36'sb100001000011110101010001111011111011;
        end
        11616: begin
            cosine_reg0 <= 36'sb110111110110000010001111111000111001;
            sine_reg0   <= 36'sb100001000011101000011101011100001000;
        end
        11617: begin
            cosine_reg0 <= 36'sb110111110110110010110110110011001111;
            sine_reg0   <= 36'sb100001000011011011101010001000101011;
        end
        11618: begin
            cosine_reg0 <= 36'sb110111110111100011011110000001101011;
            sine_reg0   <= 36'sb100001000011001110111000000001100100;
        end
        11619: begin
            cosine_reg0 <= 36'sb110111111000010100000101100100001011;
            sine_reg0   <= 36'sb100001000011000010000111000110110101;
        end
        11620: begin
            cosine_reg0 <= 36'sb110111111001000100101101011010101110;
            sine_reg0   <= 36'sb100001000010110101010111011000011110;
        end
        11621: begin
            cosine_reg0 <= 36'sb110111111001110101010101100101010001;
            sine_reg0   <= 36'sb100001000010101000101000110110011111;
        end
        11622: begin
            cosine_reg0 <= 36'sb110111111010100101111110000011110010;
            sine_reg0   <= 36'sb100001000010011011111011100000111001;
        end
        11623: begin
            cosine_reg0 <= 36'sb110111111011010110100110110110010000;
            sine_reg0   <= 36'sb100001000010001111001111010111101101;
        end
        11624: begin
            cosine_reg0 <= 36'sb110111111100000111001111111100101001;
            sine_reg0   <= 36'sb100001000010000010100100011010111010;
        end
        11625: begin
            cosine_reg0 <= 36'sb110111111100110111111001010110111011;
            sine_reg0   <= 36'sb100001000001110101111010101010100001;
        end
        11626: begin
            cosine_reg0 <= 36'sb110111111101101000100011000101000011;
            sine_reg0   <= 36'sb100001000001101001010010000110100011;
        end
        11627: begin
            cosine_reg0 <= 36'sb110111111110011001001101000111000001;
            sine_reg0   <= 36'sb100001000001011100101010101111000001;
        end
        11628: begin
            cosine_reg0 <= 36'sb110111111111001001110111011100110010;
            sine_reg0   <= 36'sb100001000001010000000100100011111010;
        end
        11629: begin
            cosine_reg0 <= 36'sb110111111111111010100010000110010101;
            sine_reg0   <= 36'sb100001000001000011011111100101001111;
        end
        11630: begin
            cosine_reg0 <= 36'sb111000000000101011001101000011100111;
            sine_reg0   <= 36'sb100001000000110110111011110011000010;
        end
        11631: begin
            cosine_reg0 <= 36'sb111000000001011011111000010100100111;
            sine_reg0   <= 36'sb100001000000101010011001001101010001;
        end
        11632: begin
            cosine_reg0 <= 36'sb111000000010001100100011111001010010;
            sine_reg0   <= 36'sb100001000000011101110111110011111110;
        end
        11633: begin
            cosine_reg0 <= 36'sb111000000010111101001111110001101000;
            sine_reg0   <= 36'sb100001000000010001010111100111001001;
        end
        11634: begin
            cosine_reg0 <= 36'sb111000000011101101111011111101100101;
            sine_reg0   <= 36'sb100001000000000100111000100110110011;
        end
        11635: begin
            cosine_reg0 <= 36'sb111000000100011110101000011101001001;
            sine_reg0   <= 36'sb100000111111111000011010110010111100;
        end
        11636: begin
            cosine_reg0 <= 36'sb111000000101001111010101010000010000;
            sine_reg0   <= 36'sb100000111111101011111110001011100101;
        end
        11637: begin
            cosine_reg0 <= 36'sb111000000110000000000010010110111010;
            sine_reg0   <= 36'sb100000111111011111100010110000101110;
        end
        11638: begin
            cosine_reg0 <= 36'sb111000000110110000101111110001000101;
            sine_reg0   <= 36'sb100000111111010011001000100010010111;
        end
        11639: begin
            cosine_reg0 <= 36'sb111000000111100001011101011110101110;
            sine_reg0   <= 36'sb100000111111000110101111100000100001;
        end
        11640: begin
            cosine_reg0 <= 36'sb111000001000010010001011011111110100;
            sine_reg0   <= 36'sb100000111110111010010111101011001101;
        end
        11641: begin
            cosine_reg0 <= 36'sb111000001001000010111001110100010101;
            sine_reg0   <= 36'sb100000111110101110000001000010011011;
        end
        11642: begin
            cosine_reg0 <= 36'sb111000001001110011101000011100001111;
            sine_reg0   <= 36'sb100000111110100001101011100110001011;
        end
        11643: begin
            cosine_reg0 <= 36'sb111000001010100100010111010111100000;
            sine_reg0   <= 36'sb100000111110010101010111010110011111;
        end
        11644: begin
            cosine_reg0 <= 36'sb111000001011010101000110100110000110;
            sine_reg0   <= 36'sb100000111110001001000100010011010101;
        end
        11645: begin
            cosine_reg0 <= 36'sb111000001100000101110110001000000000;
            sine_reg0   <= 36'sb100000111101111100110010011100110000;
        end
        11646: begin
            cosine_reg0 <= 36'sb111000001100110110100101111101001011;
            sine_reg0   <= 36'sb100000111101110000100001110010101111;
        end
        11647: begin
            cosine_reg0 <= 36'sb111000001101100111010110000101100110;
            sine_reg0   <= 36'sb100000111101100100010010010101010011;
        end
        11648: begin
            cosine_reg0 <= 36'sb111000001110011000000110100001001110;
            sine_reg0   <= 36'sb100000111101011000000100000100011100;
        end
        11649: begin
            cosine_reg0 <= 36'sb111000001111001000110111010000000010;
            sine_reg0   <= 36'sb100000111101001011110111000000001011;
        end
        11650: begin
            cosine_reg0 <= 36'sb111000001111111001101000010010000001;
            sine_reg0   <= 36'sb100000111100111111101011001000100001;
        end
        11651: begin
            cosine_reg0 <= 36'sb111000010000101010011001100111000111;
            sine_reg0   <= 36'sb100000111100110011100000011101011101;
        end
        11652: begin
            cosine_reg0 <= 36'sb111000010001011011001011001111010011;
            sine_reg0   <= 36'sb100000111100100111010110111111000000;
        end
        11653: begin
            cosine_reg0 <= 36'sb111000010010001011111101001010100100;
            sine_reg0   <= 36'sb100000111100011011001110101101001011;
        end
        11654: begin
            cosine_reg0 <= 36'sb111000010010111100101111011000110111;
            sine_reg0   <= 36'sb100000111100001111000111100111111110;
        end
        11655: begin
            cosine_reg0 <= 36'sb111000010011101101100001111010001011;
            sine_reg0   <= 36'sb100000111100000011000001101111011010;
        end
        11656: begin
            cosine_reg0 <= 36'sb111000010100011110010100101110011101;
            sine_reg0   <= 36'sb100000111011110110111101000011011111;
        end
        11657: begin
            cosine_reg0 <= 36'sb111000010101001111000111110101101101;
            sine_reg0   <= 36'sb100000111011101010111001100100001101;
        end
        11658: begin
            cosine_reg0 <= 36'sb111000010101111111111011001111110111;
            sine_reg0   <= 36'sb100000111011011110110111010001100101;
        end
        11659: begin
            cosine_reg0 <= 36'sb111000010110110000101110111100111010;
            sine_reg0   <= 36'sb100000111011010010110110001011101000;
        end
        11660: begin
            cosine_reg0 <= 36'sb111000010111100001100010111100110100;
            sine_reg0   <= 36'sb100000111011000110110110010010010110;
        end
        11661: begin
            cosine_reg0 <= 36'sb111000011000010010010111001111100100;
            sine_reg0   <= 36'sb100000111010111010110111100101101111;
        end
        11662: begin
            cosine_reg0 <= 36'sb111000011001000011001011110101000111;
            sine_reg0   <= 36'sb100000111010101110111010000101110100;
        end
        11663: begin
            cosine_reg0 <= 36'sb111000011001110100000000101101011011;
            sine_reg0   <= 36'sb100000111010100010111101110010100101;
        end
        11664: begin
            cosine_reg0 <= 36'sb111000011010100100110101111000011111;
            sine_reg0   <= 36'sb100000111010010111000010101100000011;
        end
        11665: begin
            cosine_reg0 <= 36'sb111000011011010101101011010110010001;
            sine_reg0   <= 36'sb100000111010001011001000110010001111;
        end
        11666: begin
            cosine_reg0 <= 36'sb111000011100000110100001000110101111;
            sine_reg0   <= 36'sb100000111001111111010000000101001000;
        end
        11667: begin
            cosine_reg0 <= 36'sb111000011100110111010111001001110110;
            sine_reg0   <= 36'sb100000111001110011011000100100101111;
        end
        11668: begin
            cosine_reg0 <= 36'sb111000011101101000001101011111100110;
            sine_reg0   <= 36'sb100000111001100111100010010001000100;
        end
        11669: begin
            cosine_reg0 <= 36'sb111000011110011001000100000111111100;
            sine_reg0   <= 36'sb100000111001011011101101001010001001;
        end
        11670: begin
            cosine_reg0 <= 36'sb111000011111001001111011000010110110;
            sine_reg0   <= 36'sb100000111001001111111001001111111110;
        end
        11671: begin
            cosine_reg0 <= 36'sb111000011111111010110010010000010011;
            sine_reg0   <= 36'sb100000111001000100000110100010100010;
        end
        11672: begin
            cosine_reg0 <= 36'sb111000100000101011101001110000010000;
            sine_reg0   <= 36'sb100000111000111000010101000001110111;
        end
        11673: begin
            cosine_reg0 <= 36'sb111000100001011100100001100010101100;
            sine_reg0   <= 36'sb100000111000101100100100101101111101;
        end
        11674: begin
            cosine_reg0 <= 36'sb111000100010001101011001100111100101;
            sine_reg0   <= 36'sb100000111000100000110101100110110100;
        end
        11675: begin
            cosine_reg0 <= 36'sb111000100010111110010001111110111000;
            sine_reg0   <= 36'sb100000111000010101000111101100011100;
        end
        11676: begin
            cosine_reg0 <= 36'sb111000100011101111001010101000100101;
            sine_reg0   <= 36'sb100000111000001001011010111110111000;
        end
        11677: begin
            cosine_reg0 <= 36'sb111000100100100000000011100100101001;
            sine_reg0   <= 36'sb100000110111111101101111011110000101;
        end
        11678: begin
            cosine_reg0 <= 36'sb111000100101010000111100110011000010;
            sine_reg0   <= 36'sb100000110111110010000101001010000110;
        end
        11679: begin
            cosine_reg0 <= 36'sb111000100110000001110110010011101110;
            sine_reg0   <= 36'sb100000110111100110011100000010111011;
        end
        11680: begin
            cosine_reg0 <= 36'sb111000100110110010110000000110101100;
            sine_reg0   <= 36'sb100000110111011010110100001000100011;
        end
        11681: begin
            cosine_reg0 <= 36'sb111000100111100011101010001011111001;
            sine_reg0   <= 36'sb100000110111001111001101011011000000;
        end
        11682: begin
            cosine_reg0 <= 36'sb111000101000010100100100100011010100;
            sine_reg0   <= 36'sb100000110111000011100111111010010011;
        end
        11683: begin
            cosine_reg0 <= 36'sb111000101001000101011111001100111011;
            sine_reg0   <= 36'sb100000110110111000000011100110011010;
        end
        11684: begin
            cosine_reg0 <= 36'sb111000101001110110011010001000101100;
            sine_reg0   <= 36'sb100000110110101100100000011111010111;
        end
        11685: begin
            cosine_reg0 <= 36'sb111000101010100111010101010110100101;
            sine_reg0   <= 36'sb100000110110100000111110100101001011;
        end
        11686: begin
            cosine_reg0 <= 36'sb111000101011011000010000110110100100;
            sine_reg0   <= 36'sb100000110110010101011101110111110101;
        end
        11687: begin
            cosine_reg0 <= 36'sb111000101100001001001100101000101000;
            sine_reg0   <= 36'sb100000110110001001111110010111010110;
        end
        11688: begin
            cosine_reg0 <= 36'sb111000101100111010001000101100101101;
            sine_reg0   <= 36'sb100000110101111110100000000011101111;
        end
        11689: begin
            cosine_reg0 <= 36'sb111000101101101011000101000010110100;
            sine_reg0   <= 36'sb100000110101110011000010111101000001;
        end
        11690: begin
            cosine_reg0 <= 36'sb111000101110011100000001101010111001;
            sine_reg0   <= 36'sb100000110101100111100111000011001010;
        end
        11691: begin
            cosine_reg0 <= 36'sb111000101111001100111110100100111010;
            sine_reg0   <= 36'sb100000110101011100001100010110001101;
        end
        11692: begin
            cosine_reg0 <= 36'sb111000101111111101111011110000110111;
            sine_reg0   <= 36'sb100000110101010000110010110110001001;
        end
        11693: begin
            cosine_reg0 <= 36'sb111000110000101110111001001110101100;
            sine_reg0   <= 36'sb100000110101000101011010100010111110;
        end
        11694: begin
            cosine_reg0 <= 36'sb111000110001011111110110111110011000;
            sine_reg0   <= 36'sb100000110100111010000011011100101110;
        end
        11695: begin
            cosine_reg0 <= 36'sb111000110010010000110100111111111010;
            sine_reg0   <= 36'sb100000110100101110101101100011011001;
        end
        11696: begin
            cosine_reg0 <= 36'sb111000110011000001110011010011001111;
            sine_reg0   <= 36'sb100000110100100011011000110110111111;
        end
        11697: begin
            cosine_reg0 <= 36'sb111000110011110010110001111000010101;
            sine_reg0   <= 36'sb100000110100011000000101010111100000;
        end
        11698: begin
            cosine_reg0 <= 36'sb111000110100100011110000101111001011;
            sine_reg0   <= 36'sb100000110100001100110011000100111110;
        end
        11699: begin
            cosine_reg0 <= 36'sb111000110101010100101111110111101111;
            sine_reg0   <= 36'sb100000110100000001100001111111010111;
        end
        11700: begin
            cosine_reg0 <= 36'sb111000110110000101101111010001111110;
            sine_reg0   <= 36'sb100000110011110110010010000110101110;
        end
        11701: begin
            cosine_reg0 <= 36'sb111000110110110110101110111101110111;
            sine_reg0   <= 36'sb100000110011101011000011011011000010;
        end
        11702: begin
            cosine_reg0 <= 36'sb111000110111100111101110111011011000;
            sine_reg0   <= 36'sb100000110011011111110101111100010100;
        end
        11703: begin
            cosine_reg0 <= 36'sb111000111000011000101111001010011111;
            sine_reg0   <= 36'sb100000110011010100101001101010100100;
        end
        11704: begin
            cosine_reg0 <= 36'sb111000111001001001101111101011001010;
            sine_reg0   <= 36'sb100000110011001001011110100101110010;
        end
        11705: begin
            cosine_reg0 <= 36'sb111000111001111010110000011101011000;
            sine_reg0   <= 36'sb100000110010111110010100101110000000;
        end
        11706: begin
            cosine_reg0 <= 36'sb111000111010101011110001100001000110;
            sine_reg0   <= 36'sb100000110010110011001100000011001101;
        end
        11707: begin
            cosine_reg0 <= 36'sb111000111011011100110010110110010010;
            sine_reg0   <= 36'sb100000110010101000000100100101011010;
        end
        11708: begin
            cosine_reg0 <= 36'sb111000111100001101110100011100111011;
            sine_reg0   <= 36'sb100000110010011100111110010100100111;
        end
        11709: begin
            cosine_reg0 <= 36'sb111000111100111110110110010100111111;
            sine_reg0   <= 36'sb100000110010010001111001010000110101;
        end
        11710: begin
            cosine_reg0 <= 36'sb111000111101101111111000011110011100;
            sine_reg0   <= 36'sb100000110010000110110101011010000100;
        end
        11711: begin
            cosine_reg0 <= 36'sb111000111110100000111010111001010000;
            sine_reg0   <= 36'sb100000110001111011110010110000010101;
        end
        11712: begin
            cosine_reg0 <= 36'sb111000111111010001111101100101011000;
            sine_reg0   <= 36'sb100000110001110000110001010011101000;
        end
        11713: begin
            cosine_reg0 <= 36'sb111001000000000011000000100010110100;
            sine_reg0   <= 36'sb100000110001100101110001000011111101;
        end
        11714: begin
            cosine_reg0 <= 36'sb111001000000110100000011110001100001;
            sine_reg0   <= 36'sb100000110001011010110010000001010101;
        end
        11715: begin
            cosine_reg0 <= 36'sb111001000001100101000111010001011110;
            sine_reg0   <= 36'sb100000110001001111110100001011110001;
        end
        11716: begin
            cosine_reg0 <= 36'sb111001000010010110001011000010101000;
            sine_reg0   <= 36'sb100000110001000100110111100011010000;
        end
        11717: begin
            cosine_reg0 <= 36'sb111001000011000111001111000100111110;
            sine_reg0   <= 36'sb100000110000111001111100000111110011;
        end
        11718: begin
            cosine_reg0 <= 36'sb111001000011111000010011011000011101;
            sine_reg0   <= 36'sb100000110000101111000001111001011011;
        end
        11719: begin
            cosine_reg0 <= 36'sb111001000100101001010111111101000100;
            sine_reg0   <= 36'sb100000110000100100001000111000001000;
        end
        11720: begin
            cosine_reg0 <= 36'sb111001000101011010011100110010110001;
            sine_reg0   <= 36'sb100000110000011001010001000011111010;
        end
        11721: begin
            cosine_reg0 <= 36'sb111001000110001011100001111001100010;
            sine_reg0   <= 36'sb100000110000001110011010011100110010;
        end
        11722: begin
            cosine_reg0 <= 36'sb111001000110111100100111010001010110;
            sine_reg0   <= 36'sb100000110000000011100101000010110000;
        end
        11723: begin
            cosine_reg0 <= 36'sb111001000111101101101100111010001001;
            sine_reg0   <= 36'sb100000101111111000110000110101110101;
        end
        11724: begin
            cosine_reg0 <= 36'sb111001001000011110110010110011111011;
            sine_reg0   <= 36'sb100000101111101101111101110110000010;
        end
        11725: begin
            cosine_reg0 <= 36'sb111001001001001111111000111110101001;
            sine_reg0   <= 36'sb100000101111100011001100000011010101;
        end
        11726: begin
            cosine_reg0 <= 36'sb111001001010000000111111011010010010;
            sine_reg0   <= 36'sb100000101111011000011011011101110001;
        end
        11727: begin
            cosine_reg0 <= 36'sb111001001010110010000110000110110100;
            sine_reg0   <= 36'sb100000101111001101101100000101010101;
        end
        11728: begin
            cosine_reg0 <= 36'sb111001001011100011001101000100001100;
            sine_reg0   <= 36'sb100000101111000010111101111010000001;
        end
        11729: begin
            cosine_reg0 <= 36'sb111001001100010100010100010010011010;
            sine_reg0   <= 36'sb100000101110111000010000111011110111;
        end
        11730: begin
            cosine_reg0 <= 36'sb111001001101000101011011110001011010;
            sine_reg0   <= 36'sb100000101110101101100101001010110110;
        end
        11731: begin
            cosine_reg0 <= 36'sb111001001101110110100011100001001011;
            sine_reg0   <= 36'sb100000101110100010111010100110111111;
        end
        11732: begin
            cosine_reg0 <= 36'sb111001001110100111101011100001101100;
            sine_reg0   <= 36'sb100000101110011000010001010000010011;
        end
        11733: begin
            cosine_reg0 <= 36'sb111001001111011000110011110010111010;
            sine_reg0   <= 36'sb100000101110001101101001000110110010;
        end
        11734: begin
            cosine_reg0 <= 36'sb111001010000001001111100010100110011;
            sine_reg0   <= 36'sb100000101110000011000010001010011011;
        end
        11735: begin
            cosine_reg0 <= 36'sb111001010000111011000101000111010110;
            sine_reg0   <= 36'sb100000101101111000011100011011010000;
        end
        11736: begin
            cosine_reg0 <= 36'sb111001010001101100001110001010100001;
            sine_reg0   <= 36'sb100000101101101101110111111001010010;
        end
        11737: begin
            cosine_reg0 <= 36'sb111001010010011101010111011110010001;
            sine_reg0   <= 36'sb100000101101100011010100100100100000;
        end
        11738: begin
            cosine_reg0 <= 36'sb111001010011001110100001000010100101;
            sine_reg0   <= 36'sb100000101101011000110010011100111010;
        end
        11739: begin
            cosine_reg0 <= 36'sb111001010011111111101010110111011100;
            sine_reg0   <= 36'sb100000101101001110010001100010100010;
        end
        11740: begin
            cosine_reg0 <= 36'sb111001010100110000110100111100110010;
            sine_reg0   <= 36'sb100000101101000011110001110101011000;
        end
        11741: begin
            cosine_reg0 <= 36'sb111001010101100001111111010010100110;
            sine_reg0   <= 36'sb100000101100111001010011010101011011;
        end
        11742: begin
            cosine_reg0 <= 36'sb111001010110010011001001111000110111;
            sine_reg0   <= 36'sb100000101100101110110110000010101101;
        end
        11743: begin
            cosine_reg0 <= 36'sb111001010111000100010100101111100010;
            sine_reg0   <= 36'sb100000101100100100011001111101001110;
        end
        11744: begin
            cosine_reg0 <= 36'sb111001010111110101011111110110100101;
            sine_reg0   <= 36'sb100000101100011001111111000100111110;
        end
        11745: begin
            cosine_reg0 <= 36'sb111001011000100110101011001101111111;
            sine_reg0   <= 36'sb100000101100001111100101011001111110;
        end
        11746: begin
            cosine_reg0 <= 36'sb111001011001010111110110110101101110;
            sine_reg0   <= 36'sb100000101100000101001100111100001110;
        end
        11747: begin
            cosine_reg0 <= 36'sb111001011010001001000010101101110000;
            sine_reg0   <= 36'sb100000101011111010110101101011101110;
        end
        11748: begin
            cosine_reg0 <= 36'sb111001011010111010001110110110000010;
            sine_reg0   <= 36'sb100000101011110000011111101000100000;
        end
        11749: begin
            cosine_reg0 <= 36'sb111001011011101011011011001110100011;
            sine_reg0   <= 36'sb100000101011100110001010110010100010;
        end
        11750: begin
            cosine_reg0 <= 36'sb111001011100011100100111110111010010;
            sine_reg0   <= 36'sb100000101011011011110111001001110110;
        end
        11751: begin
            cosine_reg0 <= 36'sb111001011101001101110100110000001100;
            sine_reg0   <= 36'sb100000101011010001100100101110011100;
        end
        11752: begin
            cosine_reg0 <= 36'sb111001011101111111000001111001001111;
            sine_reg0   <= 36'sb100000101011000111010011100000010101;
        end
        11753: begin
            cosine_reg0 <= 36'sb111001011110110000001111010010011001;
            sine_reg0   <= 36'sb100000101010111101000011011111100001;
        end
        11754: begin
            cosine_reg0 <= 36'sb111001011111100001011100111011101001;
            sine_reg0   <= 36'sb100000101010110010110100101100000000;
        end
        11755: begin
            cosine_reg0 <= 36'sb111001100000010010101010110100111101;
            sine_reg0   <= 36'sb100000101010101000100111000101110010;
        end
        11756: begin
            cosine_reg0 <= 36'sb111001100001000011111000111110010010;
            sine_reg0   <= 36'sb100000101010011110011010101100111001;
        end
        11757: begin
            cosine_reg0 <= 36'sb111001100001110101000111010111100111;
            sine_reg0   <= 36'sb100000101010010100001111100001010011;
        end
        11758: begin
            cosine_reg0 <= 36'sb111001100010100110010110000000111010;
            sine_reg0   <= 36'sb100000101010001010000101100011000011;
        end
        11759: begin
            cosine_reg0 <= 36'sb111001100011010111100100111010001001;
            sine_reg0   <= 36'sb100000101001111111111100110010001000;
        end
        11760: begin
            cosine_reg0 <= 36'sb111001100100001000110100000011010010;
            sine_reg0   <= 36'sb100000101001110101110101001110100011;
        end
        11761: begin
            cosine_reg0 <= 36'sb111001100100111010000011011100010100;
            sine_reg0   <= 36'sb100000101001101011101110111000010011;
        end
        11762: begin
            cosine_reg0 <= 36'sb111001100101101011010011000101001100;
            sine_reg0   <= 36'sb100000101001100001101001101111011010;
        end
        11763: begin
            cosine_reg0 <= 36'sb111001100110011100100010111101111000;
            sine_reg0   <= 36'sb100000101001010111100101110011111000;
        end
        11764: begin
            cosine_reg0 <= 36'sb111001100111001101110011000110010111;
            sine_reg0   <= 36'sb100000101001001101100011000101101101;
        end
        11765: begin
            cosine_reg0 <= 36'sb111001100111111111000011011110100110;
            sine_reg0   <= 36'sb100000101001000011100001100100111010;
        end
        11766: begin
            cosine_reg0 <= 36'sb111001101000110000010100000110100100;
            sine_reg0   <= 36'sb100000101000111001100001010001011110;
        end
        11767: begin
            cosine_reg0 <= 36'sb111001101001100001100100111110001111;
            sine_reg0   <= 36'sb100000101000101111100010001011011011;
        end
        11768: begin
            cosine_reg0 <= 36'sb111001101010010010110110000101100101;
            sine_reg0   <= 36'sb100000101000100101100100010010110000;
        end
        11769: begin
            cosine_reg0 <= 36'sb111001101011000100000111011100100100;
            sine_reg0   <= 36'sb100000101000011011100111100111011111;
        end
        11770: begin
            cosine_reg0 <= 36'sb111001101011110101011001000011001010;
            sine_reg0   <= 36'sb100000101000010001101100001001100111;
        end
        11771: begin
            cosine_reg0 <= 36'sb111001101100100110101010111001010101;
            sine_reg0   <= 36'sb100000101000000111110001111001001001;
        end
        11772: begin
            cosine_reg0 <= 36'sb111001101101010111111100111111000100;
            sine_reg0   <= 36'sb100000100111111101111000110110000101;
        end
        11773: begin
            cosine_reg0 <= 36'sb111001101110001001001111010100010100;
            sine_reg0   <= 36'sb100000100111110100000001000000011011;
        end
        11774: begin
            cosine_reg0 <= 36'sb111001101110111010100001111001000011;
            sine_reg0   <= 36'sb100000100111101010001010011000001101;
        end
        11775: begin
            cosine_reg0 <= 36'sb111001101111101011110100101101010001;
            sine_reg0   <= 36'sb100000100111100000010100111101011010;
        end
        11776: begin
            cosine_reg0 <= 36'sb111001110000011101000111110000111010;
            sine_reg0   <= 36'sb100000100111010110100000110000000011;
        end
        11777: begin
            cosine_reg0 <= 36'sb111001110001001110011011000011111100;
            sine_reg0   <= 36'sb100000100111001100101101110000001000;
        end
        11778: begin
            cosine_reg0 <= 36'sb111001110001111111101110100110010111;
            sine_reg0   <= 36'sb100000100111000010111011111101101010;
        end
        11779: begin
            cosine_reg0 <= 36'sb111001110010110001000010011000001000;
            sine_reg0   <= 36'sb100000100110111001001011011000101000;
        end
        11780: begin
            cosine_reg0 <= 36'sb111001110011100010010110011001001101;
            sine_reg0   <= 36'sb100000100110101111011100000001000100;
        end
        11781: begin
            cosine_reg0 <= 36'sb111001110100010011101010101001100100;
            sine_reg0   <= 36'sb100000100110100101101101110110111101;
        end
        11782: begin
            cosine_reg0 <= 36'sb111001110101000100111111001001001100;
            sine_reg0   <= 36'sb100000100110011100000000111010010101;
        end
        11783: begin
            cosine_reg0 <= 36'sb111001110101110110010011111000000001;
            sine_reg0   <= 36'sb100000100110010010010101001011001010;
        end
        11784: begin
            cosine_reg0 <= 36'sb111001110110100111101000110110000100;
            sine_reg0   <= 36'sb100000100110001000101010101001011111;
        end
        11785: begin
            cosine_reg0 <= 36'sb111001110111011000111110000011010001;
            sine_reg0   <= 36'sb100000100101111111000001010101010011;
        end
        11786: begin
            cosine_reg0 <= 36'sb111001111000001010010011011111100111;
            sine_reg0   <= 36'sb100000100101110101011001001110100110;
        end
        11787: begin
            cosine_reg0 <= 36'sb111001111000111011101001001011000011;
            sine_reg0   <= 36'sb100000100101101011110010010101011001;
        end
        11788: begin
            cosine_reg0 <= 36'sb111001111001101100111111000101100101;
            sine_reg0   <= 36'sb100000100101100010001100101001101100;
        end
        11789: begin
            cosine_reg0 <= 36'sb111001111010011110010101001111001010;
            sine_reg0   <= 36'sb100000100101011000101000001011100000;
        end
        11790: begin
            cosine_reg0 <= 36'sb111001111011001111101011100111101111;
            sine_reg0   <= 36'sb100000100101001111000100111010110101;
        end
        11791: begin
            cosine_reg0 <= 36'sb111001111100000001000010001111010100;
            sine_reg0   <= 36'sb100000100101000101100010110111101011;
        end
        11792: begin
            cosine_reg0 <= 36'sb111001111100110010011001000101110110;
            sine_reg0   <= 36'sb100000100100111100000010000010000100;
        end
        11793: begin
            cosine_reg0 <= 36'sb111001111101100011110000001011010100;
            sine_reg0   <= 36'sb100000100100110010100010011001111110;
        end
        11794: begin
            cosine_reg0 <= 36'sb111001111110010101000111011111101011;
            sine_reg0   <= 36'sb100000100100101001000011111111011010;
        end
        11795: begin
            cosine_reg0 <= 36'sb111001111111000110011111000010111010;
            sine_reg0   <= 36'sb100000100100011111100110110010011010;
        end
        11796: begin
            cosine_reg0 <= 36'sb111001111111110111110110110100111110;
            sine_reg0   <= 36'sb100000100100010110001010110010111100;
        end
        11797: begin
            cosine_reg0 <= 36'sb111010000000101001001110110101110111;
            sine_reg0   <= 36'sb100000100100001100110000000001000011;
        end
        11798: begin
            cosine_reg0 <= 36'sb111010000001011010100111000101100001;
            sine_reg0   <= 36'sb100000100100000011010110011100101101;
        end
        11799: begin
            cosine_reg0 <= 36'sb111010000010001011111111100011111011;
            sine_reg0   <= 36'sb100000100011111001111110000101111011;
        end
        11800: begin
            cosine_reg0 <= 36'sb111010000010111101011000010001000011;
            sine_reg0   <= 36'sb100000100011110000100110111100101110;
        end
        11801: begin
            cosine_reg0 <= 36'sb111010000011101110110001001100110111;
            sine_reg0   <= 36'sb100000100011100111010001000001000110;
        end
        11802: begin
            cosine_reg0 <= 36'sb111010000100100000001010010111010110;
            sine_reg0   <= 36'sb100000100011011101111100010011000100;
        end
        11803: begin
            cosine_reg0 <= 36'sb111010000101010001100011110000011101;
            sine_reg0   <= 36'sb100000100011010100101000110010100111;
        end
        11804: begin
            cosine_reg0 <= 36'sb111010000110000010111101011000001011;
            sine_reg0   <= 36'sb100000100011001011010110011111110000;
        end
        11805: begin
            cosine_reg0 <= 36'sb111010000110110100010111001110011101;
            sine_reg0   <= 36'sb100000100011000010000101011010100000;
        end
        11806: begin
            cosine_reg0 <= 36'sb111010000111100101110001010011010001;
            sine_reg0   <= 36'sb100000100010111000110101100010110110;
        end
        11807: begin
            cosine_reg0 <= 36'sb111010001000010111001011100110100111;
            sine_reg0   <= 36'sb100000100010101111100110111000110100;
        end
        11808: begin
            cosine_reg0 <= 36'sb111010001001001000100110001000011011;
            sine_reg0   <= 36'sb100000100010100110011001011100011001;
        end
        11809: begin
            cosine_reg0 <= 36'sb111010001001111010000000111000101100;
            sine_reg0   <= 36'sb100000100010011101001101001101100110;
        end
        11810: begin
            cosine_reg0 <= 36'sb111010001010101011011011110111011001;
            sine_reg0   <= 36'sb100000100010010100000010001100011011;
        end
        11811: begin
            cosine_reg0 <= 36'sb111010001011011100110111000100011110;
            sine_reg0   <= 36'sb100000100010001010111000011000111001;
        end
        11812: begin
            cosine_reg0 <= 36'sb111010001100001110010010011111111011;
            sine_reg0   <= 36'sb100000100010000001101111110010111111;
        end
        11813: begin
            cosine_reg0 <= 36'sb111010001100111111101110001001101101;
            sine_reg0   <= 36'sb100000100001111000101000011010101111;
        end
        11814: begin
            cosine_reg0 <= 36'sb111010001101110001001010000001110010;
            sine_reg0   <= 36'sb100000100001101111100010010000001001;
        end
        11815: begin
            cosine_reg0 <= 36'sb111010001110100010100110001000001001;
            sine_reg0   <= 36'sb100000100001100110011101010011001101;
        end
        11816: begin
            cosine_reg0 <= 36'sb111010001111010100000010011100110000;
            sine_reg0   <= 36'sb100000100001011101011001100011111010;
        end
        11817: begin
            cosine_reg0 <= 36'sb111010010000000101011110111111100100;
            sine_reg0   <= 36'sb100000100001010100010111000010010011;
        end
        11818: begin
            cosine_reg0 <= 36'sb111010010000110110111011110000100100;
            sine_reg0   <= 36'sb100000100001001011010101101110010111;
        end
        11819: begin
            cosine_reg0 <= 36'sb111010010001101000011000101111101110;
            sine_reg0   <= 36'sb100000100001000010010101101000000110;
        end
        11820: begin
            cosine_reg0 <= 36'sb111010010010011001110101111101000000;
            sine_reg0   <= 36'sb100000100000111001010110101111100000;
        end
        11821: begin
            cosine_reg0 <= 36'sb111010010011001011010011011000011000;
            sine_reg0   <= 36'sb100000100000110000011001000100100111;
        end
        11822: begin
            cosine_reg0 <= 36'sb111010010011111100110001000001110100;
            sine_reg0   <= 36'sb100000100000100111011100100111011010;
        end
        11823: begin
            cosine_reg0 <= 36'sb111010010100101110001110111001010010;
            sine_reg0   <= 36'sb100000100000011110100001010111111010;
        end
        11824: begin
            cosine_reg0 <= 36'sb111010010101011111101100111110110001;
            sine_reg0   <= 36'sb100000100000010101100111010110000111;
        end
        11825: begin
            cosine_reg0 <= 36'sb111010010110010001001011010010001110;
            sine_reg0   <= 36'sb100000100000001100101110100010000010;
        end
        11826: begin
            cosine_reg0 <= 36'sb111010010111000010101001110011101000;
            sine_reg0   <= 36'sb100000100000000011110110111011101010;
        end
        11827: begin
            cosine_reg0 <= 36'sb111010010111110100001000100010111100;
            sine_reg0   <= 36'sb100000011111111011000000100011000001;
        end
        11828: begin
            cosine_reg0 <= 36'sb111010011000100101100111100000001001;
            sine_reg0   <= 36'sb100000011111110010001011011000000110;
        end
        11829: begin
            cosine_reg0 <= 36'sb111010011001010111000110101011001101;
            sine_reg0   <= 36'sb100000011111101001010111011010111001;
        end
        11830: begin
            cosine_reg0 <= 36'sb111010011010001000100110000100000110;
            sine_reg0   <= 36'sb100000011111100000100100101011011100;
        end
        11831: begin
            cosine_reg0 <= 36'sb111010011010111010000101101010110001;
            sine_reg0   <= 36'sb100000011111010111110011001001101111;
        end
        11832: begin
            cosine_reg0 <= 36'sb111010011011101011100101011111001110;
            sine_reg0   <= 36'sb100000011111001111000010110101110001;
        end
        11833: begin
            cosine_reg0 <= 36'sb111010011100011101000101100001011010;
            sine_reg0   <= 36'sb100000011111000110010011101111100011;
        end
        11834: begin
            cosine_reg0 <= 36'sb111010011101001110100101110001010100;
            sine_reg0   <= 36'sb100000011110111101100101110111000110;
        end
        11835: begin
            cosine_reg0 <= 36'sb111010011110000000000110001110111000;
            sine_reg0   <= 36'sb100000011110110100111001001100011010;
        end
        11836: begin
            cosine_reg0 <= 36'sb111010011110110001100110111010000111;
            sine_reg0   <= 36'sb100000011110101100001101101111011111;
        end
        11837: begin
            cosine_reg0 <= 36'sb111010011111100011000111110010111100;
            sine_reg0   <= 36'sb100000011110100011100011100000010101;
        end
        11838: begin
            cosine_reg0 <= 36'sb111010100000010100101000111001011000;
            sine_reg0   <= 36'sb100000011110011010111010011110111101;
        end
        11839: begin
            cosine_reg0 <= 36'sb111010100001000110001010001101010111;
            sine_reg0   <= 36'sb100000011110010010010010101011011000;
        end
        11840: begin
            cosine_reg0 <= 36'sb111010100001110111101011101110110111;
            sine_reg0   <= 36'sb100000011110001001101100000101100101;
        end
        11841: begin
            cosine_reg0 <= 36'sb111010100010101001001101011101111000;
            sine_reg0   <= 36'sb100000011110000001000110101101100100;
        end
        11842: begin
            cosine_reg0 <= 36'sb111010100011011010101111011010010111;
            sine_reg0   <= 36'sb100000011101111000100010100011010111;
        end
        11843: begin
            cosine_reg0 <= 36'sb111010100100001100010001100100010010;
            sine_reg0   <= 36'sb100000011101101111111111100110111110;
        end
        11844: begin
            cosine_reg0 <= 36'sb111010100100111101110011111011100111;
            sine_reg0   <= 36'sb100000011101100111011101111000011000;
        end
        11845: begin
            cosine_reg0 <= 36'sb111010100101101111010110100000010100;
            sine_reg0   <= 36'sb100000011101011110111101010111100111;
        end
        11846: begin
            cosine_reg0 <= 36'sb111010100110100000111001010010011000;
            sine_reg0   <= 36'sb100000011101010110011110000100101010;
        end
        11847: begin
            cosine_reg0 <= 36'sb111010100111010010011100010001110000;
            sine_reg0   <= 36'sb100000011101001101111111111111100001;
        end
        11848: begin
            cosine_reg0 <= 36'sb111010101000000011111111011110011011;
            sine_reg0   <= 36'sb100000011101000101100011001000001110;
        end
        11849: begin
            cosine_reg0 <= 36'sb111010101000110101100010111000010110;
            sine_reg0   <= 36'sb100000011100111101000111011110110001;
        end
        11850: begin
            cosine_reg0 <= 36'sb111010101001100111000110011111100000;
            sine_reg0   <= 36'sb100000011100110100101101000011001001;
        end
        11851: begin
            cosine_reg0 <= 36'sb111010101010011000101010010011110111;
            sine_reg0   <= 36'sb100000011100101100010011110101010111;
        end
        11852: begin
            cosine_reg0 <= 36'sb111010101011001010001110010101011001;
            sine_reg0   <= 36'sb100000011100100011111011110101011100;
        end
        11853: begin
            cosine_reg0 <= 36'sb111010101011111011110010100100000100;
            sine_reg0   <= 36'sb100000011100011011100101000011010111;
        end
        11854: begin
            cosine_reg0 <= 36'sb111010101100101101010110111111110101;
            sine_reg0   <= 36'sb100000011100010011001111011111001010;
        end
        11855: begin
            cosine_reg0 <= 36'sb111010101101011110111011101000101100;
            sine_reg0   <= 36'sb100000011100001010111011001000110100;
        end
        11856: begin
            cosine_reg0 <= 36'sb111010101110010000100000011110100111;
            sine_reg0   <= 36'sb100000011100000010101000000000010101;
        end
        11857: begin
            cosine_reg0 <= 36'sb111010101111000010000101100001100010;
            sine_reg0   <= 36'sb100000011011111010010110000101101111;
        end
        11858: begin
            cosine_reg0 <= 36'sb111010101111110011101010110001011101;
            sine_reg0   <= 36'sb100000011011110010000101011001000001;
        end
        11859: begin
            cosine_reg0 <= 36'sb111010110000100101010000001110010110;
            sine_reg0   <= 36'sb100000011011101001110101111010001100;
        end
        11860: begin
            cosine_reg0 <= 36'sb111010110001010110110101111000001010;
            sine_reg0   <= 36'sb100000011011100001100111101001010000;
        end
        11861: begin
            cosine_reg0 <= 36'sb111010110010001000011011101110111000;
            sine_reg0   <= 36'sb100000011011011001011010100110001101;
        end
        11862: begin
            cosine_reg0 <= 36'sb111010110010111010000001110010011110;
            sine_reg0   <= 36'sb100000011011010001001110110001000100;
        end
        11863: begin
            cosine_reg0 <= 36'sb111010110011101011101000000010111001;
            sine_reg0   <= 36'sb100000011011001001000100001001110101;
        end
        11864: begin
            cosine_reg0 <= 36'sb111010110100011101001110100000001001;
            sine_reg0   <= 36'sb100000011011000000111010110000100000;
        end
        11865: begin
            cosine_reg0 <= 36'sb111010110101001110110101001010001010;
            sine_reg0   <= 36'sb100000011010111000110010100101000101;
        end
        11866: begin
            cosine_reg0 <= 36'sb111010110110000000011100000000111100;
            sine_reg0   <= 36'sb100000011010110000101011100111100110;
        end
        11867: begin
            cosine_reg0 <= 36'sb111010110110110010000011000100011100;
            sine_reg0   <= 36'sb100000011010101000100101111000000001;
        end
        11868: begin
            cosine_reg0 <= 36'sb111010110111100011101010010100101000;
            sine_reg0   <= 36'sb100000011010100000100001010110011001;
        end
        11869: begin
            cosine_reg0 <= 36'sb111010111000010101010001110001011110;
            sine_reg0   <= 36'sb100000011010011000011110000010101100;
        end
        11870: begin
            cosine_reg0 <= 36'sb111010111001000110111001011010111110;
            sine_reg0   <= 36'sb100000011010010000011011111100111011;
        end
        11871: begin
            cosine_reg0 <= 36'sb111010111001111000100001010001000011;
            sine_reg0   <= 36'sb100000011010001000011011000101000110;
        end
        11872: begin
            cosine_reg0 <= 36'sb111010111010101010001001010011101110;
            sine_reg0   <= 36'sb100000011010000000011011011011001111;
        end
        11873: begin
            cosine_reg0 <= 36'sb111010111011011011110001100010111011;
            sine_reg0   <= 36'sb100000011001111000011100111111010100;
        end
        11874: begin
            cosine_reg0 <= 36'sb111010111100001101011001111110101001;
            sine_reg0   <= 36'sb100000011001110000011111110001010111;
        end
        11875: begin
            cosine_reg0 <= 36'sb111010111100111111000010100110110101;
            sine_reg0   <= 36'sb100000011001101000100011110001011000;
        end
        11876: begin
            cosine_reg0 <= 36'sb111010111101110000101011011011011111;
            sine_reg0   <= 36'sb100000011001100000101000111111010110;
        end
        11877: begin
            cosine_reg0 <= 36'sb111010111110100010010100011100100100;
            sine_reg0   <= 36'sb100000011001011000101111011011010011;
        end
        11878: begin
            cosine_reg0 <= 36'sb111010111111010011111101101010000010;
            sine_reg0   <= 36'sb100000011001010000110111000101001110;
        end
        11879: begin
            cosine_reg0 <= 36'sb111011000000000101100111000011111000;
            sine_reg0   <= 36'sb100000011001001000111111111101001001;
        end
        11880: begin
            cosine_reg0 <= 36'sb111011000000110111010000101010000010;
            sine_reg0   <= 36'sb100000011001000001001010000011000010;
        end
        11881: begin
            cosine_reg0 <= 36'sb111011000001101000111010011100100001;
            sine_reg0   <= 36'sb100000011000111001010101010110111011;
        end
        11882: begin
            cosine_reg0 <= 36'sb111011000010011010100100011011010000;
            sine_reg0   <= 36'sb100000011000110001100001111000110100;
        end
        11883: begin
            cosine_reg0 <= 36'sb111011000011001100001110100110010000;
            sine_reg0   <= 36'sb100000011000101001101111101000101101;
        end
        11884: begin
            cosine_reg0 <= 36'sb111011000011111101111000111101011101;
            sine_reg0   <= 36'sb100000011000100001111110100110100110;
        end
        11885: begin
            cosine_reg0 <= 36'sb111011000100101111100011100000110101;
            sine_reg0   <= 36'sb100000011000011010001110110010100000;
        end
        11886: begin
            cosine_reg0 <= 36'sb111011000101100001001110010000011000;
            sine_reg0   <= 36'sb100000011000010010100000001100011011;
        end
        11887: begin
            cosine_reg0 <= 36'sb111011000110010010111001001100000011;
            sine_reg0   <= 36'sb100000011000001010110010110100011000;
        end
        11888: begin
            cosine_reg0 <= 36'sb111011000111000100100100010011110011;
            sine_reg0   <= 36'sb100000011000000011000110101010010110;
        end
        11889: begin
            cosine_reg0 <= 36'sb111011000111110110001111100111101000;
            sine_reg0   <= 36'sb100000010111111011011011101110010101;
        end
        11890: begin
            cosine_reg0 <= 36'sb111011001000100111111011000111011111;
            sine_reg0   <= 36'sb100000010111110011110010000000010111;
        end
        11891: begin
            cosine_reg0 <= 36'sb111011001001011001100110110011010110;
            sine_reg0   <= 36'sb100000010111101100001001100000011100;
        end
        11892: begin
            cosine_reg0 <= 36'sb111011001010001011010010101011001100;
            sine_reg0   <= 36'sb100000010111100100100010001110100011;
        end
        11893: begin
            cosine_reg0 <= 36'sb111011001010111100111110101110111110;
            sine_reg0   <= 36'sb100000010111011100111100001010101110;
        end
        11894: begin
            cosine_reg0 <= 36'sb111011001011101110101010111110101011;
            sine_reg0   <= 36'sb100000010111010101010111010100111100;
        end
        11895: begin
            cosine_reg0 <= 36'sb111011001100100000010111011010010000;
            sine_reg0   <= 36'sb100000010111001101110011101101001101;
        end
        11896: begin
            cosine_reg0 <= 36'sb111011001101010010000100000001101100;
            sine_reg0   <= 36'sb100000010111000110010001010011100010;
        end
        11897: begin
            cosine_reg0 <= 36'sb111011001110000011110000110100111101;
            sine_reg0   <= 36'sb100000010110111110110000000111111100;
        end
        11898: begin
            cosine_reg0 <= 36'sb111011001110110101011101110100000000;
            sine_reg0   <= 36'sb100000010110110111010000001010011010;
        end
        11899: begin
            cosine_reg0 <= 36'sb111011001111100111001010111110110101;
            sine_reg0   <= 36'sb100000010110101111110001011010111101;
        end
        11900: begin
            cosine_reg0 <= 36'sb111011010000011000111000010101011000;
            sine_reg0   <= 36'sb100000010110101000010011111001100101;
        end
        11901: begin
            cosine_reg0 <= 36'sb111011010001001010100101110111101001;
            sine_reg0   <= 36'sb100000010110100000110111100110010011;
        end
        11902: begin
            cosine_reg0 <= 36'sb111011010001111100010011100101100101;
            sine_reg0   <= 36'sb100000010110011001011100100001000110;
        end
        11903: begin
            cosine_reg0 <= 36'sb111011010010101110000001011111001011;
            sine_reg0   <= 36'sb100000010110010010000010101001111111;
        end
        11904: begin
            cosine_reg0 <= 36'sb111011010011011111101111100100010111;
            sine_reg0   <= 36'sb100000010110001010101010000000111111;
        end
        11905: begin
            cosine_reg0 <= 36'sb111011010100010001011101110101001001;
            sine_reg0   <= 36'sb100000010110000011010010100110000101;
        end
        11906: begin
            cosine_reg0 <= 36'sb111011010101000011001100010001011111;
            sine_reg0   <= 36'sb100000010101111011111100011001010010;
        end
        11907: begin
            cosine_reg0 <= 36'sb111011010101110100111010111001010110;
            sine_reg0   <= 36'sb100000010101110100100111011010100110;
        end
        11908: begin
            cosine_reg0 <= 36'sb111011010110100110101001101100101101;
            sine_reg0   <= 36'sb100000010101101101010011101010000001;
        end
        11909: begin
            cosine_reg0 <= 36'sb111011010111011000011000101011100010;
            sine_reg0   <= 36'sb100000010101100110000001000111100100;
        end
        11910: begin
            cosine_reg0 <= 36'sb111011011000001010000111110101110011;
            sine_reg0   <= 36'sb100000010101011110101111110011001111;
        end
        11911: begin
            cosine_reg0 <= 36'sb111011011000111011110111001011011110;
            sine_reg0   <= 36'sb100000010101010111011111101101000010;
        end
        11912: begin
            cosine_reg0 <= 36'sb111011011001101101100110101100100000;
            sine_reg0   <= 36'sb100000010101010000010000110100111110;
        end
        11913: begin
            cosine_reg0 <= 36'sb111011011010011111010110011000111001;
            sine_reg0   <= 36'sb100000010101001001000011001011000010;
        end
        11914: begin
            cosine_reg0 <= 36'sb111011011011010001000110010000100110;
            sine_reg0   <= 36'sb100000010101000001110110101111010000;
        end
        11915: begin
            cosine_reg0 <= 36'sb111011011100000010110110010011100110;
            sine_reg0   <= 36'sb100000010100111010101011100001100111;
        end
        11916: begin
            cosine_reg0 <= 36'sb111011011100110100100110100001110101;
            sine_reg0   <= 36'sb100000010100110011100001100010000111;
        end
        11917: begin
            cosine_reg0 <= 36'sb111011011101100110010110111011010011;
            sine_reg0   <= 36'sb100000010100101100011000110000110010;
        end
        11918: begin
            cosine_reg0 <= 36'sb111011011110011000000111011111111110;
            sine_reg0   <= 36'sb100000010100100101010001001101100110;
        end
        11919: begin
            cosine_reg0 <= 36'sb111011011111001001111000001111110011;
            sine_reg0   <= 36'sb100000010100011110001010111000100101;
        end
        11920: begin
            cosine_reg0 <= 36'sb111011011111111011101001001010110001;
            sine_reg0   <= 36'sb100000010100010111000101110001101111;
        end
        11921: begin
            cosine_reg0 <= 36'sb111011100000101101011010010000110110;
            sine_reg0   <= 36'sb100000010100010000000001111001000100;
        end
        11922: begin
            cosine_reg0 <= 36'sb111011100001011111001011100010000000;
            sine_reg0   <= 36'sb100000010100001000111111001110100100;
        end
        11923: begin
            cosine_reg0 <= 36'sb111011100010010000111100111110001100;
            sine_reg0   <= 36'sb100000010100000001111101110010010000;
        end
        11924: begin
            cosine_reg0 <= 36'sb111011100011000010101110100101011010;
            sine_reg0   <= 36'sb100000010011111010111101100100000111;
        end
        11925: begin
            cosine_reg0 <= 36'sb111011100011110100100000010111100111;
            sine_reg0   <= 36'sb100000010011110011111110100100001011;
        end
        11926: begin
            cosine_reg0 <= 36'sb111011100100100110010010010100110001;
            sine_reg0   <= 36'sb100000010011101101000000110010011011;
        end
        11927: begin
            cosine_reg0 <= 36'sb111011100101011000000100011100110110;
            sine_reg0   <= 36'sb100000010011100110000100001110110111;
        end
        11928: begin
            cosine_reg0 <= 36'sb111011100110001001110110101111110100;
            sine_reg0   <= 36'sb100000010011011111001000111001100001;
        end
        11929: begin
            cosine_reg0 <= 36'sb111011100110111011101001001101101010;
            sine_reg0   <= 36'sb100000010011011000001110110010010111;
        end
        11930: begin
            cosine_reg0 <= 36'sb111011100111101101011011110110010110;
            sine_reg0   <= 36'sb100000010011010001010101111001011011;
        end
        11931: begin
            cosine_reg0 <= 36'sb111011101000011111001110101001110101;
            sine_reg0   <= 36'sb100000010011001010011110001110101101;
        end
        11932: begin
            cosine_reg0 <= 36'sb111011101001010001000001101000000101;
            sine_reg0   <= 36'sb100000010011000011100111110010001100;
        end
        11933: begin
            cosine_reg0 <= 36'sb111011101010000010110100110001000110;
            sine_reg0   <= 36'sb100000010010111100110010100011111010;
        end
        11934: begin
            cosine_reg0 <= 36'sb111011101010110100101000000100110100;
            sine_reg0   <= 36'sb100000010010110101111110100011110110;
        end
        11935: begin
            cosine_reg0 <= 36'sb111011101011100110011011100011001110;
            sine_reg0   <= 36'sb100000010010101111001011110010000001;
        end
        11936: begin
            cosine_reg0 <= 36'sb111011101100011000001111001100010010;
            sine_reg0   <= 36'sb100000010010101000011010001110011100;
        end
        11937: begin
            cosine_reg0 <= 36'sb111011101101001010000010111111111111;
            sine_reg0   <= 36'sb100000010010100001101001111001000101;
        end
        11938: begin
            cosine_reg0 <= 36'sb111011101101111011110110111110010001;
            sine_reg0   <= 36'sb100000010010011010111010110001111110;
        end
        11939: begin
            cosine_reg0 <= 36'sb111011101110101101101011000111001000;
            sine_reg0   <= 36'sb100000010010010100001100111001000110;
        end
        11940: begin
            cosine_reg0 <= 36'sb111011101111011111011111011010100001;
            sine_reg0   <= 36'sb100000010010001101100000001110011111;
        end
        11941: begin
            cosine_reg0 <= 36'sb111011110000010001010011111000011010;
            sine_reg0   <= 36'sb100000010010000110110100110010001000;
        end
        11942: begin
            cosine_reg0 <= 36'sb111011110001000011001000100000110010;
            sine_reg0   <= 36'sb100000010010000000001010100100000010;
        end
        11943: begin
            cosine_reg0 <= 36'sb111011110001110100111101010011100110;
            sine_reg0   <= 36'sb100000010001111001100001100100001100;
        end
        11944: begin
            cosine_reg0 <= 36'sb111011110010100110110010010000110101;
            sine_reg0   <= 36'sb100000010001110010111001110010100111;
        end
        11945: begin
            cosine_reg0 <= 36'sb111011110011011000100111011000011101;
            sine_reg0   <= 36'sb100000010001101100010011001111010100;
        end
        11946: begin
            cosine_reg0 <= 36'sb111011110100001010011100101010011011;
            sine_reg0   <= 36'sb100000010001100101101101111010010010;
        end
        11947: begin
            cosine_reg0 <= 36'sb111011110100111100010010000110101110;
            sine_reg0   <= 36'sb100000010001011111001001110011100011;
        end
        11948: begin
            cosine_reg0 <= 36'sb111011110101101110000111101101010101;
            sine_reg0   <= 36'sb100000010001011000100110111011000101;
        end
        11949: begin
            cosine_reg0 <= 36'sb111011110110011111111101011110001100;
            sine_reg0   <= 36'sb100000010001010010000101010000111010;
        end
        11950: begin
            cosine_reg0 <= 36'sb111011110111010001110011011001010010;
            sine_reg0   <= 36'sb100000010001001011100100110101000001;
        end
        11951: begin
            cosine_reg0 <= 36'sb111011111000000011101001011110100110;
            sine_reg0   <= 36'sb100000010001000101000101100111011011;
        end
        11952: begin
            cosine_reg0 <= 36'sb111011111000110101011111101110000100;
            sine_reg0   <= 36'sb100000010000111110100111101000001000;
        end
        11953: begin
            cosine_reg0 <= 36'sb111011111001100111010110000111101101;
            sine_reg0   <= 36'sb100000010000111000001010110111001000;
        end
        11954: begin
            cosine_reg0 <= 36'sb111011111010011001001100101011011100;
            sine_reg0   <= 36'sb100000010000110001101111010100011101;
        end
        11955: begin
            cosine_reg0 <= 36'sb111011111011001011000011011001010001;
            sine_reg0   <= 36'sb100000010000101011010101000000000100;
        end
        11956: begin
            cosine_reg0 <= 36'sb111011111011111100111010010001001010;
            sine_reg0   <= 36'sb100000010000100100111011111010000000;
        end
        11957: begin
            cosine_reg0 <= 36'sb111011111100101110110001010011000100;
            sine_reg0   <= 36'sb100000010000011110100100000010010001;
        end
        11958: begin
            cosine_reg0 <= 36'sb111011111101100000101000011110111110;
            sine_reg0   <= 36'sb100000010000011000001101011000110110;
        end
        11959: begin
            cosine_reg0 <= 36'sb111011111110010010011111110100110110;
            sine_reg0   <= 36'sb100000010000010001110111111101110000;
        end
        11960: begin
            cosine_reg0 <= 36'sb111011111111000100010111010100101001;
            sine_reg0   <= 36'sb100000010000001011100011110000111110;
        end
        11961: begin
            cosine_reg0 <= 36'sb111011111111110110001110111110010111;
            sine_reg0   <= 36'sb100000010000000101010000110010100010;
        end
        11962: begin
            cosine_reg0 <= 36'sb111100000000101000000110110001111100;
            sine_reg0   <= 36'sb100000001111111110111111000010011100;
        end
        11963: begin
            cosine_reg0 <= 36'sb111100000001011001111110101111011000;
            sine_reg0   <= 36'sb100000001111111000101110100000101100;
        end
        11964: begin
            cosine_reg0 <= 36'sb111100000010001011110110110110101000;
            sine_reg0   <= 36'sb100000001111110010011111001101010001;
        end
        11965: begin
            cosine_reg0 <= 36'sb111100000010111101101111000111101010;
            sine_reg0   <= 36'sb100000001111101100010001001000001101;
        end
        11966: begin
            cosine_reg0 <= 36'sb111100000011101111100111100010011101;
            sine_reg0   <= 36'sb100000001111100110000100010001011111;
        end
        11967: begin
            cosine_reg0 <= 36'sb111100000100100001100000000110111101;
            sine_reg0   <= 36'sb100000001111011111111000101001001000;
        end
        11968: begin
            cosine_reg0 <= 36'sb111100000101010011011000110101001011;
            sine_reg0   <= 36'sb100000001111011001101110001111001001;
        end
        11969: begin
            cosine_reg0 <= 36'sb111100000110000101010001101101000011;
            sine_reg0   <= 36'sb100000001111010011100101000011100000;
        end
        11970: begin
            cosine_reg0 <= 36'sb111100000110110111001010101110100011;
            sine_reg0   <= 36'sb100000001111001101011101000110001111;
        end
        11971: begin
            cosine_reg0 <= 36'sb111100000111101001000011111001101011;
            sine_reg0   <= 36'sb100000001111000111010110010111010101;
        end
        11972: begin
            cosine_reg0 <= 36'sb111100001000011010111101001110010111;
            sine_reg0   <= 36'sb100000001111000001010000110110110100;
        end
        11973: begin
            cosine_reg0 <= 36'sb111100001001001100110110101100100110;
            sine_reg0   <= 36'sb100000001110111011001100100100101010;
        end
        11974: begin
            cosine_reg0 <= 36'sb111100001001111110110000010100010110;
            sine_reg0   <= 36'sb100000001110110101001001100000111001;
        end
        11975: begin
            cosine_reg0 <= 36'sb111100001010110000101010000101100101;
            sine_reg0   <= 36'sb100000001110101111000111101011100001;
        end
        11976: begin
            cosine_reg0 <= 36'sb111100001011100010100100000000010001;
            sine_reg0   <= 36'sb100000001110101001000111000100100010;
        end
        11977: begin
            cosine_reg0 <= 36'sb111100001100010100011110000100011000;
            sine_reg0   <= 36'sb100000001110100011000111101011111011;
        end
        11978: begin
            cosine_reg0 <= 36'sb111100001101000110011000010001111001;
            sine_reg0   <= 36'sb100000001110011101001001100001101110;
        end
        11979: begin
            cosine_reg0 <= 36'sb111100001101111000010010101000110001;
            sine_reg0   <= 36'sb100000001110010111001100100101111011;
        end
        11980: begin
            cosine_reg0 <= 36'sb111100001110101010001101001000111110;
            sine_reg0   <= 36'sb100000001110010001010000111000100001;
        end
        11981: begin
            cosine_reg0 <= 36'sb111100001111011100000111110010011111;
            sine_reg0   <= 36'sb100000001110001011010110011001100010;
        end
        11982: begin
            cosine_reg0 <= 36'sb111100010000001110000010100101010001;
            sine_reg0   <= 36'sb100000001110000101011101001000111100;
        end
        11983: begin
            cosine_reg0 <= 36'sb111100010000111111111101100001010011;
            sine_reg0   <= 36'sb100000001101111111100101000110110001;
        end
        11984: begin
            cosine_reg0 <= 36'sb111100010001110001111000100110100011;
            sine_reg0   <= 36'sb100000001101111001101110010011000001;
        end
        11985: begin
            cosine_reg0 <= 36'sb111100010010100011110011110100111110;
            sine_reg0   <= 36'sb100000001101110011111000101101101100;
        end
        11986: begin
            cosine_reg0 <= 36'sb111100010011010101101111001100100011;
            sine_reg0   <= 36'sb100000001101101110000100010110110010;
        end
        11987: begin
            cosine_reg0 <= 36'sb111100010100000111101010101101010001;
            sine_reg0   <= 36'sb100000001101101000010001001110010011;
        end
        11988: begin
            cosine_reg0 <= 36'sb111100010100111001100110010111000100;
            sine_reg0   <= 36'sb100000001101100010011111010100010000;
        end
        11989: begin
            cosine_reg0 <= 36'sb111100010101101011100010001001111011;
            sine_reg0   <= 36'sb100000001101011100101110101000101001;
        end
        11990: begin
            cosine_reg0 <= 36'sb111100010110011101011110000101110101;
            sine_reg0   <= 36'sb100000001101010110111111001011011110;
        end
        11991: begin
            cosine_reg0 <= 36'sb111100010111001111011010001010101111;
            sine_reg0   <= 36'sb100000001101010001010000111100101111;
        end
        11992: begin
            cosine_reg0 <= 36'sb111100011000000001010110011000100111;
            sine_reg0   <= 36'sb100000001101001011100011111100011101;
        end
        11993: begin
            cosine_reg0 <= 36'sb111100011000110011010010101111011011;
            sine_reg0   <= 36'sb100000001101000101111000001010100111;
        end
        11994: begin
            cosine_reg0 <= 36'sb111100011001100101001111001111001010;
            sine_reg0   <= 36'sb100000001101000000001101100111001110;
        end
        11995: begin
            cosine_reg0 <= 36'sb111100011010010111001011110111110001;
            sine_reg0   <= 36'sb100000001100111010100100010010010011;
        end
        11996: begin
            cosine_reg0 <= 36'sb111100011011001001001000101001001111;
            sine_reg0   <= 36'sb100000001100110100111100001011110100;
        end
        11997: begin
            cosine_reg0 <= 36'sb111100011011111011000101100011100010;
            sine_reg0   <= 36'sb100000001100101111010101010011110100;
        end
        11998: begin
            cosine_reg0 <= 36'sb111100011100101101000010100110101000;
            sine_reg0   <= 36'sb100000001100101001101111101010010001;
        end
        11999: begin
            cosine_reg0 <= 36'sb111100011101011110111111110010011110;
            sine_reg0   <= 36'sb100000001100100100001011001111001100;
        end
        12000: begin
            cosine_reg0 <= 36'sb111100011110010000111101000111000011;
            sine_reg0   <= 36'sb100000001100011110101000000010100110;
        end
        12001: begin
            cosine_reg0 <= 36'sb111100011111000010111010100100010101;
            sine_reg0   <= 36'sb100000001100011001000110000100011101;
        end
        12002: begin
            cosine_reg0 <= 36'sb111100011111110100111000001010010011;
            sine_reg0   <= 36'sb100000001100010011100101010100110100;
        end
        12003: begin
            cosine_reg0 <= 36'sb111100100000100110110101111000111001;
            sine_reg0   <= 36'sb100000001100001110000101110011101001;
        end
        12004: begin
            cosine_reg0 <= 36'sb111100100001011000110011110000000111;
            sine_reg0   <= 36'sb100000001100001000100111100000111110;
        end
        12005: begin
            cosine_reg0 <= 36'sb111100100010001010110001101111111001;
            sine_reg0   <= 36'sb100000001100000011001010011100110010;
        end
        12006: begin
            cosine_reg0 <= 36'sb111100100010111100101111111000010000;
            sine_reg0   <= 36'sb100000001011111101101110100111000101;
        end
        12007: begin
            cosine_reg0 <= 36'sb111100100011101110101110001001000111;
            sine_reg0   <= 36'sb100000001011111000010011111111111000;
        end
        12008: begin
            cosine_reg0 <= 36'sb111100100100100000101100100010011110;
            sine_reg0   <= 36'sb100000001011110010111010100111001011;
        end
        12009: begin
            cosine_reg0 <= 36'sb111100100101010010101011000100010011;
            sine_reg0   <= 36'sb100000001011101101100010011100111110;
        end
        12010: begin
            cosine_reg0 <= 36'sb111100100110000100101001101110100011;
            sine_reg0   <= 36'sb100000001011101000001011100001010001;
        end
        12011: begin
            cosine_reg0 <= 36'sb111100100110110110101000100001001101;
            sine_reg0   <= 36'sb100000001011100010110101110100000101;
        end
        12012: begin
            cosine_reg0 <= 36'sb111100100111101000100111011100001111;
            sine_reg0   <= 36'sb100000001011011101100001010101011010;
        end
        12013: begin
            cosine_reg0 <= 36'sb111100101000011010100110011111100111;
            sine_reg0   <= 36'sb100000001011011000001110000101010000;
        end
        12014: begin
            cosine_reg0 <= 36'sb111100101001001100100101101011010010;
            sine_reg0   <= 36'sb100000001011010010111100000011100111;
        end
        12015: begin
            cosine_reg0 <= 36'sb111100101001111110100100111111010000;
            sine_reg0   <= 36'sb100000001011001101101011010000011111;
        end
        12016: begin
            cosine_reg0 <= 36'sb111100101010110000100100011011011110;
            sine_reg0   <= 36'sb100000001011001000011011101011111000;
        end
        12017: begin
            cosine_reg0 <= 36'sb111100101011100010100011111111111010;
            sine_reg0   <= 36'sb100000001011000011001101010101110100;
        end
        12018: begin
            cosine_reg0 <= 36'sb111100101100010100100011101100100010;
            sine_reg0   <= 36'sb100000001010111110000000001110010010;
        end
        12019: begin
            cosine_reg0 <= 36'sb111100101101000110100011100001010100;
            sine_reg0   <= 36'sb100000001010111000110100010101010001;
        end
        12020: begin
            cosine_reg0 <= 36'sb111100101101111000100011011110001111;
            sine_reg0   <= 36'sb100000001010110011101001101010110011;
        end
        12021: begin
            cosine_reg0 <= 36'sb111100101110101010100011100011010000;
            sine_reg0   <= 36'sb100000001010101110100000001110111000;
        end
        12022: begin
            cosine_reg0 <= 36'sb111100101111011100100011110000010110;
            sine_reg0   <= 36'sb100000001010101001011000000001011111;
        end
        12023: begin
            cosine_reg0 <= 36'sb111100110000001110100100000101011110;
            sine_reg0   <= 36'sb100000001010100100010001000010101010;
        end
        12024: begin
            cosine_reg0 <= 36'sb111100110001000000100100100010100111;
            sine_reg0   <= 36'sb100000001010011111001011010010010111;
        end
        12025: begin
            cosine_reg0 <= 36'sb111100110001110010100101000111101111;
            sine_reg0   <= 36'sb100000001010011010000110110000101000;
        end
        12026: begin
            cosine_reg0 <= 36'sb111100110010100100100101110100110011;
            sine_reg0   <= 36'sb100000001010010101000011011101011100;
        end
        12027: begin
            cosine_reg0 <= 36'sb111100110011010110100110101001110010;
            sine_reg0   <= 36'sb100000001010010000000001011000110101;
        end
        12028: begin
            cosine_reg0 <= 36'sb111100110100001000100111100110101011;
            sine_reg0   <= 36'sb100000001010001011000000100010110001;
        end
        12029: begin
            cosine_reg0 <= 36'sb111100110100111010101000101011011010;
            sine_reg0   <= 36'sb100000001010000110000000111011010001;
        end
        12030: begin
            cosine_reg0 <= 36'sb111100110101101100101001110111111110;
            sine_reg0   <= 36'sb100000001010000001000010100010010110;
        end
        12031: begin
            cosine_reg0 <= 36'sb111100110110011110101011001100010110;
            sine_reg0   <= 36'sb100000001001111100000101010111111111;
        end
        12032: begin
            cosine_reg0 <= 36'sb111100110111010000101100101000011111;
            sine_reg0   <= 36'sb100000001001110111001001011100001101;
        end
        12033: begin
            cosine_reg0 <= 36'sb111100111000000010101110001100010111;
            sine_reg0   <= 36'sb100000001001110010001110101110111111;
        end
        12034: begin
            cosine_reg0 <= 36'sb111100111000110100101111110111111100;
            sine_reg0   <= 36'sb100000001001101101010101010000010111;
        end
        12035: begin
            cosine_reg0 <= 36'sb111100111001100110110001101011001101;
            sine_reg0   <= 36'sb100000001001101000011101000000010100;
        end
        12036: begin
            cosine_reg0 <= 36'sb111100111010011000110011100110001000;
            sine_reg0   <= 36'sb100000001001100011100101111110110111;
        end
        12037: begin
            cosine_reg0 <= 36'sb111100111011001010110101101000101010;
            sine_reg0   <= 36'sb100000001001011110110000001011111111;
        end
        12038: begin
            cosine_reg0 <= 36'sb111100111011111100110111110010110001;
            sine_reg0   <= 36'sb100000001001011001111011100111101101;
        end
        12039: begin
            cosine_reg0 <= 36'sb111100111100101110111010000100011101;
            sine_reg0   <= 36'sb100000001001010101001000010010000010;
        end
        12040: begin
            cosine_reg0 <= 36'sb111100111101100000111100011101101010;
            sine_reg0   <= 36'sb100000001001010000010110001010111100;
        end
        12041: begin
            cosine_reg0 <= 36'sb111100111110010010111110111110010111;
            sine_reg0   <= 36'sb100000001001001011100101010010011101;
        end
        12042: begin
            cosine_reg0 <= 36'sb111100111111000101000001100110100010;
            sine_reg0   <= 36'sb100000001001000110110101101000100100;
        end
        12043: begin
            cosine_reg0 <= 36'sb111100111111110111000100010110001001;
            sine_reg0   <= 36'sb100000001001000010000111001101010010;
        end
        12044: begin
            cosine_reg0 <= 36'sb111101000000101001000111001101001010;
            sine_reg0   <= 36'sb100000001000111101011010000000100111;
        end
        12045: begin
            cosine_reg0 <= 36'sb111101000001011011001010001011100100;
            sine_reg0   <= 36'sb100000001000111000101110000010100011;
        end
        12046: begin
            cosine_reg0 <= 36'sb111101000010001101001101010001010011;
            sine_reg0   <= 36'sb100000001000110100000011010011000111;
        end
        12047: begin
            cosine_reg0 <= 36'sb111101000010111111010000011110010111;
            sine_reg0   <= 36'sb100000001000101111011001110010010010;
        end
        12048: begin
            cosine_reg0 <= 36'sb111101000011110001010011110010101101;
            sine_reg0   <= 36'sb100000001000101010110001100000000101;
        end
        12049: begin
            cosine_reg0 <= 36'sb111101000100100011010111001110010100;
            sine_reg0   <= 36'sb100000001000100110001010011100011111;
        end
        12050: begin
            cosine_reg0 <= 36'sb111101000101010101011010110001001001;
            sine_reg0   <= 36'sb100000001000100001100100100111100010;
        end
        12051: begin
            cosine_reg0 <= 36'sb111101000110000111011110011011001011;
            sine_reg0   <= 36'sb100000001000011101000000000001001100;
        end
        12052: begin
            cosine_reg0 <= 36'sb111101000110111001100010001100010111;
            sine_reg0   <= 36'sb100000001000011000011100101001011111;
        end
        12053: begin
            cosine_reg0 <= 36'sb111101000111101011100110000100101100;
            sine_reg0   <= 36'sb100000001000010011111010100000011011;
        end
        12054: begin
            cosine_reg0 <= 36'sb111101001000011101101010000100001000;
            sine_reg0   <= 36'sb100000001000001111011001100101111111;
        end
        12055: begin
            cosine_reg0 <= 36'sb111101001001001111101110001010101001;
            sine_reg0   <= 36'sb100000001000001010111001111010001101;
        end
        12056: begin
            cosine_reg0 <= 36'sb111101001010000001110010011000001100;
            sine_reg0   <= 36'sb100000001000000110011011011101000011;
        end
        12057: begin
            cosine_reg0 <= 36'sb111101001010110011110110101100110001;
            sine_reg0   <= 36'sb100000001000000001111110001110100011;
        end
        12058: begin
            cosine_reg0 <= 36'sb111101001011100101111011001000010101;
            sine_reg0   <= 36'sb100000000111111101100010001110101100;
        end
        12059: begin
            cosine_reg0 <= 36'sb111101001100010111111111101010110101;
            sine_reg0   <= 36'sb100000000111111001000111011101011111;
        end
        12060: begin
            cosine_reg0 <= 36'sb111101001101001010000100010100010010;
            sine_reg0   <= 36'sb100000000111110100101101111010111011;
        end
        12061: begin
            cosine_reg0 <= 36'sb111101001101111100001001000100100111;
            sine_reg0   <= 36'sb100000000111110000010101100111000001;
        end
        12062: begin
            cosine_reg0 <= 36'sb111101001110101110001101111011110100;
            sine_reg0   <= 36'sb100000000111101011111110100001110010;
        end
        12063: begin
            cosine_reg0 <= 36'sb111101001111100000010010111001110110;
            sine_reg0   <= 36'sb100000000111100111101000101011001100;
        end
        12064: begin
            cosine_reg0 <= 36'sb111101010000010010010111111110101011;
            sine_reg0   <= 36'sb100000000111100011010100000011010010;
        end
        12065: begin
            cosine_reg0 <= 36'sb111101010001000100011101001010010010;
            sine_reg0   <= 36'sb100000000111011111000000101010000001;
        end
        12066: begin
            cosine_reg0 <= 36'sb111101010001110110100010011100101001;
            sine_reg0   <= 36'sb100000000111011010101110011111011100;
        end
        12067: begin
            cosine_reg0 <= 36'sb111101010010101000100111110101101110;
            sine_reg0   <= 36'sb100000000111010110011101100011100001;
        end
        12068: begin
            cosine_reg0 <= 36'sb111101010011011010101101010101011110;
            sine_reg0   <= 36'sb100000000111010010001101110110010010;
        end
        12069: begin
            cosine_reg0 <= 36'sb111101010100001100110010111011111000;
            sine_reg0   <= 36'sb100000000111001101111111010111101110;
        end
        12070: begin
            cosine_reg0 <= 36'sb111101010100111110111000101000111010;
            sine_reg0   <= 36'sb100000000111001001110010000111110101;
        end
        12071: begin
            cosine_reg0 <= 36'sb111101010101110000111110011100100010;
            sine_reg0   <= 36'sb100000000111000101100110000110101000;
        end
        12072: begin
            cosine_reg0 <= 36'sb111101010110100011000100010110101110;
            sine_reg0   <= 36'sb100000000111000001011011010100000111;
        end
        12073: begin
            cosine_reg0 <= 36'sb111101010111010101001010010111011100;
            sine_reg0   <= 36'sb100000000110111101010001110000010001;
        end
        12074: begin
            cosine_reg0 <= 36'sb111101011000000111010000011110101010;
            sine_reg0   <= 36'sb100000000110111001001001011011001000;
        end
        12075: begin
            cosine_reg0 <= 36'sb111101011000111001010110101100010110;
            sine_reg0   <= 36'sb100000000110110101000010010100101010;
        end
        12076: begin
            cosine_reg0 <= 36'sb111101011001101011011101000000011111;
            sine_reg0   <= 36'sb100000000110110000111100011100111010;
        end
        12077: begin
            cosine_reg0 <= 36'sb111101011010011101100011011011000010;
            sine_reg0   <= 36'sb100000000110101100110111110011110101;
        end
        12078: begin
            cosine_reg0 <= 36'sb111101011011001111101001111011111110;
            sine_reg0   <= 36'sb100000000110101000110100011001011110;
        end
        12079: begin
            cosine_reg0 <= 36'sb111101011100000001110000100011010000;
            sine_reg0   <= 36'sb100000000110100100110010001101110011;
        end
        12080: begin
            cosine_reg0 <= 36'sb111101011100110011110111010000110111;
            sine_reg0   <= 36'sb100000000110100000110001010000110101;
        end
        12081: begin
            cosine_reg0 <= 36'sb111101011101100101111110000100110000;
            sine_reg0   <= 36'sb100000000110011100110001100010100101;
        end
        12082: begin
            cosine_reg0 <= 36'sb111101011110011000000100111110111010;
            sine_reg0   <= 36'sb100000000110011000110011000011000010;
        end
        12083: begin
            cosine_reg0 <= 36'sb111101011111001010001011111111010011;
            sine_reg0   <= 36'sb100000000110010100110101110010001100;
        end
        12084: begin
            cosine_reg0 <= 36'sb111101011111111100010011000101111001;
            sine_reg0   <= 36'sb100000000110010000111001110000000100;
        end
        12085: begin
            cosine_reg0 <= 36'sb111101100000101110011010010010101010;
            sine_reg0   <= 36'sb100000000110001100111110111100101010;
        end
        12086: begin
            cosine_reg0 <= 36'sb111101100001100000100001100101100011;
            sine_reg0   <= 36'sb100000000110001001000101010111111101;
        end
        12087: begin
            cosine_reg0 <= 36'sb111101100010010010101000111110100100;
            sine_reg0   <= 36'sb100000000110000101001101000001111111;
        end
        12088: begin
            cosine_reg0 <= 36'sb111101100011000100110000011101101010;
            sine_reg0   <= 36'sb100000000110000001010101111010101111;
        end
        12089: begin
            cosine_reg0 <= 36'sb111101100011110110111000000010110011;
            sine_reg0   <= 36'sb100000000101111101100000000010001101;
        end
        12090: begin
            cosine_reg0 <= 36'sb111101100100101000111111101101111101;
            sine_reg0   <= 36'sb100000000101111001101011011000011010;
        end
        12091: begin
            cosine_reg0 <= 36'sb111101100101011011000111011111000111;
            sine_reg0   <= 36'sb100000000101110101110111111101010110;
        end
        12092: begin
            cosine_reg0 <= 36'sb111101100110001101001111010110001110;
            sine_reg0   <= 36'sb100000000101110010000101110001000000;
        end
        12093: begin
            cosine_reg0 <= 36'sb111101100110111111010111010011010001;
            sine_reg0   <= 36'sb100000000101101110010100110011011001;
        end
        12094: begin
            cosine_reg0 <= 36'sb111101100111110001011111010110001101;
            sine_reg0   <= 36'sb100000000101101010100101000100100010;
        end
        12095: begin
            cosine_reg0 <= 36'sb111101101000100011100111011111000000;
            sine_reg0   <= 36'sb100000000101100110110110100100011010;
        end
        12096: begin
            cosine_reg0 <= 36'sb111101101001010101101111101101101010;
            sine_reg0   <= 36'sb100000000101100011001001010011000001;
        end
        12097: begin
            cosine_reg0 <= 36'sb111101101010000111111000000010000111;
            sine_reg0   <= 36'sb100000000101011111011101010000010111;
        end
        12098: begin
            cosine_reg0 <= 36'sb111101101010111010000000011100010110;
            sine_reg0   <= 36'sb100000000101011011110010011100011110;
        end
        12099: begin
            cosine_reg0 <= 36'sb111101101011101100001000111100010100;
            sine_reg0   <= 36'sb100000000101011000001000110111010100;
        end
        12100: begin
            cosine_reg0 <= 36'sb111101101100011110010001100010000001;
            sine_reg0   <= 36'sb100000000101010100100000100000111010;
        end
        12101: begin
            cosine_reg0 <= 36'sb111101101101010000011010001101011010;
            sine_reg0   <= 36'sb100000000101010000111001011001010000;
        end
        12102: begin
            cosine_reg0 <= 36'sb111101101110000010100010111110011101;
            sine_reg0   <= 36'sb100000000101001101010011100000010111;
        end
        12103: begin
            cosine_reg0 <= 36'sb111101101110110100101011110101001000;
            sine_reg0   <= 36'sb100000000101001001101110110110001110;
        end
        12104: begin
            cosine_reg0 <= 36'sb111101101111100110110100110001011001;
            sine_reg0   <= 36'sb100000000101000110001011011010110101;
        end
        12105: begin
            cosine_reg0 <= 36'sb111101110000011000111101110011001110;
            sine_reg0   <= 36'sb100000000101000010101001001110001101;
        end
        12106: begin
            cosine_reg0 <= 36'sb111101110001001011000110111010100110;
            sine_reg0   <= 36'sb100000000100111111001000010000010110;
        end
        12107: begin
            cosine_reg0 <= 36'sb111101110001111101010000000111011110;
            sine_reg0   <= 36'sb100000000100111011101000100001010000;
        end
        12108: begin
            cosine_reg0 <= 36'sb111101110010101111011001011001110101;
            sine_reg0   <= 36'sb100000000100111000001010000000111011;
        end
        12109: begin
            cosine_reg0 <= 36'sb111101110011100001100010110001101000;
            sine_reg0   <= 36'sb100000000100110100101100101111010111;
        end
        12110: begin
            cosine_reg0 <= 36'sb111101110100010011101100001110110110;
            sine_reg0   <= 36'sb100000000100110001010000101100100100;
        end
        12111: begin
            cosine_reg0 <= 36'sb111101110101000101110101110001011100;
            sine_reg0   <= 36'sb100000000100101101110101111000100011;
        end
        12112: begin
            cosine_reg0 <= 36'sb111101110101110111111111011001011001;
            sine_reg0   <= 36'sb100000000100101010011100010011010011;
        end
        12113: begin
            cosine_reg0 <= 36'sb111101110110101010001001000110101011;
            sine_reg0   <= 36'sb100000000100100111000011111100110110;
        end
        12114: begin
            cosine_reg0 <= 36'sb111101110111011100010010111001010000;
            sine_reg0   <= 36'sb100000000100100011101100110101001010;
        end
        12115: begin
            cosine_reg0 <= 36'sb111101111000001110011100110001000110;
            sine_reg0   <= 36'sb100000000100100000010110111100010000;
        end
        12116: begin
            cosine_reg0 <= 36'sb111101111001000000100110101110001011;
            sine_reg0   <= 36'sb100000000100011101000010010010001000;
        end
        12117: begin
            cosine_reg0 <= 36'sb111101111001110010110000110000011101;
            sine_reg0   <= 36'sb100000000100011001101110110110110010;
        end
        12118: begin
            cosine_reg0 <= 36'sb111101111010100100111010110111111010;
            sine_reg0   <= 36'sb100000000100010110011100101010001111;
        end
        12119: begin
            cosine_reg0 <= 36'sb111101111011010111000101000100100000;
            sine_reg0   <= 36'sb100000000100010011001011101100011110;
        end
        12120: begin
            cosine_reg0 <= 36'sb111101111100001001001111010110001110;
            sine_reg0   <= 36'sb100000000100001111111011111101100000;
        end
        12121: begin
            cosine_reg0 <= 36'sb111101111100111011011001101101000001;
            sine_reg0   <= 36'sb100000000100001100101101011101010101;
        end
        12122: begin
            cosine_reg0 <= 36'sb111101111101101101100100001000110111;
            sine_reg0   <= 36'sb100000000100001001100000001011111101;
        end
        12123: begin
            cosine_reg0 <= 36'sb111101111110011111101110101001101111;
            sine_reg0   <= 36'sb100000000100000110010100001001010111;
        end
        12124: begin
            cosine_reg0 <= 36'sb111101111111010001111001001111100110;
            sine_reg0   <= 36'sb100000000100000011001001010101100101;
        end
        12125: begin
            cosine_reg0 <= 36'sb111110000000000100000011111010011011;
            sine_reg0   <= 36'sb100000000011111111111111110000100110;
        end
        12126: begin
            cosine_reg0 <= 36'sb111110000000110110001110101010001100;
            sine_reg0   <= 36'sb100000000011111100110111011010011010;
        end
        12127: begin
            cosine_reg0 <= 36'sb111110000001101000011001011110110110;
            sine_reg0   <= 36'sb100000000011111001110000010011000010;
        end
        12128: begin
            cosine_reg0 <= 36'sb111110000010011010100100011000011000;
            sine_reg0   <= 36'sb100000000011110110101010011010011101;
        end
        12129: begin
            cosine_reg0 <= 36'sb111110000011001100101111010110110000;
            sine_reg0   <= 36'sb100000000011110011100101110000101101;
        end
        12130: begin
            cosine_reg0 <= 36'sb111110000011111110111010011001111100;
            sine_reg0   <= 36'sb100000000011110000100010010101110000;
        end
        12131: begin
            cosine_reg0 <= 36'sb111110000100110001000101100001111010;
            sine_reg0   <= 36'sb100000000011101101100000001001100110;
        end
        12132: begin
            cosine_reg0 <= 36'sb111110000101100011010000101110101000;
            sine_reg0   <= 36'sb100000000011101010011111001100010001;
        end
        12133: begin
            cosine_reg0 <= 36'sb111110000110010101011100000000000100;
            sine_reg0   <= 36'sb100000000011100111011111011101110001;
        end
        12134: begin
            cosine_reg0 <= 36'sb111110000111000111100111010110001101;
            sine_reg0   <= 36'sb100000000011100100100000111110000100;
        end
        12135: begin
            cosine_reg0 <= 36'sb111110000111111001110010110000111111;
            sine_reg0   <= 36'sb100000000011100001100011101101001100;
        end
        12136: begin
            cosine_reg0 <= 36'sb111110001000101011111110010000011010;
            sine_reg0   <= 36'sb100000000011011110100111101011001001;
        end
        12137: begin
            cosine_reg0 <= 36'sb111110001001011110001001110100011011;
            sine_reg0   <= 36'sb100000000011011011101100110111111010;
        end
        12138: begin
            cosine_reg0 <= 36'sb111110001010010000010101011101000001;
            sine_reg0   <= 36'sb100000000011011000110011010011100000;
        end
        12139: begin
            cosine_reg0 <= 36'sb111110001011000010100001001010001001;
            sine_reg0   <= 36'sb100000000011010101111010111101111011;
        end
        12140: begin
            cosine_reg0 <= 36'sb111110001011110100101100111011110010;
            sine_reg0   <= 36'sb100000000011010011000011110111001010;
        end
        12141: begin
            cosine_reg0 <= 36'sb111110001100100110111000110001111010;
            sine_reg0   <= 36'sb100000000011010000001101111111001111;
        end
        12142: begin
            cosine_reg0 <= 36'sb111110001101011001000100101100011110;
            sine_reg0   <= 36'sb100000000011001101011001010110001001;
        end
        12143: begin
            cosine_reg0 <= 36'sb111110001110001011010000101011011101;
            sine_reg0   <= 36'sb100000000011001010100101111011111001;
        end
        12144: begin
            cosine_reg0 <= 36'sb111110001110111101011100101110110101;
            sine_reg0   <= 36'sb100000000011000111110011110000011110;
        end
        12145: begin
            cosine_reg0 <= 36'sb111110001111101111101000110110100100;
            sine_reg0   <= 36'sb100000000011000101000010110011111000;
        end
        12146: begin
            cosine_reg0 <= 36'sb111110010000100001110101000010101000;
            sine_reg0   <= 36'sb100000000011000010010011000110001000;
        end
        12147: begin
            cosine_reg0 <= 36'sb111110010001010100000001010010111110;
            sine_reg0   <= 36'sb100000000010111111100100100111001110;
        end
        12148: begin
            cosine_reg0 <= 36'sb111110010010000110001101100111100110;
            sine_reg0   <= 36'sb100000000010111100110111010111001001;
        end
        12149: begin
            cosine_reg0 <= 36'sb111110010010111000011010000000011110;
            sine_reg0   <= 36'sb100000000010111010001011010101111011;
        end
        12150: begin
            cosine_reg0 <= 36'sb111110010011101010100110011101100010;
            sine_reg0   <= 36'sb100000000010110111100000100011100011;
        end
        12151: begin
            cosine_reg0 <= 36'sb111110010100011100110010111110110010;
            sine_reg0   <= 36'sb100000000010110100110111000000000000;
        end
        12152: begin
            cosine_reg0 <= 36'sb111110010101001110111111100100001011;
            sine_reg0   <= 36'sb100000000010110010001110101011010101;
        end
        12153: begin
            cosine_reg0 <= 36'sb111110010110000001001100001101101011;
            sine_reg0   <= 36'sb100000000010101111100111100101011111;
        end
        12154: begin
            cosine_reg0 <= 36'sb111110010110110011011000111011010001;
            sine_reg0   <= 36'sb100000000010101101000001101110100000;
        end
        12155: begin
            cosine_reg0 <= 36'sb111110010111100101100101101100111011;
            sine_reg0   <= 36'sb100000000010101010011101000110010111;
        end
        12156: begin
            cosine_reg0 <= 36'sb111110011000010111110010100010100110;
            sine_reg0   <= 36'sb100000000010100111111001101101000101;
        end
        12157: begin
            cosine_reg0 <= 36'sb111110011001001001111111011100010001;
            sine_reg0   <= 36'sb100000000010100101010111100010101010;
        end
        12158: begin
            cosine_reg0 <= 36'sb111110011001111100001100011001111001;
            sine_reg0   <= 36'sb100000000010100010110110100111000110;
        end
        12159: begin
            cosine_reg0 <= 36'sb111110011010101110011001011011011110;
            sine_reg0   <= 36'sb100000000010100000010110111010011001;
        end
        12160: begin
            cosine_reg0 <= 36'sb111110011011100000100110100000111100;
            sine_reg0   <= 36'sb100000000010011101111000011100100011;
        end
        12161: begin
            cosine_reg0 <= 36'sb111110011100010010110011101010010010;
            sine_reg0   <= 36'sb100000000010011011011011001101100100;
        end
        12162: begin
            cosine_reg0 <= 36'sb111110011101000101000000110111011110;
            sine_reg0   <= 36'sb100000000010011000111111001101011100;
        end
        12163: begin
            cosine_reg0 <= 36'sb111110011101110111001110001000011111;
            sine_reg0   <= 36'sb100000000010010110100100011100001011;
        end
        12164: begin
            cosine_reg0 <= 36'sb111110011110101001011011011101010001;
            sine_reg0   <= 36'sb100000000010010100001010111001110010;
        end
        12165: begin
            cosine_reg0 <= 36'sb111110011111011011101000110101110100;
            sine_reg0   <= 36'sb100000000010010001110010100110010001;
        end
        12166: begin
            cosine_reg0 <= 36'sb111110100000001101110110010010000101;
            sine_reg0   <= 36'sb100000000010001111011011100001100111;
        end
        12167: begin
            cosine_reg0 <= 36'sb111110100001000000000011110010000010;
            sine_reg0   <= 36'sb100000000010001101000101101011110101;
        end
        12168: begin
            cosine_reg0 <= 36'sb111110100001110010010001010101101010;
            sine_reg0   <= 36'sb100000000010001010110001000100111010;
        end
        12169: begin
            cosine_reg0 <= 36'sb111110100010100100011110111100111010;
            sine_reg0   <= 36'sb100000000010001000011101101100111000;
        end
        12170: begin
            cosine_reg0 <= 36'sb111110100011010110101100100111110001;
            sine_reg0   <= 36'sb100000000010000110001011100011101101;
        end
        12171: begin
            cosine_reg0 <= 36'sb111110100100001000111010010110001100;
            sine_reg0   <= 36'sb100000000010000011111010101001011011;
        end
        12172: begin
            cosine_reg0 <= 36'sb111110100100111011001000001000001010;
            sine_reg0   <= 36'sb100000000010000001101010111110000000;
        end
        12173: begin
            cosine_reg0 <= 36'sb111110100101101101010101111101101001;
            sine_reg0   <= 36'sb100000000001111111011100100001011110;
        end
        12174: begin
            cosine_reg0 <= 36'sb111110100110011111100011110110100110;
            sine_reg0   <= 36'sb100000000001111101001111010011110100;
        end
        12175: begin
            cosine_reg0 <= 36'sb111110100111010001110001110011000001;
            sine_reg0   <= 36'sb100000000001111011000011010101000011;
        end
        12176: begin
            cosine_reg0 <= 36'sb111110101000000011111111110010110110;
            sine_reg0   <= 36'sb100000000001111000111000100101001010;
        end
        12177: begin
            cosine_reg0 <= 36'sb111110101000110110001101110110000100;
            sine_reg0   <= 36'sb100000000001110110101111000100001010;
        end
        12178: begin
            cosine_reg0 <= 36'sb111110101001101000011011111100101001;
            sine_reg0   <= 36'sb100000000001110100100110110010000010;
        end
        12179: begin
            cosine_reg0 <= 36'sb111110101010011010101010000110100100;
            sine_reg0   <= 36'sb100000000001110010011111101110110011;
        end
        12180: begin
            cosine_reg0 <= 36'sb111110101011001100111000010011110001;
            sine_reg0   <= 36'sb100000000001110000011001111010011101;
        end
        12181: begin
            cosine_reg0 <= 36'sb111110101011111111000110100100010000;
            sine_reg0   <= 36'sb100000000001101110010101010101000000;
        end
        12182: begin
            cosine_reg0 <= 36'sb111110101100110001010100110111111110;
            sine_reg0   <= 36'sb100000000001101100010001111110011100;
        end
        12183: begin
            cosine_reg0 <= 36'sb111110101101100011100011001110111001;
            sine_reg0   <= 36'sb100000000001101010001111110110110001;
        end
        12184: begin
            cosine_reg0 <= 36'sb111110101110010101110001101001000000;
            sine_reg0   <= 36'sb100000000001101000001110111101111111;
        end
        12185: begin
            cosine_reg0 <= 36'sb111110101111001000000000000110010000;
            sine_reg0   <= 36'sb100000000001100110001111010100000110;
        end
        12186: begin
            cosine_reg0 <= 36'sb111110101111111010001110100110101000;
            sine_reg0   <= 36'sb100000000001100100010000111001000111;
        end
        12187: begin
            cosine_reg0 <= 36'sb111110110000101100011101001010000110;
            sine_reg0   <= 36'sb100000000001100010010011101101000001;
        end
        12188: begin
            cosine_reg0 <= 36'sb111110110001011110101011110000100111;
            sine_reg0   <= 36'sb100000000001100000010111101111110100;
        end
        12189: begin
            cosine_reg0 <= 36'sb111110110010010000111010011010001010;
            sine_reg0   <= 36'sb100000000001011110011101000001100001;
        end
        12190: begin
            cosine_reg0 <= 36'sb111110110011000011001001000110101101;
            sine_reg0   <= 36'sb100000000001011100100011100010000111;
        end
        12191: begin
            cosine_reg0 <= 36'sb111110110011110101010111110110001101;
            sine_reg0   <= 36'sb100000000001011010101011010001100111;
        end
        12192: begin
            cosine_reg0 <= 36'sb111110110100100111100110101000101010;
            sine_reg0   <= 36'sb100000000001011000110100010000000001;
        end
        12193: begin
            cosine_reg0 <= 36'sb111110110101011001110101011110000000;
            sine_reg0   <= 36'sb100000000001010110111110011101010101;
        end
        12194: begin
            cosine_reg0 <= 36'sb111110110110001100000100010110001111;
            sine_reg0   <= 36'sb100000000001010101001001111001100011;
        end
        12195: begin
            cosine_reg0 <= 36'sb111110110110111110010011010001010011;
            sine_reg0   <= 36'sb100000000001010011010110100100101010;
        end
        12196: begin
            cosine_reg0 <= 36'sb111110110111110000100010001111001100;
            sine_reg0   <= 36'sb100000000001010001100100011110101100;
        end
        12197: begin
            cosine_reg0 <= 36'sb111110111000100010110001001111110111;
            sine_reg0   <= 36'sb100000000001001111110011100111100111;
        end
        12198: begin
            cosine_reg0 <= 36'sb111110111001010101000000010011010011;
            sine_reg0   <= 36'sb100000000001001110000011111111011101;
        end
        12199: begin
            cosine_reg0 <= 36'sb111110111010000111001111011001011101;
            sine_reg0   <= 36'sb100000000001001100010101100110001101;
        end
        12200: begin
            cosine_reg0 <= 36'sb111110111010111001011110100010010011;
            sine_reg0   <= 36'sb100000000001001010101000011011111000;
        end
        12201: begin
            cosine_reg0 <= 36'sb111110111011101011101101101101110100;
            sine_reg0   <= 36'sb100000000001001000111100100000011100;
        end
        12202: begin
            cosine_reg0 <= 36'sb111110111100011101111100111011111101;
            sine_reg0   <= 36'sb100000000001000111010001110011111011;
        end
        12203: begin
            cosine_reg0 <= 36'sb111110111101010000001100001100101101;
            sine_reg0   <= 36'sb100000000001000101101000010110010101;
        end
        12204: begin
            cosine_reg0 <= 36'sb111110111110000010011011100000000010;
            sine_reg0   <= 36'sb100000000001000100000000000111101001;
        end
        12205: begin
            cosine_reg0 <= 36'sb111110111110110100101010110101111001;
            sine_reg0   <= 36'sb100000000001000010011001000111111000;
        end
        12206: begin
            cosine_reg0 <= 36'sb111110111111100110111010001110010001;
            sine_reg0   <= 36'sb100000000001000000110011010111000001;
        end
        12207: begin
            cosine_reg0 <= 36'sb111111000000011001001001101001001000;
            sine_reg0   <= 36'sb100000000000111111001110110101000110;
        end
        12208: begin
            cosine_reg0 <= 36'sb111111000001001011011001000110011100;
            sine_reg0   <= 36'sb100000000000111101101011100010000101;
        end
        12209: begin
            cosine_reg0 <= 36'sb111111000001111101101000100110001011;
            sine_reg0   <= 36'sb100000000000111100001001011101111110;
        end
        12210: begin
            cosine_reg0 <= 36'sb111111000010101111111000001000010100;
            sine_reg0   <= 36'sb100000000000111010101000101000110011;
        end
        12211: begin
            cosine_reg0 <= 36'sb111111000011100010000111101100110011;
            sine_reg0   <= 36'sb100000000000111001001001000010100011;
        end
        12212: begin
            cosine_reg0 <= 36'sb111111000100010100010111010011100111;
            sine_reg0   <= 36'sb100000000000110111101010101011001110;
        end
        12213: begin
            cosine_reg0 <= 36'sb111111000101000110100110111100101111;
            sine_reg0   <= 36'sb100000000000110110001101100010110100;
        end
        12214: begin
            cosine_reg0 <= 36'sb111111000101111000110110101000001000;
            sine_reg0   <= 36'sb100000000000110100110001101001010101;
        end
        12215: begin
            cosine_reg0 <= 36'sb111111000110101011000110010101110000;
            sine_reg0   <= 36'sb100000000000110011010110111110110001;
        end
        12216: begin
            cosine_reg0 <= 36'sb111111000111011101010110000101100110;
            sine_reg0   <= 36'sb100000000000110001111101100011001000;
        end
        12217: begin
            cosine_reg0 <= 36'sb111111001000001111100101110111101000;
            sine_reg0   <= 36'sb100000000000110000100101010110011011;
        end
        12218: begin
            cosine_reg0 <= 36'sb111111001001000001110101101011110011;
            sine_reg0   <= 36'sb100000000000101111001110011000101001;
        end
        12219: begin
            cosine_reg0 <= 36'sb111111001001110100000101100010000101;
            sine_reg0   <= 36'sb100000000000101101111000101001110011;
        end
        12220: begin
            cosine_reg0 <= 36'sb111111001010100110010101011010011101;
            sine_reg0   <= 36'sb100000000000101100100100001001111000;
        end
        12221: begin
            cosine_reg0 <= 36'sb111111001011011000100101010100111001;
            sine_reg0   <= 36'sb100000000000101011010000111000111000;
        end
        12222: begin
            cosine_reg0 <= 36'sb111111001100001010110101010001010111;
            sine_reg0   <= 36'sb100000000000101001111110110110110101;
        end
        12223: begin
            cosine_reg0 <= 36'sb111111001100111101000101001111110101;
            sine_reg0   <= 36'sb100000000000101000101110000011101100;
        end
        12224: begin
            cosine_reg0 <= 36'sb111111001101101111010101010000010001;
            sine_reg0   <= 36'sb100000000000100111011110011111100000;
        end
        12225: begin
            cosine_reg0 <= 36'sb111111001110100001100101010010101000;
            sine_reg0   <= 36'sb100000000000100110010000001010001111;
        end
        12226: begin
            cosine_reg0 <= 36'sb111111001111010011110101010110111010;
            sine_reg0   <= 36'sb100000000000100101000011000011111010;
        end
        12227: begin
            cosine_reg0 <= 36'sb111111010000000110000101011101000100;
            sine_reg0   <= 36'sb100000000000100011110111001100100001;
        end
        12228: begin
            cosine_reg0 <= 36'sb111111010000111000010101100101000100;
            sine_reg0   <= 36'sb100000000000100010101100100100000011;
        end
        12229: begin
            cosine_reg0 <= 36'sb111111010001101010100101101110111001;
            sine_reg0   <= 36'sb100000000000100001100011001010100010;
        end
        12230: begin
            cosine_reg0 <= 36'sb111111010010011100110101111010011111;
            sine_reg0   <= 36'sb100000000000100000011010111111111100;
        end
        12231: begin
            cosine_reg0 <= 36'sb111111010011001111000110000111110111;
            sine_reg0   <= 36'sb100000000000011111010100000100010010;
        end
        12232: begin
            cosine_reg0 <= 36'sb111111010100000001010110010110111100;
            sine_reg0   <= 36'sb100000000000011110001110010111100101;
        end
        12233: begin
            cosine_reg0 <= 36'sb111111010100110011100110100111101110;
            sine_reg0   <= 36'sb100000000000011101001001111001110011;
        end
        12234: begin
            cosine_reg0 <= 36'sb111111010101100101110110111010001011;
            sine_reg0   <= 36'sb100000000000011100000110101010111110;
        end
        12235: begin
            cosine_reg0 <= 36'sb111111010110011000000111001110010000;
            sine_reg0   <= 36'sb100000000000011011000100101011000101;
        end
        12236: begin
            cosine_reg0 <= 36'sb111111010111001010010111100011111100;
            sine_reg0   <= 36'sb100000000000011010000011111010001000;
        end
        12237: begin
            cosine_reg0 <= 36'sb111111010111111100100111111011001101;
            sine_reg0   <= 36'sb100000000000011001000100011000000111;
        end
        12238: begin
            cosine_reg0 <= 36'sb111111011000101110111000010100000000;
            sine_reg0   <= 36'sb100000000000011000000110000101000010;
        end
        12239: begin
            cosine_reg0 <= 36'sb111111011001100001001000101110010101;
            sine_reg0   <= 36'sb100000000000010111001001000000111010;
        end
        12240: begin
            cosine_reg0 <= 36'sb111111011010010011011001001010001000;
            sine_reg0   <= 36'sb100000000000010110001101001011101110;
        end
        12241: begin
            cosine_reg0 <= 36'sb111111011011000101101001100111011001;
            sine_reg0   <= 36'sb100000000000010101010010100101011111;
        end
        12242: begin
            cosine_reg0 <= 36'sb111111011011110111111010000110000100;
            sine_reg0   <= 36'sb100000000000010100011001001110001100;
        end
        12243: begin
            cosine_reg0 <= 36'sb111111011100101010001010100110001001;
            sine_reg0   <= 36'sb100000000000010011100001000101110101;
        end
        12244: begin
            cosine_reg0 <= 36'sb111111011101011100011011000111100101;
            sine_reg0   <= 36'sb100000000000010010101010001100011011;
        end
        12245: begin
            cosine_reg0 <= 36'sb111111011110001110101011101010010110;
            sine_reg0   <= 36'sb100000000000010001110100100001111101;
        end
        12246: begin
            cosine_reg0 <= 36'sb111111011111000000111100001110011010;
            sine_reg0   <= 36'sb100000000000010001000000000110011100;
        end
        12247: begin
            cosine_reg0 <= 36'sb111111011111110011001100110011110000;
            sine_reg0   <= 36'sb100000000000010000001100111001111000;
        end
        12248: begin
            cosine_reg0 <= 36'sb111111100000100101011101011010010101;
            sine_reg0   <= 36'sb100000000000001111011010111100010000;
        end
        12249: begin
            cosine_reg0 <= 36'sb111111100001010111101110000010001000;
            sine_reg0   <= 36'sb100000000000001110101010001101100100;
        end
        12250: begin
            cosine_reg0 <= 36'sb111111100010001001111110101011000110;
            sine_reg0   <= 36'sb100000000000001101111010101101110110;
        end
        12251: begin
            cosine_reg0 <= 36'sb111111100010111100001111010101001110;
            sine_reg0   <= 36'sb100000000000001101001100011101000100;
        end
        12252: begin
            cosine_reg0 <= 36'sb111111100011101110100000000000011110;
            sine_reg0   <= 36'sb100000000000001100011111011011001111;
        end
        12253: begin
            cosine_reg0 <= 36'sb111111100100100000110000101100110100;
            sine_reg0   <= 36'sb100000000000001011110011101000010110;
        end
        12254: begin
            cosine_reg0 <= 36'sb111111100101010011000001011010001101;
            sine_reg0   <= 36'sb100000000000001011001001000100011011;
        end
        12255: begin
            cosine_reg0 <= 36'sb111111100110000101010010001000101000;
            sine_reg0   <= 36'sb100000000000001010011111101111011100;
        end
        12256: begin
            cosine_reg0 <= 36'sb111111100110110111100010111000000011;
            sine_reg0   <= 36'sb100000000000001001110111101001011010;
        end
        12257: begin
            cosine_reg0 <= 36'sb111111100111101001110011101000011100;
            sine_reg0   <= 36'sb100000000000001001010000110010010101;
        end
        12258: begin
            cosine_reg0 <= 36'sb111111101000011100000100011001110001;
            sine_reg0   <= 36'sb100000000000001000101011001010001101;
        end
        12259: begin
            cosine_reg0 <= 36'sb111111101001001110010101001100000001;
            sine_reg0   <= 36'sb100000000000001000000110110001000001;
        end
        12260: begin
            cosine_reg0 <= 36'sb111111101010000000100101111111001000;
            sine_reg0   <= 36'sb100000000000000111100011100110110011;
        end
        12261: begin
            cosine_reg0 <= 36'sb111111101010110010110110110011000110;
            sine_reg0   <= 36'sb100000000000000111000001101011100010;
        end
        12262: begin
            cosine_reg0 <= 36'sb111111101011100101000111100111111000;
            sine_reg0   <= 36'sb100000000000000110100000111111001101;
        end
        12263: begin
            cosine_reg0 <= 36'sb111111101100010111011000011101011101;
            sine_reg0   <= 36'sb100000000000000110000001100001110110;
        end
        12264: begin
            cosine_reg0 <= 36'sb111111101101001001101001010011110010;
            sine_reg0   <= 36'sb100000000000000101100011010011011011;
        end
        12265: begin
            cosine_reg0 <= 36'sb111111101101111011111010001010110101;
            sine_reg0   <= 36'sb100000000000000101000110010011111110;
        end
        12266: begin
            cosine_reg0 <= 36'sb111111101110101110001011000010100101;
            sine_reg0   <= 36'sb100000000000000100101010100011011101;
        end
        12267: begin
            cosine_reg0 <= 36'sb111111101111100000011011111011000000;
            sine_reg0   <= 36'sb100000000000000100010000000001111010;
        end
        12268: begin
            cosine_reg0 <= 36'sb111111110000010010101100110100000011;
            sine_reg0   <= 36'sb100000000000000011110110101111010100;
        end
        12269: begin
            cosine_reg0 <= 36'sb111111110001000100111101101101101101;
            sine_reg0   <= 36'sb100000000000000011011110101011101010;
        end
        12270: begin
            cosine_reg0 <= 36'sb111111110001110111001110100111111100;
            sine_reg0   <= 36'sb100000000000000011000111110110111110;
        end
        12271: begin
            cosine_reg0 <= 36'sb111111110010101001011111100010101110;
            sine_reg0   <= 36'sb100000000000000010110010010001001111;
        end
        12272: begin
            cosine_reg0 <= 36'sb111111110011011011110000011110000001;
            sine_reg0   <= 36'sb100000000000000010011101111010011101;
        end
        12273: begin
            cosine_reg0 <= 36'sb111111110100001110000001011001110011;
            sine_reg0   <= 36'sb100000000000000010001010110010101001;
        end
        12274: begin
            cosine_reg0 <= 36'sb111111110101000000010010010110000001;
            sine_reg0   <= 36'sb100000000000000001111000111001110001;
        end
        12275: begin
            cosine_reg0 <= 36'sb111111110101110010100011010010101011;
            sine_reg0   <= 36'sb100000000000000001101000001111110111;
        end
        12276: begin
            cosine_reg0 <= 36'sb111111110110100100110100001111101111;
            sine_reg0   <= 36'sb100000000000000001011000110100111001;
        end
        12277: begin
            cosine_reg0 <= 36'sb111111110111010111000101001101001001;
            sine_reg0   <= 36'sb100000000000000001001010101000111001;
        end
        12278: begin
            cosine_reg0 <= 36'sb111111111000001001010110001010111001;
            sine_reg0   <= 36'sb100000000000000000111101101011110111;
        end
        12279: begin
            cosine_reg0 <= 36'sb111111111000111011100111001000111100;
            sine_reg0   <= 36'sb100000000000000000110001111101110001;
        end
        12280: begin
            cosine_reg0 <= 36'sb111111111001101101111000000111010000;
            sine_reg0   <= 36'sb100000000000000000100111011110101000;
        end
        12281: begin
            cosine_reg0 <= 36'sb111111111010100000001001000101110100;
            sine_reg0   <= 36'sb100000000000000000011110001110011101;
        end
        12282: begin
            cosine_reg0 <= 36'sb111111111011010010011010000100100110;
            sine_reg0   <= 36'sb100000000000000000010110001101001111;
        end
        12283: begin
            cosine_reg0 <= 36'sb111111111100000100101011000011100011;
            sine_reg0   <= 36'sb100000000000000000001111011010111110;
        end
        12284: begin
            cosine_reg0 <= 36'sb111111111100110110111100000010101010;
            sine_reg0   <= 36'sb100000000000000000001001110111101011;
        end
        12285: begin
            cosine_reg0 <= 36'sb111111111101101001001101000001111001;
            sine_reg0   <= 36'sb100000000000000000000101100011010101;
        end
        12286: begin
            cosine_reg0 <= 36'sb111111111110011011011110000001001101;
            sine_reg0   <= 36'sb100000000000000000000010011101111011;
        end
        12287: begin
            cosine_reg0 <= 36'sb111111111111001101101111000000100110;
            sine_reg0   <= 36'sb100000000000000000000000100111100000;
        end
        12288: begin
            cosine_reg0 <= 36'sb0;
            sine_reg0   <= 36'sb100000000000000000000000000000000001;
        end
        12289: begin
            cosine_reg0 <= 36'sb110010010000111111011010;
            sine_reg0   <= 36'sb100000000000000000000000100111100000;
        end
        12290: begin
            cosine_reg0 <= 36'sb1100100100001111110110011;
            sine_reg0   <= 36'sb100000000000000000000010011101111011;
        end
        12291: begin
            cosine_reg0 <= 36'sb10010110110010111110000111;
            sine_reg0   <= 36'sb100000000000000000000101100011010101;
        end
        12292: begin
            cosine_reg0 <= 36'sb11001001000011111101010110;
            sine_reg0   <= 36'sb100000000000000000001001110111101011;
        end
        12293: begin
            cosine_reg0 <= 36'sb11111011010100111100011101;
            sine_reg0   <= 36'sb100000000000000000001111011010111110;
        end
        12294: begin
            cosine_reg0 <= 36'sb100101101100101111011011010;
            sine_reg0   <= 36'sb100000000000000000010110001101001111;
        end
        12295: begin
            cosine_reg0 <= 36'sb101011111110110111010001100;
            sine_reg0   <= 36'sb100000000000000000011110001110011101;
        end
        12296: begin
            cosine_reg0 <= 36'sb110010010000111111000110000;
            sine_reg0   <= 36'sb100000000000000000100111011110101000;
        end
        12297: begin
            cosine_reg0 <= 36'sb111000100011000110111000100;
            sine_reg0   <= 36'sb100000000000000000110001111101110001;
        end
        12298: begin
            cosine_reg0 <= 36'sb111110110101001110101000111;
            sine_reg0   <= 36'sb100000000000000000111101101011110111;
        end
        12299: begin
            cosine_reg0 <= 36'sb1000101000111010110010110111;
            sine_reg0   <= 36'sb100000000000000001001010101000111001;
        end
        12300: begin
            cosine_reg0 <= 36'sb1001011011001011110000010001;
            sine_reg0   <= 36'sb100000000000000001011000110100111001;
        end
        12301: begin
            cosine_reg0 <= 36'sb1010001101011100101101010101;
            sine_reg0   <= 36'sb100000000000000001101000001111110111;
        end
        12302: begin
            cosine_reg0 <= 36'sb1010111111101101101001111111;
            sine_reg0   <= 36'sb100000000000000001111000111001110001;
        end
        12303: begin
            cosine_reg0 <= 36'sb1011110001111110100110001101;
            sine_reg0   <= 36'sb100000000000000010001010110010101001;
        end
        12304: begin
            cosine_reg0 <= 36'sb1100100100001111100001111111;
            sine_reg0   <= 36'sb100000000000000010011101111010011101;
        end
        12305: begin
            cosine_reg0 <= 36'sb1101010110100000011101010010;
            sine_reg0   <= 36'sb100000000000000010110010010001001111;
        end
        12306: begin
            cosine_reg0 <= 36'sb1110001000110001011000000100;
            sine_reg0   <= 36'sb100000000000000011000111110110111110;
        end
        12307: begin
            cosine_reg0 <= 36'sb1110111011000010010010010011;
            sine_reg0   <= 36'sb100000000000000011011110101011101010;
        end
        12308: begin
            cosine_reg0 <= 36'sb1111101101010011001011111101;
            sine_reg0   <= 36'sb100000000000000011110110101111010100;
        end
        12309: begin
            cosine_reg0 <= 36'sb10000011111100100000101000000;
            sine_reg0   <= 36'sb100000000000000100010000000001111010;
        end
        12310: begin
            cosine_reg0 <= 36'sb10001010001110100111101011011;
            sine_reg0   <= 36'sb100000000000000100101010100011011101;
        end
        12311: begin
            cosine_reg0 <= 36'sb10010000100000101110101001011;
            sine_reg0   <= 36'sb100000000000000101000110010011111110;
        end
        12312: begin
            cosine_reg0 <= 36'sb10010110110010110101100001110;
            sine_reg0   <= 36'sb100000000000000101100011010011011011;
        end
        12313: begin
            cosine_reg0 <= 36'sb10011101000100111100010100011;
            sine_reg0   <= 36'sb100000000000000110000001100001110110;
        end
        12314: begin
            cosine_reg0 <= 36'sb10100011010111000011000001000;
            sine_reg0   <= 36'sb100000000000000110100000111111001101;
        end
        12315: begin
            cosine_reg0 <= 36'sb10101001101001001001100111010;
            sine_reg0   <= 36'sb100000000000000111000001101011100010;
        end
        12316: begin
            cosine_reg0 <= 36'sb10101111111011010000000111000;
            sine_reg0   <= 36'sb100000000000000111100011100110110011;
        end
        12317: begin
            cosine_reg0 <= 36'sb10110110001101010110011111111;
            sine_reg0   <= 36'sb100000000000001000000110110001000001;
        end
        12318: begin
            cosine_reg0 <= 36'sb10111100011111011100110001111;
            sine_reg0   <= 36'sb100000000000001000101011001010001101;
        end
        12319: begin
            cosine_reg0 <= 36'sb11000010110001100010111100100;
            sine_reg0   <= 36'sb100000000000001001010000110010010101;
        end
        12320: begin
            cosine_reg0 <= 36'sb11001001000011101000111111101;
            sine_reg0   <= 36'sb100000000000001001110111101001011010;
        end
        12321: begin
            cosine_reg0 <= 36'sb11001111010101101110111011000;
            sine_reg0   <= 36'sb100000000000001010011111101111011100;
        end
        12322: begin
            cosine_reg0 <= 36'sb11010101100111110100101110011;
            sine_reg0   <= 36'sb100000000000001011001001000100011011;
        end
        12323: begin
            cosine_reg0 <= 36'sb11011011111001111010011001100;
            sine_reg0   <= 36'sb100000000000001011110011101000010110;
        end
        12324: begin
            cosine_reg0 <= 36'sb11100010001011111111111100010;
            sine_reg0   <= 36'sb100000000000001100011111011011001111;
        end
        12325: begin
            cosine_reg0 <= 36'sb11101000011110000101010110010;
            sine_reg0   <= 36'sb100000000000001101001100011101000100;
        end
        12326: begin
            cosine_reg0 <= 36'sb11101110110000001010100111010;
            sine_reg0   <= 36'sb100000000000001101111010101101110110;
        end
        12327: begin
            cosine_reg0 <= 36'sb11110101000010001111101111000;
            sine_reg0   <= 36'sb100000000000001110101010001101100100;
        end
        12328: begin
            cosine_reg0 <= 36'sb11111011010100010100101101011;
            sine_reg0   <= 36'sb100000000000001111011010111100010000;
        end
        12329: begin
            cosine_reg0 <= 36'sb100000001100110011001100010000;
            sine_reg0   <= 36'sb100000000000010000001100111001111000;
        end
        12330: begin
            cosine_reg0 <= 36'sb100000111111000011110001100110;
            sine_reg0   <= 36'sb100000000000010001000000000110011100;
        end
        12331: begin
            cosine_reg0 <= 36'sb100001110001010100010101101010;
            sine_reg0   <= 36'sb100000000000010001110100100001111101;
        end
        12332: begin
            cosine_reg0 <= 36'sb100010100011100100111000011011;
            sine_reg0   <= 36'sb100000000000010010101010001100011011;
        end
        12333: begin
            cosine_reg0 <= 36'sb100011010101110101011001110111;
            sine_reg0   <= 36'sb100000000000010011100001000101110101;
        end
        12334: begin
            cosine_reg0 <= 36'sb100100001000000101111001111100;
            sine_reg0   <= 36'sb100000000000010100011001001110001100;
        end
        12335: begin
            cosine_reg0 <= 36'sb100100111010010110011000100111;
            sine_reg0   <= 36'sb100000000000010101010010100101011111;
        end
        12336: begin
            cosine_reg0 <= 36'sb100101101100100110110101111000;
            sine_reg0   <= 36'sb100000000000010110001101001011101110;
        end
        12337: begin
            cosine_reg0 <= 36'sb100110011110110111010001101011;
            sine_reg0   <= 36'sb100000000000010111001001000000111010;
        end
        12338: begin
            cosine_reg0 <= 36'sb100111010001000111101100000000;
            sine_reg0   <= 36'sb100000000000011000000110000101000010;
        end
        12339: begin
            cosine_reg0 <= 36'sb101000000011011000000100110011;
            sine_reg0   <= 36'sb100000000000011001000100011000000111;
        end
        12340: begin
            cosine_reg0 <= 36'sb101000110101101000011100000100;
            sine_reg0   <= 36'sb100000000000011010000011111010001000;
        end
        12341: begin
            cosine_reg0 <= 36'sb101001100111111000110001110000;
            sine_reg0   <= 36'sb100000000000011011000100101011000101;
        end
        12342: begin
            cosine_reg0 <= 36'sb101010011010001001000101110101;
            sine_reg0   <= 36'sb100000000000011100000110101010111110;
        end
        12343: begin
            cosine_reg0 <= 36'sb101011001100011001011000010010;
            sine_reg0   <= 36'sb100000000000011101001001111001110011;
        end
        12344: begin
            cosine_reg0 <= 36'sb101011111110101001101001000100;
            sine_reg0   <= 36'sb100000000000011110001110010111100101;
        end
        12345: begin
            cosine_reg0 <= 36'sb101100110000111001111000001001;
            sine_reg0   <= 36'sb100000000000011111010100000100010010;
        end
        12346: begin
            cosine_reg0 <= 36'sb101101100011001010000101100001;
            sine_reg0   <= 36'sb100000000000100000011010111111111100;
        end
        12347: begin
            cosine_reg0 <= 36'sb101110010101011010010001000111;
            sine_reg0   <= 36'sb100000000000100001100011001010100010;
        end
        12348: begin
            cosine_reg0 <= 36'sb101111000111101010011010111100;
            sine_reg0   <= 36'sb100000000000100010101100100100000011;
        end
        12349: begin
            cosine_reg0 <= 36'sb101111111001111010100010111100;
            sine_reg0   <= 36'sb100000000000100011110111001100100001;
        end
        12350: begin
            cosine_reg0 <= 36'sb110000101100001010101001000110;
            sine_reg0   <= 36'sb100000000000100101000011000011111010;
        end
        12351: begin
            cosine_reg0 <= 36'sb110001011110011010101101011000;
            sine_reg0   <= 36'sb100000000000100110010000001010001111;
        end
        12352: begin
            cosine_reg0 <= 36'sb110010010000101010101111101111;
            sine_reg0   <= 36'sb100000000000100111011110011111100000;
        end
        12353: begin
            cosine_reg0 <= 36'sb110011000010111010110000001011;
            sine_reg0   <= 36'sb100000000000101000101110000011101100;
        end
        12354: begin
            cosine_reg0 <= 36'sb110011110101001010101110101001;
            sine_reg0   <= 36'sb100000000000101001111110110110110101;
        end
        12355: begin
            cosine_reg0 <= 36'sb110100100111011010101011000111;
            sine_reg0   <= 36'sb100000000000101011010000111000111000;
        end
        12356: begin
            cosine_reg0 <= 36'sb110101011001101010100101100011;
            sine_reg0   <= 36'sb100000000000101100100100001001111000;
        end
        12357: begin
            cosine_reg0 <= 36'sb110110001011111010011101111011;
            sine_reg0   <= 36'sb100000000000101101111000101001110011;
        end
        12358: begin
            cosine_reg0 <= 36'sb110110111110001010010100001101;
            sine_reg0   <= 36'sb100000000000101111001110011000101001;
        end
        12359: begin
            cosine_reg0 <= 36'sb110111110000011010001000011000;
            sine_reg0   <= 36'sb100000000000110000100101010110011011;
        end
        12360: begin
            cosine_reg0 <= 36'sb111000100010101001111010011010;
            sine_reg0   <= 36'sb100000000000110001111101100011001000;
        end
        12361: begin
            cosine_reg0 <= 36'sb111001010100111001101010010000;
            sine_reg0   <= 36'sb100000000000110011010110111110110001;
        end
        12362: begin
            cosine_reg0 <= 36'sb111010000111001001010111111000;
            sine_reg0   <= 36'sb100000000000110100110001101001010101;
        end
        12363: begin
            cosine_reg0 <= 36'sb111010111001011001000011010001;
            sine_reg0   <= 36'sb100000000000110110001101100010110100;
        end
        12364: begin
            cosine_reg0 <= 36'sb111011101011101000101100011001;
            sine_reg0   <= 36'sb100000000000110111101010101011001110;
        end
        12365: begin
            cosine_reg0 <= 36'sb111100011101111000010011001101;
            sine_reg0   <= 36'sb100000000000111001001001000010100011;
        end
        12366: begin
            cosine_reg0 <= 36'sb111101010000000111110111101100;
            sine_reg0   <= 36'sb100000000000111010101000101000110011;
        end
        12367: begin
            cosine_reg0 <= 36'sb111110000010010111011001110101;
            sine_reg0   <= 36'sb100000000000111100001001011101111110;
        end
        12368: begin
            cosine_reg0 <= 36'sb111110110100100110111001100100;
            sine_reg0   <= 36'sb100000000000111101101011100010000101;
        end
        12369: begin
            cosine_reg0 <= 36'sb111111100110110110010110111000;
            sine_reg0   <= 36'sb100000000000111111001110110101000110;
        end
        12370: begin
            cosine_reg0 <= 36'sb1000000011001000101110001101111;
            sine_reg0   <= 36'sb100000000001000000110011010111000001;
        end
        12371: begin
            cosine_reg0 <= 36'sb1000001001011010101001010000111;
            sine_reg0   <= 36'sb100000000001000010011001000111111000;
        end
        12372: begin
            cosine_reg0 <= 36'sb1000001111101100100011111111110;
            sine_reg0   <= 36'sb100000000001000100000000000111101001;
        end
        12373: begin
            cosine_reg0 <= 36'sb1000010101111110011110011010011;
            sine_reg0   <= 36'sb100000000001000101101000010110010101;
        end
        12374: begin
            cosine_reg0 <= 36'sb1000011100010000011000100000011;
            sine_reg0   <= 36'sb100000000001000111010001110011111011;
        end
        12375: begin
            cosine_reg0 <= 36'sb1000100010100010010010010001100;
            sine_reg0   <= 36'sb100000000001001000111100100000011100;
        end
        12376: begin
            cosine_reg0 <= 36'sb1000101000110100001011101101101;
            sine_reg0   <= 36'sb100000000001001010101000011011111000;
        end
        12377: begin
            cosine_reg0 <= 36'sb1000101111000110000100110100011;
            sine_reg0   <= 36'sb100000000001001100010101100110001101;
        end
        12378: begin
            cosine_reg0 <= 36'sb1000110101010111111101100101101;
            sine_reg0   <= 36'sb100000000001001110000011111111011101;
        end
        12379: begin
            cosine_reg0 <= 36'sb1000111011101001110110000001001;
            sine_reg0   <= 36'sb100000000001001111110011100111100111;
        end
        12380: begin
            cosine_reg0 <= 36'sb1001000001111011101110000110100;
            sine_reg0   <= 36'sb100000000001010001100100011110101100;
        end
        12381: begin
            cosine_reg0 <= 36'sb1001001000001101100101110101101;
            sine_reg0   <= 36'sb100000000001010011010110100100101010;
        end
        12382: begin
            cosine_reg0 <= 36'sb1001001110011111011101001110001;
            sine_reg0   <= 36'sb100000000001010101001001111001100011;
        end
        12383: begin
            cosine_reg0 <= 36'sb1001010100110001010100010000000;
            sine_reg0   <= 36'sb100000000001010110111110011101010101;
        end
        12384: begin
            cosine_reg0 <= 36'sb1001011011000011001010111010110;
            sine_reg0   <= 36'sb100000000001011000110100010000000001;
        end
        12385: begin
            cosine_reg0 <= 36'sb1001100001010101000001001110011;
            sine_reg0   <= 36'sb100000000001011010101011010001100111;
        end
        12386: begin
            cosine_reg0 <= 36'sb1001100111100110110111001010011;
            sine_reg0   <= 36'sb100000000001011100100011100010000111;
        end
        12387: begin
            cosine_reg0 <= 36'sb1001101101111000101100101110110;
            sine_reg0   <= 36'sb100000000001011110011101000001100001;
        end
        12388: begin
            cosine_reg0 <= 36'sb1001110100001010100001111011001;
            sine_reg0   <= 36'sb100000000001100000010111101111110100;
        end
        12389: begin
            cosine_reg0 <= 36'sb1001111010011100010110101111010;
            sine_reg0   <= 36'sb100000000001100010010011101101000001;
        end
        12390: begin
            cosine_reg0 <= 36'sb1010000000101110001011001011000;
            sine_reg0   <= 36'sb100000000001100100010000111001000111;
        end
        12391: begin
            cosine_reg0 <= 36'sb1010000110111111111111001110000;
            sine_reg0   <= 36'sb100000000001100110001111010100000110;
        end
        12392: begin
            cosine_reg0 <= 36'sb1010001101010001110010111000000;
            sine_reg0   <= 36'sb100000000001101000001110111101111111;
        end
        12393: begin
            cosine_reg0 <= 36'sb1010010011100011100110001000111;
            sine_reg0   <= 36'sb100000000001101010001111110110110001;
        end
        12394: begin
            cosine_reg0 <= 36'sb1010011001110101011001000000010;
            sine_reg0   <= 36'sb100000000001101100010001111110011100;
        end
        12395: begin
            cosine_reg0 <= 36'sb1010100000000111001011011110000;
            sine_reg0   <= 36'sb100000000001101110010101010101000000;
        end
        12396: begin
            cosine_reg0 <= 36'sb1010100110011000111101100001111;
            sine_reg0   <= 36'sb100000000001110000011001111010011101;
        end
        12397: begin
            cosine_reg0 <= 36'sb1010101100101010101111001011100;
            sine_reg0   <= 36'sb100000000001110010011111101110110011;
        end
        12398: begin
            cosine_reg0 <= 36'sb1010110010111100100000011010111;
            sine_reg0   <= 36'sb100000000001110100100110110010000010;
        end
        12399: begin
            cosine_reg0 <= 36'sb1010111001001110010001001111100;
            sine_reg0   <= 36'sb100000000001110110101111000100001010;
        end
        12400: begin
            cosine_reg0 <= 36'sb1010111111100000000001101001010;
            sine_reg0   <= 36'sb100000000001111000111000100101001010;
        end
        12401: begin
            cosine_reg0 <= 36'sb1011000101110001110001100111111;
            sine_reg0   <= 36'sb100000000001111011000011010101000011;
        end
        12402: begin
            cosine_reg0 <= 36'sb1011001100000011100001001011010;
            sine_reg0   <= 36'sb100000000001111101001111010011110100;
        end
        12403: begin
            cosine_reg0 <= 36'sb1011010010010101010000010010111;
            sine_reg0   <= 36'sb100000000001111111011100100001011110;
        end
        12404: begin
            cosine_reg0 <= 36'sb1011011000100110111110111110110;
            sine_reg0   <= 36'sb100000000010000001101010111110000000;
        end
        12405: begin
            cosine_reg0 <= 36'sb1011011110111000101101001110100;
            sine_reg0   <= 36'sb100000000010000011111010101001011011;
        end
        12406: begin
            cosine_reg0 <= 36'sb1011100101001010011011000001111;
            sine_reg0   <= 36'sb100000000010000110001011100011101101;
        end
        12407: begin
            cosine_reg0 <= 36'sb1011101011011100001000011000110;
            sine_reg0   <= 36'sb100000000010001000011101101100111000;
        end
        12408: begin
            cosine_reg0 <= 36'sb1011110001101101110101010010110;
            sine_reg0   <= 36'sb100000000010001010110001000100111010;
        end
        12409: begin
            cosine_reg0 <= 36'sb1011110111111111100001101111110;
            sine_reg0   <= 36'sb100000000010001101000101101011110101;
        end
        12410: begin
            cosine_reg0 <= 36'sb1011111110010001001101101111011;
            sine_reg0   <= 36'sb100000000010001111011011100001100111;
        end
        12411: begin
            cosine_reg0 <= 36'sb1100000100100010111001010001100;
            sine_reg0   <= 36'sb100000000010010001110010100110010001;
        end
        12412: begin
            cosine_reg0 <= 36'sb1100001010110100100100010101111;
            sine_reg0   <= 36'sb100000000010010100001010111001110010;
        end
        12413: begin
            cosine_reg0 <= 36'sb1100010001000110001110111100001;
            sine_reg0   <= 36'sb100000000010010110100100011100001011;
        end
        12414: begin
            cosine_reg0 <= 36'sb1100010111010111111001000100010;
            sine_reg0   <= 36'sb100000000010011000111111001101011100;
        end
        12415: begin
            cosine_reg0 <= 36'sb1100011101101001100010101101110;
            sine_reg0   <= 36'sb100000000010011011011011001101100100;
        end
        12416: begin
            cosine_reg0 <= 36'sb1100100011111011001011111000100;
            sine_reg0   <= 36'sb100000000010011101111000011100100011;
        end
        12417: begin
            cosine_reg0 <= 36'sb1100101010001100110100100100010;
            sine_reg0   <= 36'sb100000000010100000010110111010011001;
        end
        12418: begin
            cosine_reg0 <= 36'sb1100110000011110011100110000111;
            sine_reg0   <= 36'sb100000000010100010110110100111000110;
        end
        12419: begin
            cosine_reg0 <= 36'sb1100110110110000000100011101111;
            sine_reg0   <= 36'sb100000000010100101010111100010101010;
        end
        12420: begin
            cosine_reg0 <= 36'sb1100111101000001101011101011010;
            sine_reg0   <= 36'sb100000000010100111111001101101000101;
        end
        12421: begin
            cosine_reg0 <= 36'sb1101000011010011010010011000101;
            sine_reg0   <= 36'sb100000000010101010011101000110010111;
        end
        12422: begin
            cosine_reg0 <= 36'sb1101001001100100111000100101111;
            sine_reg0   <= 36'sb100000000010101101000001101110100000;
        end
        12423: begin
            cosine_reg0 <= 36'sb1101001111110110011110010010101;
            sine_reg0   <= 36'sb100000000010101111100111100101011111;
        end
        12424: begin
            cosine_reg0 <= 36'sb1101010110001000000011011110101;
            sine_reg0   <= 36'sb100000000010110010001110101011010101;
        end
        12425: begin
            cosine_reg0 <= 36'sb1101011100011001101000001001110;
            sine_reg0   <= 36'sb100000000010110100110111000000000000;
        end
        12426: begin
            cosine_reg0 <= 36'sb1101100010101011001100010011110;
            sine_reg0   <= 36'sb100000000010110111100000100011100011;
        end
        12427: begin
            cosine_reg0 <= 36'sb1101101000111100101111111100010;
            sine_reg0   <= 36'sb100000000010111010001011010101111011;
        end
        12428: begin
            cosine_reg0 <= 36'sb1101101111001110010011000011010;
            sine_reg0   <= 36'sb100000000010111100110111010111001001;
        end
        12429: begin
            cosine_reg0 <= 36'sb1101110101011111110101101000010;
            sine_reg0   <= 36'sb100000000010111111100100100111001110;
        end
        12430: begin
            cosine_reg0 <= 36'sb1101111011110001010111101011000;
            sine_reg0   <= 36'sb100000000011000010010011000110001000;
        end
        12431: begin
            cosine_reg0 <= 36'sb1110000010000010111001001011100;
            sine_reg0   <= 36'sb100000000011000101000010110011111000;
        end
        12432: begin
            cosine_reg0 <= 36'sb1110001000010100011010001001011;
            sine_reg0   <= 36'sb100000000011000111110011110000011110;
        end
        12433: begin
            cosine_reg0 <= 36'sb1110001110100101111010100100011;
            sine_reg0   <= 36'sb100000000011001010100101111011111001;
        end
        12434: begin
            cosine_reg0 <= 36'sb1110010100110111011010011100010;
            sine_reg0   <= 36'sb100000000011001101011001010110001001;
        end
        12435: begin
            cosine_reg0 <= 36'sb1110011011001000111001110000110;
            sine_reg0   <= 36'sb100000000011010000001101111111001111;
        end
        12436: begin
            cosine_reg0 <= 36'sb1110100001011010011000100001110;
            sine_reg0   <= 36'sb100000000011010011000011110111001010;
        end
        12437: begin
            cosine_reg0 <= 36'sb1110100111101011110110101110111;
            sine_reg0   <= 36'sb100000000011010101111010111101111011;
        end
        12438: begin
            cosine_reg0 <= 36'sb1110101101111101010100010111111;
            sine_reg0   <= 36'sb100000000011011000110011010011100000;
        end
        12439: begin
            cosine_reg0 <= 36'sb1110110100001110110001011100101;
            sine_reg0   <= 36'sb100000000011011011101100110111111010;
        end
        12440: begin
            cosine_reg0 <= 36'sb1110111010100000001101111100110;
            sine_reg0   <= 36'sb100000000011011110100111101011001001;
        end
        12441: begin
            cosine_reg0 <= 36'sb1111000000110001101001111000001;
            sine_reg0   <= 36'sb100000000011100001100011101101001100;
        end
        12442: begin
            cosine_reg0 <= 36'sb1111000111000011000101001110011;
            sine_reg0   <= 36'sb100000000011100100100000111110000100;
        end
        12443: begin
            cosine_reg0 <= 36'sb1111001101010100011111111111100;
            sine_reg0   <= 36'sb100000000011100111011111011101110001;
        end
        12444: begin
            cosine_reg0 <= 36'sb1111010011100101111010001011000;
            sine_reg0   <= 36'sb100000000011101010011111001100010001;
        end
        12445: begin
            cosine_reg0 <= 36'sb1111011001110111010011110000110;
            sine_reg0   <= 36'sb100000000011101101100000001001100110;
        end
        12446: begin
            cosine_reg0 <= 36'sb1111100000001000101100110000100;
            sine_reg0   <= 36'sb100000000011110000100010010101110000;
        end
        12447: begin
            cosine_reg0 <= 36'sb1111100110011010000101001010000;
            sine_reg0   <= 36'sb100000000011110011100101110000101101;
        end
        12448: begin
            cosine_reg0 <= 36'sb1111101100101011011100111101000;
            sine_reg0   <= 36'sb100000000011110110101010011010011101;
        end
        12449: begin
            cosine_reg0 <= 36'sb1111110010111100110100001001010;
            sine_reg0   <= 36'sb100000000011111001110000010011000010;
        end
        12450: begin
            cosine_reg0 <= 36'sb1111111001001110001010101110100;
            sine_reg0   <= 36'sb100000000011111100110111011010011010;
        end
        12451: begin
            cosine_reg0 <= 36'sb1111111111011111100000101100101;
            sine_reg0   <= 36'sb100000000011111111111111110000100110;
        end
        12452: begin
            cosine_reg0 <= 36'sb10000000101110000110110000011010;
            sine_reg0   <= 36'sb100000000100000011001001010101100101;
        end
        12453: begin
            cosine_reg0 <= 36'sb10000001100000010001010110010001;
            sine_reg0   <= 36'sb100000000100000110010100001001010111;
        end
        12454: begin
            cosine_reg0 <= 36'sb10000010010010011011110111001001;
            sine_reg0   <= 36'sb100000000100001001100000001011111101;
        end
        12455: begin
            cosine_reg0 <= 36'sb10000011000100100110010010111111;
            sine_reg0   <= 36'sb100000000100001100101101011101010101;
        end
        12456: begin
            cosine_reg0 <= 36'sb10000011110110110000101001110010;
            sine_reg0   <= 36'sb100000000100001111111011111101100000;
        end
        12457: begin
            cosine_reg0 <= 36'sb10000100101000111010111011100000;
            sine_reg0   <= 36'sb100000000100010011001011101100011110;
        end
        12458: begin
            cosine_reg0 <= 36'sb10000101011011000101001000000110;
            sine_reg0   <= 36'sb100000000100010110011100101010001111;
        end
        12459: begin
            cosine_reg0 <= 36'sb10000110001101001111001111100011;
            sine_reg0   <= 36'sb100000000100011001101110110110110010;
        end
        12460: begin
            cosine_reg0 <= 36'sb10000110111111011001010001110101;
            sine_reg0   <= 36'sb100000000100011101000010010010001000;
        end
        12461: begin
            cosine_reg0 <= 36'sb10000111110001100011001110111010;
            sine_reg0   <= 36'sb100000000100100000010110111100010000;
        end
        12462: begin
            cosine_reg0 <= 36'sb10001000100011101101000110110000;
            sine_reg0   <= 36'sb100000000100100011101100110101001010;
        end
        12463: begin
            cosine_reg0 <= 36'sb10001001010101110110111001010101;
            sine_reg0   <= 36'sb100000000100100111000011111100110110;
        end
        12464: begin
            cosine_reg0 <= 36'sb10001010001000000000100110100111;
            sine_reg0   <= 36'sb100000000100101010011100010011010011;
        end
        12465: begin
            cosine_reg0 <= 36'sb10001010111010001010001110100100;
            sine_reg0   <= 36'sb100000000100101101110101111000100011;
        end
        12466: begin
            cosine_reg0 <= 36'sb10001011101100010011110001001010;
            sine_reg0   <= 36'sb100000000100110001010000101100100100;
        end
        12467: begin
            cosine_reg0 <= 36'sb10001100011110011101001110011000;
            sine_reg0   <= 36'sb100000000100110100101100101111010111;
        end
        12468: begin
            cosine_reg0 <= 36'sb10001101010000100110100110001011;
            sine_reg0   <= 36'sb100000000100111000001010000000111011;
        end
        12469: begin
            cosine_reg0 <= 36'sb10001110000010101111111000100010;
            sine_reg0   <= 36'sb100000000100111011101000100001010000;
        end
        12470: begin
            cosine_reg0 <= 36'sb10001110110100111001000101011010;
            sine_reg0   <= 36'sb100000000100111111001000010000010110;
        end
        12471: begin
            cosine_reg0 <= 36'sb10001111100111000010001100110010;
            sine_reg0   <= 36'sb100000000101000010101001001110001101;
        end
        12472: begin
            cosine_reg0 <= 36'sb10010000011001001011001110100111;
            sine_reg0   <= 36'sb100000000101000110001011011010110101;
        end
        12473: begin
            cosine_reg0 <= 36'sb10010001001011010100001010111000;
            sine_reg0   <= 36'sb100000000101001001101110110110001110;
        end
        12474: begin
            cosine_reg0 <= 36'sb10010001111101011101000001100011;
            sine_reg0   <= 36'sb100000000101001101010011100000010111;
        end
        12475: begin
            cosine_reg0 <= 36'sb10010010101111100101110010100110;
            sine_reg0   <= 36'sb100000000101010000111001011001010000;
        end
        12476: begin
            cosine_reg0 <= 36'sb10010011100001101110011101111111;
            sine_reg0   <= 36'sb100000000101010100100000100000111010;
        end
        12477: begin
            cosine_reg0 <= 36'sb10010100010011110111000011101100;
            sine_reg0   <= 36'sb100000000101011000001000110111010100;
        end
        12478: begin
            cosine_reg0 <= 36'sb10010101000101111111100011101010;
            sine_reg0   <= 36'sb100000000101011011110010011100011110;
        end
        12479: begin
            cosine_reg0 <= 36'sb10010101111000000111111101111001;
            sine_reg0   <= 36'sb100000000101011111011101010000010111;
        end
        12480: begin
            cosine_reg0 <= 36'sb10010110101010010000010010010110;
            sine_reg0   <= 36'sb100000000101100011001001010011000001;
        end
        12481: begin
            cosine_reg0 <= 36'sb10010111011100011000100001000000;
            sine_reg0   <= 36'sb100000000101100110110110100100011010;
        end
        12482: begin
            cosine_reg0 <= 36'sb10011000001110100000101001110011;
            sine_reg0   <= 36'sb100000000101101010100101000100100010;
        end
        12483: begin
            cosine_reg0 <= 36'sb10011001000000101000101100101111;
            sine_reg0   <= 36'sb100000000101101110010100110011011001;
        end
        12484: begin
            cosine_reg0 <= 36'sb10011001110010110000101001110010;
            sine_reg0   <= 36'sb100000000101110010000101110001000000;
        end
        12485: begin
            cosine_reg0 <= 36'sb10011010100100111000100000111001;
            sine_reg0   <= 36'sb100000000101110101110111111101010110;
        end
        12486: begin
            cosine_reg0 <= 36'sb10011011010111000000010010000011;
            sine_reg0   <= 36'sb100000000101111001101011011000011010;
        end
        12487: begin
            cosine_reg0 <= 36'sb10011100001001000111111101001101;
            sine_reg0   <= 36'sb100000000101111101100000000010001101;
        end
        12488: begin
            cosine_reg0 <= 36'sb10011100111011001111100010010110;
            sine_reg0   <= 36'sb100000000110000001010101111010101111;
        end
        12489: begin
            cosine_reg0 <= 36'sb10011101101101010111000001011100;
            sine_reg0   <= 36'sb100000000110000101001101000001111111;
        end
        12490: begin
            cosine_reg0 <= 36'sb10011110011111011110011010011101;
            sine_reg0   <= 36'sb100000000110001001000101010111111101;
        end
        12491: begin
            cosine_reg0 <= 36'sb10011111010001100101101101010110;
            sine_reg0   <= 36'sb100000000110001100111110111100101010;
        end
        12492: begin
            cosine_reg0 <= 36'sb10100000000011101100111010000111;
            sine_reg0   <= 36'sb100000000110010000111001110000000100;
        end
        12493: begin
            cosine_reg0 <= 36'sb10100000110101110100000000101101;
            sine_reg0   <= 36'sb100000000110010100110101110010001100;
        end
        12494: begin
            cosine_reg0 <= 36'sb10100001100111111011000001000110;
            sine_reg0   <= 36'sb100000000110011000110011000011000010;
        end
        12495: begin
            cosine_reg0 <= 36'sb10100010011010000001111011010000;
            sine_reg0   <= 36'sb100000000110011100110001100010100101;
        end
        12496: begin
            cosine_reg0 <= 36'sb10100011001100001000101111001001;
            sine_reg0   <= 36'sb100000000110100000110001010000110101;
        end
        12497: begin
            cosine_reg0 <= 36'sb10100011111110001111011100110000;
            sine_reg0   <= 36'sb100000000110100100110010001101110011;
        end
        12498: begin
            cosine_reg0 <= 36'sb10100100110000010110000100000010;
            sine_reg0   <= 36'sb100000000110101000110100011001011110;
        end
        12499: begin
            cosine_reg0 <= 36'sb10100101100010011100100100111110;
            sine_reg0   <= 36'sb100000000110101100110111110011110101;
        end
        12500: begin
            cosine_reg0 <= 36'sb10100110010100100010111111100001;
            sine_reg0   <= 36'sb100000000110110000111100011100111010;
        end
        12501: begin
            cosine_reg0 <= 36'sb10100111000110101001010011101010;
            sine_reg0   <= 36'sb100000000110110101000010010100101010;
        end
        12502: begin
            cosine_reg0 <= 36'sb10100111111000101111100001010110;
            sine_reg0   <= 36'sb100000000110111001001001011011001000;
        end
        12503: begin
            cosine_reg0 <= 36'sb10101000101010110101101000100100;
            sine_reg0   <= 36'sb100000000110111101010001110000010001;
        end
        12504: begin
            cosine_reg0 <= 36'sb10101001011100111011101001010010;
            sine_reg0   <= 36'sb100000000111000001011011010100000111;
        end
        12505: begin
            cosine_reg0 <= 36'sb10101010001111000001100011011110;
            sine_reg0   <= 36'sb100000000111000101100110000110101000;
        end
        12506: begin
            cosine_reg0 <= 36'sb10101011000001000111010111000110;
            sine_reg0   <= 36'sb100000000111001001110010000111110101;
        end
        12507: begin
            cosine_reg0 <= 36'sb10101011110011001101000100001000;
            sine_reg0   <= 36'sb100000000111001101111111010111101110;
        end
        12508: begin
            cosine_reg0 <= 36'sb10101100100101010010101010100010;
            sine_reg0   <= 36'sb100000000111010010001101110110010010;
        end
        12509: begin
            cosine_reg0 <= 36'sb10101101010111011000001010010010;
            sine_reg0   <= 36'sb100000000111010110011101100011100001;
        end
        12510: begin
            cosine_reg0 <= 36'sb10101110001001011101100011010111;
            sine_reg0   <= 36'sb100000000111011010101110011111011100;
        end
        12511: begin
            cosine_reg0 <= 36'sb10101110111011100010110101101110;
            sine_reg0   <= 36'sb100000000111011111000000101010000001;
        end
        12512: begin
            cosine_reg0 <= 36'sb10101111101101101000000001010101;
            sine_reg0   <= 36'sb100000000111100011010100000011010010;
        end
        12513: begin
            cosine_reg0 <= 36'sb10110000011111101101000110001010;
            sine_reg0   <= 36'sb100000000111100111101000101011001100;
        end
        12514: begin
            cosine_reg0 <= 36'sb10110001010001110010000100001100;
            sine_reg0   <= 36'sb100000000111101011111110100001110010;
        end
        12515: begin
            cosine_reg0 <= 36'sb10110010000011110110111011011001;
            sine_reg0   <= 36'sb100000000111110000010101100111000001;
        end
        12516: begin
            cosine_reg0 <= 36'sb10110010110101111011101011101110;
            sine_reg0   <= 36'sb100000000111110100101101111010111011;
        end
        12517: begin
            cosine_reg0 <= 36'sb10110011101000000000010101001011;
            sine_reg0   <= 36'sb100000000111111001000111011101011111;
        end
        12518: begin
            cosine_reg0 <= 36'sb10110100011010000100110111101011;
            sine_reg0   <= 36'sb100000000111111101100010001110101100;
        end
        12519: begin
            cosine_reg0 <= 36'sb10110101001100001001010011001111;
            sine_reg0   <= 36'sb100000001000000001111110001110100011;
        end
        12520: begin
            cosine_reg0 <= 36'sb10110101111110001101100111110100;
            sine_reg0   <= 36'sb100000001000000110011011011101000011;
        end
        12521: begin
            cosine_reg0 <= 36'sb10110110110000010001110101010111;
            sine_reg0   <= 36'sb100000001000001010111001111010001101;
        end
        12522: begin
            cosine_reg0 <= 36'sb10110111100010010101111011111000;
            sine_reg0   <= 36'sb100000001000001111011001100101111111;
        end
        12523: begin
            cosine_reg0 <= 36'sb10111000010100011001111011010100;
            sine_reg0   <= 36'sb100000001000010011111010100000011011;
        end
        12524: begin
            cosine_reg0 <= 36'sb10111001000110011101110011101001;
            sine_reg0   <= 36'sb100000001000011000011100101001011111;
        end
        12525: begin
            cosine_reg0 <= 36'sb10111001111000100001100100110101;
            sine_reg0   <= 36'sb100000001000011101000000000001001100;
        end
        12526: begin
            cosine_reg0 <= 36'sb10111010101010100101001110110111;
            sine_reg0   <= 36'sb100000001000100001100100100111100010;
        end
        12527: begin
            cosine_reg0 <= 36'sb10111011011100101000110001101100;
            sine_reg0   <= 36'sb100000001000100110001010011100011111;
        end
        12528: begin
            cosine_reg0 <= 36'sb10111100001110101100001101010011;
            sine_reg0   <= 36'sb100000001000101010110001100000000101;
        end
        12529: begin
            cosine_reg0 <= 36'sb10111101000000101111100001101001;
            sine_reg0   <= 36'sb100000001000101111011001110010010010;
        end
        12530: begin
            cosine_reg0 <= 36'sb10111101110010110010101110101101;
            sine_reg0   <= 36'sb100000001000110100000011010011000111;
        end
        12531: begin
            cosine_reg0 <= 36'sb10111110100100110101110100011100;
            sine_reg0   <= 36'sb100000001000111000101110000010100011;
        end
        12532: begin
            cosine_reg0 <= 36'sb10111111010110111000110010110110;
            sine_reg0   <= 36'sb100000001000111101011010000000100111;
        end
        12533: begin
            cosine_reg0 <= 36'sb11000000001000111011101001110111;
            sine_reg0   <= 36'sb100000001001000010000111001101010010;
        end
        12534: begin
            cosine_reg0 <= 36'sb11000000111010111110011001011110;
            sine_reg0   <= 36'sb100000001001000110110101101000100100;
        end
        12535: begin
            cosine_reg0 <= 36'sb11000001101101000001000001101001;
            sine_reg0   <= 36'sb100000001001001011100101010010011101;
        end
        12536: begin
            cosine_reg0 <= 36'sb11000010011111000011100010010110;
            sine_reg0   <= 36'sb100000001001010000010110001010111100;
        end
        12537: begin
            cosine_reg0 <= 36'sb11000011010001000101111011100011;
            sine_reg0   <= 36'sb100000001001010101001000010010000010;
        end
        12538: begin
            cosine_reg0 <= 36'sb11000100000011001000001101001111;
            sine_reg0   <= 36'sb100000001001011001111011100111101101;
        end
        12539: begin
            cosine_reg0 <= 36'sb11000100110101001010010111010110;
            sine_reg0   <= 36'sb100000001001011110110000001011111111;
        end
        12540: begin
            cosine_reg0 <= 36'sb11000101100111001100011001111000;
            sine_reg0   <= 36'sb100000001001100011100101111110110111;
        end
        12541: begin
            cosine_reg0 <= 36'sb11000110011001001110010100110011;
            sine_reg0   <= 36'sb100000001001101000011101000000010100;
        end
        12542: begin
            cosine_reg0 <= 36'sb11000111001011010000001000000100;
            sine_reg0   <= 36'sb100000001001101101010101010000010111;
        end
        12543: begin
            cosine_reg0 <= 36'sb11000111111101010001110011101001;
            sine_reg0   <= 36'sb100000001001110010001110101110111111;
        end
        12544: begin
            cosine_reg0 <= 36'sb11001000101111010011010111100001;
            sine_reg0   <= 36'sb100000001001110111001001011100001101;
        end
        12545: begin
            cosine_reg0 <= 36'sb11001001100001010100110011101010;
            sine_reg0   <= 36'sb100000001001111100000101010111111111;
        end
        12546: begin
            cosine_reg0 <= 36'sb11001010010011010110001000000010;
            sine_reg0   <= 36'sb100000001010000001000010100010010110;
        end
        12547: begin
            cosine_reg0 <= 36'sb11001011000101010111010100100110;
            sine_reg0   <= 36'sb100000001010000110000000111011010001;
        end
        12548: begin
            cosine_reg0 <= 36'sb11001011110111011000011001010101;
            sine_reg0   <= 36'sb100000001010001011000000100010110001;
        end
        12549: begin
            cosine_reg0 <= 36'sb11001100101001011001010110001110;
            sine_reg0   <= 36'sb100000001010010000000001011000110101;
        end
        12550: begin
            cosine_reg0 <= 36'sb11001101011011011010001011001101;
            sine_reg0   <= 36'sb100000001010010101000011011101011100;
        end
        12551: begin
            cosine_reg0 <= 36'sb11001110001101011010111000010001;
            sine_reg0   <= 36'sb100000001010011010000110110000101000;
        end
        12552: begin
            cosine_reg0 <= 36'sb11001110111111011011011101011001;
            sine_reg0   <= 36'sb100000001010011111001011010010010111;
        end
        12553: begin
            cosine_reg0 <= 36'sb11001111110001011011111010100010;
            sine_reg0   <= 36'sb100000001010100100010001000010101010;
        end
        12554: begin
            cosine_reg0 <= 36'sb11010000100011011100001111101010;
            sine_reg0   <= 36'sb100000001010101001011000000001011111;
        end
        12555: begin
            cosine_reg0 <= 36'sb11010001010101011100011100110000;
            sine_reg0   <= 36'sb100000001010101110100000001110111000;
        end
        12556: begin
            cosine_reg0 <= 36'sb11010010000111011100100001110001;
            sine_reg0   <= 36'sb100000001010110011101001101010110011;
        end
        12557: begin
            cosine_reg0 <= 36'sb11010010111001011100011110101100;
            sine_reg0   <= 36'sb100000001010111000110100010101010001;
        end
        12558: begin
            cosine_reg0 <= 36'sb11010011101011011100010011011110;
            sine_reg0   <= 36'sb100000001010111110000000001110010010;
        end
        12559: begin
            cosine_reg0 <= 36'sb11010100011101011100000000000110;
            sine_reg0   <= 36'sb100000001011000011001101010101110100;
        end
        12560: begin
            cosine_reg0 <= 36'sb11010101001111011011100100100010;
            sine_reg0   <= 36'sb100000001011001000011011101011111000;
        end
        12561: begin
            cosine_reg0 <= 36'sb11010110000001011011000000110000;
            sine_reg0   <= 36'sb100000001011001101101011010000011111;
        end
        12562: begin
            cosine_reg0 <= 36'sb11010110110011011010010100101110;
            sine_reg0   <= 36'sb100000001011010010111100000011100111;
        end
        12563: begin
            cosine_reg0 <= 36'sb11010111100101011001100000011001;
            sine_reg0   <= 36'sb100000001011011000001110000101010000;
        end
        12564: begin
            cosine_reg0 <= 36'sb11011000010111011000100011110001;
            sine_reg0   <= 36'sb100000001011011101100001010101011010;
        end
        12565: begin
            cosine_reg0 <= 36'sb11011001001001010111011110110011;
            sine_reg0   <= 36'sb100000001011100010110101110100000101;
        end
        12566: begin
            cosine_reg0 <= 36'sb11011001111011010110010001011101;
            sine_reg0   <= 36'sb100000001011101000001011100001010001;
        end
        12567: begin
            cosine_reg0 <= 36'sb11011010101101010100111011101101;
            sine_reg0   <= 36'sb100000001011101101100010011100111110;
        end
        12568: begin
            cosine_reg0 <= 36'sb11011011011111010011011101100010;
            sine_reg0   <= 36'sb100000001011110010111010100111001011;
        end
        12569: begin
            cosine_reg0 <= 36'sb11011100010001010001110110111001;
            sine_reg0   <= 36'sb100000001011111000010011111111111000;
        end
        12570: begin
            cosine_reg0 <= 36'sb11011101000011010000000111110000;
            sine_reg0   <= 36'sb100000001011111101101110100111000101;
        end
        12571: begin
            cosine_reg0 <= 36'sb11011101110101001110010000000111;
            sine_reg0   <= 36'sb100000001100000011001010011100110010;
        end
        12572: begin
            cosine_reg0 <= 36'sb11011110100111001100001111111001;
            sine_reg0   <= 36'sb100000001100001000100111100000111110;
        end
        12573: begin
            cosine_reg0 <= 36'sb11011111011001001010000111000111;
            sine_reg0   <= 36'sb100000001100001110000101110011101001;
        end
        12574: begin
            cosine_reg0 <= 36'sb11100000001011000111110101101101;
            sine_reg0   <= 36'sb100000001100010011100101010100110100;
        end
        12575: begin
            cosine_reg0 <= 36'sb11100000111101000101011011101011;
            sine_reg0   <= 36'sb100000001100011001000110000100011101;
        end
        12576: begin
            cosine_reg0 <= 36'sb11100001101111000010111000111101;
            sine_reg0   <= 36'sb100000001100011110101000000010100110;
        end
        12577: begin
            cosine_reg0 <= 36'sb11100010100001000000001101100010;
            sine_reg0   <= 36'sb100000001100100100001011001111001100;
        end
        12578: begin
            cosine_reg0 <= 36'sb11100011010010111101011001011000;
            sine_reg0   <= 36'sb100000001100101001101111101010010001;
        end
        12579: begin
            cosine_reg0 <= 36'sb11100100000100111010011100011110;
            sine_reg0   <= 36'sb100000001100101111010101010011110100;
        end
        12580: begin
            cosine_reg0 <= 36'sb11100100110110110111010110110001;
            sine_reg0   <= 36'sb100000001100110100111100001011110100;
        end
        12581: begin
            cosine_reg0 <= 36'sb11100101101000110100001000001111;
            sine_reg0   <= 36'sb100000001100111010100100010010010011;
        end
        12582: begin
            cosine_reg0 <= 36'sb11100110011010110000110000110110;
            sine_reg0   <= 36'sb100000001101000000001101100111001110;
        end
        12583: begin
            cosine_reg0 <= 36'sb11100111001100101101010000100101;
            sine_reg0   <= 36'sb100000001101000101111000001010100111;
        end
        12584: begin
            cosine_reg0 <= 36'sb11100111111110101001100111011001;
            sine_reg0   <= 36'sb100000001101001011100011111100011101;
        end
        12585: begin
            cosine_reg0 <= 36'sb11101000110000100101110101010001;
            sine_reg0   <= 36'sb100000001101010001010000111100101111;
        end
        12586: begin
            cosine_reg0 <= 36'sb11101001100010100001111010001011;
            sine_reg0   <= 36'sb100000001101010110111111001011011110;
        end
        12587: begin
            cosine_reg0 <= 36'sb11101010010100011101110110000101;
            sine_reg0   <= 36'sb100000001101011100101110101000101001;
        end
        12588: begin
            cosine_reg0 <= 36'sb11101011000110011001101000111100;
            sine_reg0   <= 36'sb100000001101100010011111010100010000;
        end
        12589: begin
            cosine_reg0 <= 36'sb11101011111000010101010010101111;
            sine_reg0   <= 36'sb100000001101101000010001001110010011;
        end
        12590: begin
            cosine_reg0 <= 36'sb11101100101010010000110011011101;
            sine_reg0   <= 36'sb100000001101101110000100010110110010;
        end
        12591: begin
            cosine_reg0 <= 36'sb11101101011100001100001011000010;
            sine_reg0   <= 36'sb100000001101110011111000101101101100;
        end
        12592: begin
            cosine_reg0 <= 36'sb11101110001110000111011001011101;
            sine_reg0   <= 36'sb100000001101111001101110010011000001;
        end
        12593: begin
            cosine_reg0 <= 36'sb11101111000000000010011110101101;
            sine_reg0   <= 36'sb100000001101111111100101000110110001;
        end
        12594: begin
            cosine_reg0 <= 36'sb11101111110001111101011010101111;
            sine_reg0   <= 36'sb100000001110000101011101001000111100;
        end
        12595: begin
            cosine_reg0 <= 36'sb11110000100011111000001101100001;
            sine_reg0   <= 36'sb100000001110001011010110011001100010;
        end
        12596: begin
            cosine_reg0 <= 36'sb11110001010101110010110111000010;
            sine_reg0   <= 36'sb100000001110010001010000111000100001;
        end
        12597: begin
            cosine_reg0 <= 36'sb11110010000111101101010111001111;
            sine_reg0   <= 36'sb100000001110010111001100100101111011;
        end
        12598: begin
            cosine_reg0 <= 36'sb11110010111001100111101110000111;
            sine_reg0   <= 36'sb100000001110011101001001100001101110;
        end
        12599: begin
            cosine_reg0 <= 36'sb11110011101011100001111011101000;
            sine_reg0   <= 36'sb100000001110100011000111101011111011;
        end
        12600: begin
            cosine_reg0 <= 36'sb11110100011101011011111111101111;
            sine_reg0   <= 36'sb100000001110101001000111000100100010;
        end
        12601: begin
            cosine_reg0 <= 36'sb11110101001111010101111010011011;
            sine_reg0   <= 36'sb100000001110101111000111101011100001;
        end
        12602: begin
            cosine_reg0 <= 36'sb11110110000001001111101011101010;
            sine_reg0   <= 36'sb100000001110110101001001100000111001;
        end
        12603: begin
            cosine_reg0 <= 36'sb11110110110011001001010011011010;
            sine_reg0   <= 36'sb100000001110111011001100100100101010;
        end
        12604: begin
            cosine_reg0 <= 36'sb11110111100101000010110001101001;
            sine_reg0   <= 36'sb100000001111000001010000110110110100;
        end
        12605: begin
            cosine_reg0 <= 36'sb11111000010110111100000110010101;
            sine_reg0   <= 36'sb100000001111000111010110010111010101;
        end
        12606: begin
            cosine_reg0 <= 36'sb11111001001000110101010001011101;
            sine_reg0   <= 36'sb100000001111001101011101000110001111;
        end
        12607: begin
            cosine_reg0 <= 36'sb11111001111010101110010010111101;
            sine_reg0   <= 36'sb100000001111010011100101000011100000;
        end
        12608: begin
            cosine_reg0 <= 36'sb11111010101100100111001010110101;
            sine_reg0   <= 36'sb100000001111011001101110001111001001;
        end
        12609: begin
            cosine_reg0 <= 36'sb11111011011110011111111001000011;
            sine_reg0   <= 36'sb100000001111011111111000101001001000;
        end
        12610: begin
            cosine_reg0 <= 36'sb11111100010000011000011101100011;
            sine_reg0   <= 36'sb100000001111100110000100010001011111;
        end
        12611: begin
            cosine_reg0 <= 36'sb11111101000010010000111000010110;
            sine_reg0   <= 36'sb100000001111101100010001001000001101;
        end
        12612: begin
            cosine_reg0 <= 36'sb11111101110100001001001001011000;
            sine_reg0   <= 36'sb100000001111110010011111001101010001;
        end
        12613: begin
            cosine_reg0 <= 36'sb11111110100110000001010000101000;
            sine_reg0   <= 36'sb100000001111111000101110100000101100;
        end
        12614: begin
            cosine_reg0 <= 36'sb11111111010111111001001110000100;
            sine_reg0   <= 36'sb100000001111111110111111000010011100;
        end
        12615: begin
            cosine_reg0 <= 36'sb100000000001001110001000001101001;
            sine_reg0   <= 36'sb100000010000000101010000110010100010;
        end
        12616: begin
            cosine_reg0 <= 36'sb100000000111011101000101011010111;
            sine_reg0   <= 36'sb100000010000001011100011110000111110;
        end
        12617: begin
            cosine_reg0 <= 36'sb100000001101101100000001011001010;
            sine_reg0   <= 36'sb100000010000010001110111111101110000;
        end
        12618: begin
            cosine_reg0 <= 36'sb100000010011111010111100001000010;
            sine_reg0   <= 36'sb100000010000011000001101011000110110;
        end
        12619: begin
            cosine_reg0 <= 36'sb100000011010001001110101100111100;
            sine_reg0   <= 36'sb100000010000011110100100000010010001;
        end
        12620: begin
            cosine_reg0 <= 36'sb100000100000011000101101110110110;
            sine_reg0   <= 36'sb100000010000100100111011111010000000;
        end
        12621: begin
            cosine_reg0 <= 36'sb100000100110100111100100110101111;
            sine_reg0   <= 36'sb100000010000101011010101000000000100;
        end
        12622: begin
            cosine_reg0 <= 36'sb100000101100110110011010100100100;
            sine_reg0   <= 36'sb100000010000110001101111010100011101;
        end
        12623: begin
            cosine_reg0 <= 36'sb100000110011000101001111000010011;
            sine_reg0   <= 36'sb100000010000111000001010110111001000;
        end
        12624: begin
            cosine_reg0 <= 36'sb100000111001010100000010001111100;
            sine_reg0   <= 36'sb100000010000111110100111101000001000;
        end
        12625: begin
            cosine_reg0 <= 36'sb100000111111100010110100001011010;
            sine_reg0   <= 36'sb100000010001000101000101100111011011;
        end
        12626: begin
            cosine_reg0 <= 36'sb100001000101110001100100110101110;
            sine_reg0   <= 36'sb100000010001001011100100110101000001;
        end
        12627: begin
            cosine_reg0 <= 36'sb100001001100000000010100001110100;
            sine_reg0   <= 36'sb100000010001010010000101010000111010;
        end
        12628: begin
            cosine_reg0 <= 36'sb100001010010001111000010010101011;
            sine_reg0   <= 36'sb100000010001011000100110111011000101;
        end
        12629: begin
            cosine_reg0 <= 36'sb100001011000011101101111001010010;
            sine_reg0   <= 36'sb100000010001011111001001110011100011;
        end
        12630: begin
            cosine_reg0 <= 36'sb100001011110101100011010101100101;
            sine_reg0   <= 36'sb100000010001100101101101111010010010;
        end
        12631: begin
            cosine_reg0 <= 36'sb100001100100111011000100111100011;
            sine_reg0   <= 36'sb100000010001101100010011001111010100;
        end
        12632: begin
            cosine_reg0 <= 36'sb100001101011001001101101111001011;
            sine_reg0   <= 36'sb100000010001110010111001110010100111;
        end
        12633: begin
            cosine_reg0 <= 36'sb100001110001011000010101100011010;
            sine_reg0   <= 36'sb100000010001111001100001100100001100;
        end
        12634: begin
            cosine_reg0 <= 36'sb100001110111100110111011111001110;
            sine_reg0   <= 36'sb100000010010000000001010100100000010;
        end
        12635: begin
            cosine_reg0 <= 36'sb100001111101110101100000111100110;
            sine_reg0   <= 36'sb100000010010000110110100110010001000;
        end
        12636: begin
            cosine_reg0 <= 36'sb100010000100000100000100101011111;
            sine_reg0   <= 36'sb100000010010001101100000001110011111;
        end
        12637: begin
            cosine_reg0 <= 36'sb100010001010010010100111000111000;
            sine_reg0   <= 36'sb100000010010010100001100111001000110;
        end
        12638: begin
            cosine_reg0 <= 36'sb100010010000100001001000001101111;
            sine_reg0   <= 36'sb100000010010011010111010110001111110;
        end
        12639: begin
            cosine_reg0 <= 36'sb100010010110101111101000000000001;
            sine_reg0   <= 36'sb100000010010100001101001111001000101;
        end
        12640: begin
            cosine_reg0 <= 36'sb100010011100111110000110011101110;
            sine_reg0   <= 36'sb100000010010101000011010001110011100;
        end
        12641: begin
            cosine_reg0 <= 36'sb100010100011001100100011100110010;
            sine_reg0   <= 36'sb100000010010101111001011110010000001;
        end
        12642: begin
            cosine_reg0 <= 36'sb100010101001011010111111011001100;
            sine_reg0   <= 36'sb100000010010110101111110100011110110;
        end
        12643: begin
            cosine_reg0 <= 36'sb100010101111101001011001110111010;
            sine_reg0   <= 36'sb100000010010111100110010100011111010;
        end
        12644: begin
            cosine_reg0 <= 36'sb100010110101110111110010111111011;
            sine_reg0   <= 36'sb100000010011000011100111110010001100;
        end
        12645: begin
            cosine_reg0 <= 36'sb100010111100000110001010110001011;
            sine_reg0   <= 36'sb100000010011001010011110001110101101;
        end
        12646: begin
            cosine_reg0 <= 36'sb100011000010010100100001001101010;
            sine_reg0   <= 36'sb100000010011010001010101111001011011;
        end
        12647: begin
            cosine_reg0 <= 36'sb100011001000100010110110010010110;
            sine_reg0   <= 36'sb100000010011011000001110110010010111;
        end
        12648: begin
            cosine_reg0 <= 36'sb100011001110110001001010000001100;
            sine_reg0   <= 36'sb100000010011011111001000111001100001;
        end
        12649: begin
            cosine_reg0 <= 36'sb100011010100111111011100011001010;
            sine_reg0   <= 36'sb100000010011100110000100001110110111;
        end
        12650: begin
            cosine_reg0 <= 36'sb100011011011001101101101011001111;
            sine_reg0   <= 36'sb100000010011101101000000110010011011;
        end
        12651: begin
            cosine_reg0 <= 36'sb100011100001011011111101000011001;
            sine_reg0   <= 36'sb100000010011110011111110100100001011;
        end
        12652: begin
            cosine_reg0 <= 36'sb100011100111101010001011010100110;
            sine_reg0   <= 36'sb100000010011111010111101100100000111;
        end
        12653: begin
            cosine_reg0 <= 36'sb100011101101111000011000001110100;
            sine_reg0   <= 36'sb100000010100000001111101110010010000;
        end
        12654: begin
            cosine_reg0 <= 36'sb100011110100000110100011110000000;
            sine_reg0   <= 36'sb100000010100001000111111001110100100;
        end
        12655: begin
            cosine_reg0 <= 36'sb100011111010010100101101111001010;
            sine_reg0   <= 36'sb100000010100010000000001111001000100;
        end
        12656: begin
            cosine_reg0 <= 36'sb100100000000100010110110101001111;
            sine_reg0   <= 36'sb100000010100010111000101110001101111;
        end
        12657: begin
            cosine_reg0 <= 36'sb100100000110110000111110000001101;
            sine_reg0   <= 36'sb100000010100011110001010111000100101;
        end
        12658: begin
            cosine_reg0 <= 36'sb100100001100111111000100000000010;
            sine_reg0   <= 36'sb100000010100100101010001001101100110;
        end
        12659: begin
            cosine_reg0 <= 36'sb100100010011001101001000100101101;
            sine_reg0   <= 36'sb100000010100101100011000110000110010;
        end
        12660: begin
            cosine_reg0 <= 36'sb100100011001011011001011110001011;
            sine_reg0   <= 36'sb100000010100110011100001100010000111;
        end
        12661: begin
            cosine_reg0 <= 36'sb100100011111101001001101100011010;
            sine_reg0   <= 36'sb100000010100111010101011100001100111;
        end
        12662: begin
            cosine_reg0 <= 36'sb100100100101110111001101111011010;
            sine_reg0   <= 36'sb100000010101000001110110101111010000;
        end
        12663: begin
            cosine_reg0 <= 36'sb100100101100000101001100111000111;
            sine_reg0   <= 36'sb100000010101001001000011001011000010;
        end
        12664: begin
            cosine_reg0 <= 36'sb100100110010010011001010011100000;
            sine_reg0   <= 36'sb100000010101010000010000110100111110;
        end
        12665: begin
            cosine_reg0 <= 36'sb100100111000100001000110100100010;
            sine_reg0   <= 36'sb100000010101010111011111101101000010;
        end
        12666: begin
            cosine_reg0 <= 36'sb100100111110101111000001010001101;
            sine_reg0   <= 36'sb100000010101011110101111110011001111;
        end
        12667: begin
            cosine_reg0 <= 36'sb100101000100111100111010100011110;
            sine_reg0   <= 36'sb100000010101100110000001000111100100;
        end
        12668: begin
            cosine_reg0 <= 36'sb100101001011001010110010011010011;
            sine_reg0   <= 36'sb100000010101101101010011101010000001;
        end
        12669: begin
            cosine_reg0 <= 36'sb100101010001011000101000110101010;
            sine_reg0   <= 36'sb100000010101110100100111011010100110;
        end
        12670: begin
            cosine_reg0 <= 36'sb100101010111100110011101110100001;
            sine_reg0   <= 36'sb100000010101111011111100011001010010;
        end
        12671: begin
            cosine_reg0 <= 36'sb100101011101110100010001010110111;
            sine_reg0   <= 36'sb100000010110000011010010100110000101;
        end
        12672: begin
            cosine_reg0 <= 36'sb100101100100000010000011011101001;
            sine_reg0   <= 36'sb100000010110001010101010000000111111;
        end
        12673: begin
            cosine_reg0 <= 36'sb100101101010001111110100000110101;
            sine_reg0   <= 36'sb100000010110010010000010101001111111;
        end
        12674: begin
            cosine_reg0 <= 36'sb100101110000011101100011010011011;
            sine_reg0   <= 36'sb100000010110011001011100100001000110;
        end
        12675: begin
            cosine_reg0 <= 36'sb100101110110101011010001000010111;
            sine_reg0   <= 36'sb100000010110100000110111100110010011;
        end
        12676: begin
            cosine_reg0 <= 36'sb100101111100111000111101010101000;
            sine_reg0   <= 36'sb100000010110101000010011111001100101;
        end
        12677: begin
            cosine_reg0 <= 36'sb100110000011000110101000001001011;
            sine_reg0   <= 36'sb100000010110101111110001011010111101;
        end
        12678: begin
            cosine_reg0 <= 36'sb100110001001010100010001100000000;
            sine_reg0   <= 36'sb100000010110110111010000001010011010;
        end
        12679: begin
            cosine_reg0 <= 36'sb100110001111100001111001011000011;
            sine_reg0   <= 36'sb100000010110111110110000000111111100;
        end
        12680: begin
            cosine_reg0 <= 36'sb100110010101101111011111110010100;
            sine_reg0   <= 36'sb100000010111000110010001010011100010;
        end
        12681: begin
            cosine_reg0 <= 36'sb100110011011111101000100101110000;
            sine_reg0   <= 36'sb100000010111001101110011101101001101;
        end
        12682: begin
            cosine_reg0 <= 36'sb100110100010001010101000001010101;
            sine_reg0   <= 36'sb100000010111010101010111010100111100;
        end
        12683: begin
            cosine_reg0 <= 36'sb100110101000011000001010001000010;
            sine_reg0   <= 36'sb100000010111011100111100001010101110;
        end
        12684: begin
            cosine_reg0 <= 36'sb100110101110100101101010100110100;
            sine_reg0   <= 36'sb100000010111100100100010001110100011;
        end
        12685: begin
            cosine_reg0 <= 36'sb100110110100110011001001100101010;
            sine_reg0   <= 36'sb100000010111101100001001100000011100;
        end
        12686: begin
            cosine_reg0 <= 36'sb100110111011000000100111000100001;
            sine_reg0   <= 36'sb100000010111110011110010000000010111;
        end
        12687: begin
            cosine_reg0 <= 36'sb100111000001001110000011000011000;
            sine_reg0   <= 36'sb100000010111111011011011101110010101;
        end
        12688: begin
            cosine_reg0 <= 36'sb100111000111011011011101100001101;
            sine_reg0   <= 36'sb100000011000000011000110101010010110;
        end
        12689: begin
            cosine_reg0 <= 36'sb100111001101101000110110011111101;
            sine_reg0   <= 36'sb100000011000001010110010110100011000;
        end
        12690: begin
            cosine_reg0 <= 36'sb100111010011110110001101111101000;
            sine_reg0   <= 36'sb100000011000010010100000001100011011;
        end
        12691: begin
            cosine_reg0 <= 36'sb100111011010000011100011111001011;
            sine_reg0   <= 36'sb100000011000011010001110110010100000;
        end
        12692: begin
            cosine_reg0 <= 36'sb100111100000010000111000010100011;
            sine_reg0   <= 36'sb100000011000100001111110100110100110;
        end
        12693: begin
            cosine_reg0 <= 36'sb100111100110011110001011001110000;
            sine_reg0   <= 36'sb100000011000101001101111101000101101;
        end
        12694: begin
            cosine_reg0 <= 36'sb100111101100101011011100100110000;
            sine_reg0   <= 36'sb100000011000110001100001111000110100;
        end
        12695: begin
            cosine_reg0 <= 36'sb100111110010111000101100011011111;
            sine_reg0   <= 36'sb100000011000111001010101010110111011;
        end
        12696: begin
            cosine_reg0 <= 36'sb100111111001000101111010101111110;
            sine_reg0   <= 36'sb100000011001000001001010000011000010;
        end
        12697: begin
            cosine_reg0 <= 36'sb100111111111010011000111100001000;
            sine_reg0   <= 36'sb100000011001001000111111111101001001;
        end
        12698: begin
            cosine_reg0 <= 36'sb101000000101100000010010101111110;
            sine_reg0   <= 36'sb100000011001010000110111000101001110;
        end
        12699: begin
            cosine_reg0 <= 36'sb101000001011101101011100011011100;
            sine_reg0   <= 36'sb100000011001011000101111011011010011;
        end
        12700: begin
            cosine_reg0 <= 36'sb101000010001111010100100100100001;
            sine_reg0   <= 36'sb100000011001100000101000111111010110;
        end
        12701: begin
            cosine_reg0 <= 36'sb101000011000000111101011001001011;
            sine_reg0   <= 36'sb100000011001101000100011110001011000;
        end
        12702: begin
            cosine_reg0 <= 36'sb101000011110010100110000001010111;
            sine_reg0   <= 36'sb100000011001110000011111110001010111;
        end
        12703: begin
            cosine_reg0 <= 36'sb101000100100100001110011101000101;
            sine_reg0   <= 36'sb100000011001111000011100111111010100;
        end
        12704: begin
            cosine_reg0 <= 36'sb101000101010101110110101100010010;
            sine_reg0   <= 36'sb100000011010000000011011011011001111;
        end
        12705: begin
            cosine_reg0 <= 36'sb101000110000111011110101110111101;
            sine_reg0   <= 36'sb100000011010001000011011000101000110;
        end
        12706: begin
            cosine_reg0 <= 36'sb101000110111001000110100101000010;
            sine_reg0   <= 36'sb100000011010010000011011111100111011;
        end
        12707: begin
            cosine_reg0 <= 36'sb101000111101010101110001110100010;
            sine_reg0   <= 36'sb100000011010011000011110000010101100;
        end
        12708: begin
            cosine_reg0 <= 36'sb101001000011100010101101011011000;
            sine_reg0   <= 36'sb100000011010100000100001010110011001;
        end
        12709: begin
            cosine_reg0 <= 36'sb101001001001101111100111011100100;
            sine_reg0   <= 36'sb100000011010101000100101111000000001;
        end
        12710: begin
            cosine_reg0 <= 36'sb101001001111111100011111111000100;
            sine_reg0   <= 36'sb100000011010110000101011100111100110;
        end
        12711: begin
            cosine_reg0 <= 36'sb101001010110001001010110101110110;
            sine_reg0   <= 36'sb100000011010111000110010100101000101;
        end
        12712: begin
            cosine_reg0 <= 36'sb101001011100010110001011111110111;
            sine_reg0   <= 36'sb100000011011000000111010110000100000;
        end
        12713: begin
            cosine_reg0 <= 36'sb101001100010100010111111101000111;
            sine_reg0   <= 36'sb100000011011001001000100001001110101;
        end
        12714: begin
            cosine_reg0 <= 36'sb101001101000101111110001101100010;
            sine_reg0   <= 36'sb100000011011010001001110110001000100;
        end
        12715: begin
            cosine_reg0 <= 36'sb101001101110111100100010001001000;
            sine_reg0   <= 36'sb100000011011011001011010100110001101;
        end
        12716: begin
            cosine_reg0 <= 36'sb101001110101001001010000111110110;
            sine_reg0   <= 36'sb100000011011100001100111101001010000;
        end
        12717: begin
            cosine_reg0 <= 36'sb101001111011010101111110001101010;
            sine_reg0   <= 36'sb100000011011101001110101111010001100;
        end
        12718: begin
            cosine_reg0 <= 36'sb101010000001100010101001110100011;
            sine_reg0   <= 36'sb100000011011110010000101011001000001;
        end
        12719: begin
            cosine_reg0 <= 36'sb101010000111101111010011110011110;
            sine_reg0   <= 36'sb100000011011111010010110000101101111;
        end
        12720: begin
            cosine_reg0 <= 36'sb101010001101111011111100001011001;
            sine_reg0   <= 36'sb100000011100000010101000000000010101;
        end
        12721: begin
            cosine_reg0 <= 36'sb101010010100001000100010111010100;
            sine_reg0   <= 36'sb100000011100001010111011001000110100;
        end
        12722: begin
            cosine_reg0 <= 36'sb101010011010010101001000000001011;
            sine_reg0   <= 36'sb100000011100010011001111011111001010;
        end
        12723: begin
            cosine_reg0 <= 36'sb101010100000100001101011011111100;
            sine_reg0   <= 36'sb100000011100011011100101000011010111;
        end
        12724: begin
            cosine_reg0 <= 36'sb101010100110101110001101010100111;
            sine_reg0   <= 36'sb100000011100100011111011110101011100;
        end
        12725: begin
            cosine_reg0 <= 36'sb101010101100111010101101100001001;
            sine_reg0   <= 36'sb100000011100101100010011110101010111;
        end
        12726: begin
            cosine_reg0 <= 36'sb101010110011000111001100000100000;
            sine_reg0   <= 36'sb100000011100110100101101000011001001;
        end
        12727: begin
            cosine_reg0 <= 36'sb101010111001010011101000111101010;
            sine_reg0   <= 36'sb100000011100111101000111011110110001;
        end
        12728: begin
            cosine_reg0 <= 36'sb101010111111100000000100001100101;
            sine_reg0   <= 36'sb100000011101000101100011001000001110;
        end
        12729: begin
            cosine_reg0 <= 36'sb101011000101101100011101110010000;
            sine_reg0   <= 36'sb100000011101001101111111111111100001;
        end
        12730: begin
            cosine_reg0 <= 36'sb101011001011111000110101101101000;
            sine_reg0   <= 36'sb100000011101010110011110000100101010;
        end
        12731: begin
            cosine_reg0 <= 36'sb101011010010000101001011111101100;
            sine_reg0   <= 36'sb100000011101011110111101010111100111;
        end
        12732: begin
            cosine_reg0 <= 36'sb101011011000010001100000100011001;
            sine_reg0   <= 36'sb100000011101100111011101111000011000;
        end
        12733: begin
            cosine_reg0 <= 36'sb101011011110011101110011011101110;
            sine_reg0   <= 36'sb100000011101101111111111100110111110;
        end
        12734: begin
            cosine_reg0 <= 36'sb101011100100101010000100101101001;
            sine_reg0   <= 36'sb100000011101111000100010100011010111;
        end
        12735: begin
            cosine_reg0 <= 36'sb101011101010110110010100010001000;
            sine_reg0   <= 36'sb100000011110000001000110101101100100;
        end
        12736: begin
            cosine_reg0 <= 36'sb101011110001000010100010001001001;
            sine_reg0   <= 36'sb100000011110001001101100000101100101;
        end
        12737: begin
            cosine_reg0 <= 36'sb101011110111001110101110010101001;
            sine_reg0   <= 36'sb100000011110010010010010101011011000;
        end
        12738: begin
            cosine_reg0 <= 36'sb101011111101011010111000110101000;
            sine_reg0   <= 36'sb100000011110011010111010011110111101;
        end
        12739: begin
            cosine_reg0 <= 36'sb101100000011100111000001101000100;
            sine_reg0   <= 36'sb100000011110100011100011100000010101;
        end
        12740: begin
            cosine_reg0 <= 36'sb101100001001110011001000101111001;
            sine_reg0   <= 36'sb100000011110101100001101101111011111;
        end
        12741: begin
            cosine_reg0 <= 36'sb101100001111111111001110001001000;
            sine_reg0   <= 36'sb100000011110110100111001001100011010;
        end
        12742: begin
            cosine_reg0 <= 36'sb101100010110001011010001110101100;
            sine_reg0   <= 36'sb100000011110111101100101110111000110;
        end
        12743: begin
            cosine_reg0 <= 36'sb101100011100010111010011110100110;
            sine_reg0   <= 36'sb100000011111000110010011101111100011;
        end
        12744: begin
            cosine_reg0 <= 36'sb101100100010100011010100000110010;
            sine_reg0   <= 36'sb100000011111001111000010110101110001;
        end
        12745: begin
            cosine_reg0 <= 36'sb101100101000101111010010101001111;
            sine_reg0   <= 36'sb100000011111010111110011001001101111;
        end
        12746: begin
            cosine_reg0 <= 36'sb101100101110111011001111011111010;
            sine_reg0   <= 36'sb100000011111100000100100101011011100;
        end
        12747: begin
            cosine_reg0 <= 36'sb101100110101000111001010100110011;
            sine_reg0   <= 36'sb100000011111101001010111011010111001;
        end
        12748: begin
            cosine_reg0 <= 36'sb101100111011010011000011111110111;
            sine_reg0   <= 36'sb100000011111110010001011011000000110;
        end
        12749: begin
            cosine_reg0 <= 36'sb101101000001011110111011101000100;
            sine_reg0   <= 36'sb100000011111111011000000100011000001;
        end
        12750: begin
            cosine_reg0 <= 36'sb101101000111101010110001100011000;
            sine_reg0   <= 36'sb100000100000000011110110111011101010;
        end
        12751: begin
            cosine_reg0 <= 36'sb101101001101110110100101101110010;
            sine_reg0   <= 36'sb100000100000001100101110100010000010;
        end
        12752: begin
            cosine_reg0 <= 36'sb101101010100000010011000001001111;
            sine_reg0   <= 36'sb100000100000010101100111010110000111;
        end
        12753: begin
            cosine_reg0 <= 36'sb101101011010001110001000110101110;
            sine_reg0   <= 36'sb100000100000011110100001010111111010;
        end
        12754: begin
            cosine_reg0 <= 36'sb101101100000011001110111110001100;
            sine_reg0   <= 36'sb100000100000100111011100100111011010;
        end
        12755: begin
            cosine_reg0 <= 36'sb101101100110100101100100111101000;
            sine_reg0   <= 36'sb100000100000110000011001000100100111;
        end
        12756: begin
            cosine_reg0 <= 36'sb101101101100110001010000011000000;
            sine_reg0   <= 36'sb100000100000111001010110101111100000;
        end
        12757: begin
            cosine_reg0 <= 36'sb101101110010111100111010000010010;
            sine_reg0   <= 36'sb100000100001000010010101101000000110;
        end
        12758: begin
            cosine_reg0 <= 36'sb101101111001001000100001111011100;
            sine_reg0   <= 36'sb100000100001001011010101101110010111;
        end
        12759: begin
            cosine_reg0 <= 36'sb101101111111010100001000000011100;
            sine_reg0   <= 36'sb100000100001010100010111000010010011;
        end
        12760: begin
            cosine_reg0 <= 36'sb101110000101011111101100011010000;
            sine_reg0   <= 36'sb100000100001011101011001100011111010;
        end
        12761: begin
            cosine_reg0 <= 36'sb101110001011101011001110111110111;
            sine_reg0   <= 36'sb100000100001100110011101010011001101;
        end
        12762: begin
            cosine_reg0 <= 36'sb101110010001110110101111110001110;
            sine_reg0   <= 36'sb100000100001101111100010010000001001;
        end
        12763: begin
            cosine_reg0 <= 36'sb101110011000000010001110110010011;
            sine_reg0   <= 36'sb100000100001111000101000011010101111;
        end
        12764: begin
            cosine_reg0 <= 36'sb101110011110001101101100000000101;
            sine_reg0   <= 36'sb100000100010000001101111110010111111;
        end
        12765: begin
            cosine_reg0 <= 36'sb101110100100011001000111011100010;
            sine_reg0   <= 36'sb100000100010001010111000011000111001;
        end
        12766: begin
            cosine_reg0 <= 36'sb101110101010100100100001000100111;
            sine_reg0   <= 36'sb100000100010010100000010001100011011;
        end
        12767: begin
            cosine_reg0 <= 36'sb101110110000101111111000111010100;
            sine_reg0   <= 36'sb100000100010011101001101001101100110;
        end
        12768: begin
            cosine_reg0 <= 36'sb101110110110111011001110111100101;
            sine_reg0   <= 36'sb100000100010100110011001011100011001;
        end
        12769: begin
            cosine_reg0 <= 36'sb101110111101000110100011001011001;
            sine_reg0   <= 36'sb100000100010101111100110111000110100;
        end
        12770: begin
            cosine_reg0 <= 36'sb101111000011010001110101100101111;
            sine_reg0   <= 36'sb100000100010111000110101100010110110;
        end
        12771: begin
            cosine_reg0 <= 36'sb101111001001011101000110001100011;
            sine_reg0   <= 36'sb100000100011000010000101011010100000;
        end
        12772: begin
            cosine_reg0 <= 36'sb101111001111101000010100111110101;
            sine_reg0   <= 36'sb100000100011001011010110011111110000;
        end
        12773: begin
            cosine_reg0 <= 36'sb101111010101110011100001111100011;
            sine_reg0   <= 36'sb100000100011010100101000110010100111;
        end
        12774: begin
            cosine_reg0 <= 36'sb101111011011111110101101000101010;
            sine_reg0   <= 36'sb100000100011011101111100010011000100;
        end
        12775: begin
            cosine_reg0 <= 36'sb101111100010001001110110011001001;
            sine_reg0   <= 36'sb100000100011100111010001000001000110;
        end
        12776: begin
            cosine_reg0 <= 36'sb101111101000010100111101110111101;
            sine_reg0   <= 36'sb100000100011110000100110111100101110;
        end
        12777: begin
            cosine_reg0 <= 36'sb101111101110100000000011100000101;
            sine_reg0   <= 36'sb100000100011111001111110000101111011;
        end
        12778: begin
            cosine_reg0 <= 36'sb101111110100101011000111010011111;
            sine_reg0   <= 36'sb100000100100000011010110011100101101;
        end
        12779: begin
            cosine_reg0 <= 36'sb101111111010110110001001010001001;
            sine_reg0   <= 36'sb100000100100001100110000000001000011;
        end
        12780: begin
            cosine_reg0 <= 36'sb110000000001000001001001011000010;
            sine_reg0   <= 36'sb100000100100010110001010110010111100;
        end
        12781: begin
            cosine_reg0 <= 36'sb110000000111001100000111101000110;
            sine_reg0   <= 36'sb100000100100011111100110110010011010;
        end
        12782: begin
            cosine_reg0 <= 36'sb110000001101010111000100000010101;
            sine_reg0   <= 36'sb100000100100101001000011111111011010;
        end
        12783: begin
            cosine_reg0 <= 36'sb110000010011100001111110100101100;
            sine_reg0   <= 36'sb100000100100110010100010011001111110;
        end
        12784: begin
            cosine_reg0 <= 36'sb110000011001101100110111010001010;
            sine_reg0   <= 36'sb100000100100111100000010000010000100;
        end
        12785: begin
            cosine_reg0 <= 36'sb110000011111110111101110000101100;
            sine_reg0   <= 36'sb100000100101000101100010110111101011;
        end
        12786: begin
            cosine_reg0 <= 36'sb110000100110000010100011000010001;
            sine_reg0   <= 36'sb100000100101001111000100111010110101;
        end
        12787: begin
            cosine_reg0 <= 36'sb110000101100001101010110000110110;
            sine_reg0   <= 36'sb100000100101011000101000001011100000;
        end
        12788: begin
            cosine_reg0 <= 36'sb110000110010011000000111010011011;
            sine_reg0   <= 36'sb100000100101100010001100101001101100;
        end
        12789: begin
            cosine_reg0 <= 36'sb110000111000100010110110100111101;
            sine_reg0   <= 36'sb100000100101101011110010010101011001;
        end
        12790: begin
            cosine_reg0 <= 36'sb110000111110101101100100000011001;
            sine_reg0   <= 36'sb100000100101110101011001001110100110;
        end
        12791: begin
            cosine_reg0 <= 36'sb110001000100111000001111100101111;
            sine_reg0   <= 36'sb100000100101111111000001010101010011;
        end
        12792: begin
            cosine_reg0 <= 36'sb110001001011000010111001001111100;
            sine_reg0   <= 36'sb100000100110001000101010101001011111;
        end
        12793: begin
            cosine_reg0 <= 36'sb110001010001001101100000111111111;
            sine_reg0   <= 36'sb100000100110010010010101001011001010;
        end
        12794: begin
            cosine_reg0 <= 36'sb110001010111011000000110110110100;
            sine_reg0   <= 36'sb100000100110011100000000111010010101;
        end
        12795: begin
            cosine_reg0 <= 36'sb110001011101100010101010110011100;
            sine_reg0   <= 36'sb100000100110100101101101110110111101;
        end
        12796: begin
            cosine_reg0 <= 36'sb110001100011101101001100110110011;
            sine_reg0   <= 36'sb100000100110101111011100000001000100;
        end
        12797: begin
            cosine_reg0 <= 36'sb110001101001110111101100111111000;
            sine_reg0   <= 36'sb100000100110111001001011011000101000;
        end
        12798: begin
            cosine_reg0 <= 36'sb110001110000000010001011001101001;
            sine_reg0   <= 36'sb100000100111000010111011111101101010;
        end
        12799: begin
            cosine_reg0 <= 36'sb110001110110001100100111100000100;
            sine_reg0   <= 36'sb100000100111001100101101110000001000;
        end
        12800: begin
            cosine_reg0 <= 36'sb110001111100010111000001111000110;
            sine_reg0   <= 36'sb100000100111010110100000110000000011;
        end
        12801: begin
            cosine_reg0 <= 36'sb110010000010100001011010010101111;
            sine_reg0   <= 36'sb100000100111100000010100111101011010;
        end
        12802: begin
            cosine_reg0 <= 36'sb110010001000101011110000110111101;
            sine_reg0   <= 36'sb100000100111101010001010011000001101;
        end
        12803: begin
            cosine_reg0 <= 36'sb110010001110110110000101011101100;
            sine_reg0   <= 36'sb100000100111110100000001000000011011;
        end
        12804: begin
            cosine_reg0 <= 36'sb110010010101000000011000000111100;
            sine_reg0   <= 36'sb100000100111111101111000110110000101;
        end
        12805: begin
            cosine_reg0 <= 36'sb110010011011001010101000110101011;
            sine_reg0   <= 36'sb100000101000000111110001111001001001;
        end
        12806: begin
            cosine_reg0 <= 36'sb110010100001010100110111100110110;
            sine_reg0   <= 36'sb100000101000010001101100001001100111;
        end
        12807: begin
            cosine_reg0 <= 36'sb110010100111011111000100011011100;
            sine_reg0   <= 36'sb100000101000011011100111100111011111;
        end
        12808: begin
            cosine_reg0 <= 36'sb110010101101101001001111010011011;
            sine_reg0   <= 36'sb100000101000100101100100010010110000;
        end
        12809: begin
            cosine_reg0 <= 36'sb110010110011110011011000001110001;
            sine_reg0   <= 36'sb100000101000101111100010001011011011;
        end
        12810: begin
            cosine_reg0 <= 36'sb110010111001111101011111001011100;
            sine_reg0   <= 36'sb100000101000111001100001010001011110;
        end
        12811: begin
            cosine_reg0 <= 36'sb110011000000000111100100001011010;
            sine_reg0   <= 36'sb100000101001000011100001100100111010;
        end
        12812: begin
            cosine_reg0 <= 36'sb110011000110010001100111001101001;
            sine_reg0   <= 36'sb100000101001001101100011000101101101;
        end
        12813: begin
            cosine_reg0 <= 36'sb110011001100011011101000010001000;
            sine_reg0   <= 36'sb100000101001010111100101110011111000;
        end
        12814: begin
            cosine_reg0 <= 36'sb110011010010100101100111010110100;
            sine_reg0   <= 36'sb100000101001100001101001101111011010;
        end
        12815: begin
            cosine_reg0 <= 36'sb110011011000101111100100011101100;
            sine_reg0   <= 36'sb100000101001101011101110111000010011;
        end
        12816: begin
            cosine_reg0 <= 36'sb110011011110111001011111100101110;
            sine_reg0   <= 36'sb100000101001110101110101001110100011;
        end
        12817: begin
            cosine_reg0 <= 36'sb110011100101000011011000101110111;
            sine_reg0   <= 36'sb100000101001111111111100110010001000;
        end
        12818: begin
            cosine_reg0 <= 36'sb110011101011001101001111111000110;
            sine_reg0   <= 36'sb100000101010001010000101100011000011;
        end
        12819: begin
            cosine_reg0 <= 36'sb110011110001010111000101000011001;
            sine_reg0   <= 36'sb100000101010010100001111100001010011;
        end
        12820: begin
            cosine_reg0 <= 36'sb110011110111100000111000001101110;
            sine_reg0   <= 36'sb100000101010011110011010101100111001;
        end
        12821: begin
            cosine_reg0 <= 36'sb110011111101101010101001011000011;
            sine_reg0   <= 36'sb100000101010101000100111000101110010;
        end
        12822: begin
            cosine_reg0 <= 36'sb110100000011110100011000100010111;
            sine_reg0   <= 36'sb100000101010110010110100101100000000;
        end
        12823: begin
            cosine_reg0 <= 36'sb110100001001111110000101101100111;
            sine_reg0   <= 36'sb100000101010111101000011011111100001;
        end
        12824: begin
            cosine_reg0 <= 36'sb110100010000000111110000110110001;
            sine_reg0   <= 36'sb100000101011000111010011100000010101;
        end
        12825: begin
            cosine_reg0 <= 36'sb110100010110010001011001111110100;
            sine_reg0   <= 36'sb100000101011010001100100101110011100;
        end
        12826: begin
            cosine_reg0 <= 36'sb110100011100011011000001000101110;
            sine_reg0   <= 36'sb100000101011011011110111001001110110;
        end
        12827: begin
            cosine_reg0 <= 36'sb110100100010100100100110001011101;
            sine_reg0   <= 36'sb100000101011100110001010110010100010;
        end
        12828: begin
            cosine_reg0 <= 36'sb110100101000101110001001001111110;
            sine_reg0   <= 36'sb100000101011110000011111101000100000;
        end
        12829: begin
            cosine_reg0 <= 36'sb110100101110110111101010010010000;
            sine_reg0   <= 36'sb100000101011111010110101101011101110;
        end
        12830: begin
            cosine_reg0 <= 36'sb110100110101000001001001010010010;
            sine_reg0   <= 36'sb100000101100000101001100111100001110;
        end
        12831: begin
            cosine_reg0 <= 36'sb110100111011001010100110010000001;
            sine_reg0   <= 36'sb100000101100001111100101011001111110;
        end
        12832: begin
            cosine_reg0 <= 36'sb110101000001010100000001001011011;
            sine_reg0   <= 36'sb100000101100011001111111000100111110;
        end
        12833: begin
            cosine_reg0 <= 36'sb110101000111011101011010000011110;
            sine_reg0   <= 36'sb100000101100100100011001111101001110;
        end
        12834: begin
            cosine_reg0 <= 36'sb110101001101100110110000111001001;
            sine_reg0   <= 36'sb100000101100101110110110000010101101;
        end
        12835: begin
            cosine_reg0 <= 36'sb110101010011110000000101101011010;
            sine_reg0   <= 36'sb100000101100111001010011010101011011;
        end
        12836: begin
            cosine_reg0 <= 36'sb110101011001111001011000011001110;
            sine_reg0   <= 36'sb100000101101000011110001110101011000;
        end
        12837: begin
            cosine_reg0 <= 36'sb110101100000000010101001000100100;
            sine_reg0   <= 36'sb100000101101001110010001100010100010;
        end
        12838: begin
            cosine_reg0 <= 36'sb110101100110001011110111101011011;
            sine_reg0   <= 36'sb100000101101011000110010011100111010;
        end
        12839: begin
            cosine_reg0 <= 36'sb110101101100010101000100001101111;
            sine_reg0   <= 36'sb100000101101100011010100100100100000;
        end
        12840: begin
            cosine_reg0 <= 36'sb110101110010011110001110101011111;
            sine_reg0   <= 36'sb100000101101101101110111111001010010;
        end
        12841: begin
            cosine_reg0 <= 36'sb110101111000100111010111000101010;
            sine_reg0   <= 36'sb100000101101111000011100011011010000;
        end
        12842: begin
            cosine_reg0 <= 36'sb110101111110110000011101011001101;
            sine_reg0   <= 36'sb100000101110000011000010001010011011;
        end
        12843: begin
            cosine_reg0 <= 36'sb110110000100111001100001101000110;
            sine_reg0   <= 36'sb100000101110001101101001000110110010;
        end
        12844: begin
            cosine_reg0 <= 36'sb110110001011000010100011110010100;
            sine_reg0   <= 36'sb100000101110011000010001010000010011;
        end
        12845: begin
            cosine_reg0 <= 36'sb110110010001001011100011110110101;
            sine_reg0   <= 36'sb100000101110100010111010100110111111;
        end
        12846: begin
            cosine_reg0 <= 36'sb110110010111010100100001110100110;
            sine_reg0   <= 36'sb100000101110101101100101001010110110;
        end
        12847: begin
            cosine_reg0 <= 36'sb110110011101011101011101101100110;
            sine_reg0   <= 36'sb100000101110111000010000111011110111;
        end
        12848: begin
            cosine_reg0 <= 36'sb110110100011100110010111011110100;
            sine_reg0   <= 36'sb100000101111000010111101111010000001;
        end
        12849: begin
            cosine_reg0 <= 36'sb110110101001101111001111001001100;
            sine_reg0   <= 36'sb100000101111001101101100000101010101;
        end
        12850: begin
            cosine_reg0 <= 36'sb110110101111111000000100101101110;
            sine_reg0   <= 36'sb100000101111011000011011011101110001;
        end
        12851: begin
            cosine_reg0 <= 36'sb110110110110000000111000001010111;
            sine_reg0   <= 36'sb100000101111100011001100000011010101;
        end
        12852: begin
            cosine_reg0 <= 36'sb110110111100001001101001100000101;
            sine_reg0   <= 36'sb100000101111101101111101110110000010;
        end
        12853: begin
            cosine_reg0 <= 36'sb110111000010010010011000101110111;
            sine_reg0   <= 36'sb100000101111111000110000110101110101;
        end
        12854: begin
            cosine_reg0 <= 36'sb110111001000011011000101110101010;
            sine_reg0   <= 36'sb100000110000000011100101000010110000;
        end
        12855: begin
            cosine_reg0 <= 36'sb110111001110100011110000110011110;
            sine_reg0   <= 36'sb100000110000001110011010011100110010;
        end
        12856: begin
            cosine_reg0 <= 36'sb110111010100101100011001101001111;
            sine_reg0   <= 36'sb100000110000011001010001000011111010;
        end
        12857: begin
            cosine_reg0 <= 36'sb110111011010110101000000010111100;
            sine_reg0   <= 36'sb100000110000100100001000111000001000;
        end
        12858: begin
            cosine_reg0 <= 36'sb110111100000111101100100111100011;
            sine_reg0   <= 36'sb100000110000101111000001111001011011;
        end
        12859: begin
            cosine_reg0 <= 36'sb110111100111000110000111011000010;
            sine_reg0   <= 36'sb100000110000111001111100000111110011;
        end
        12860: begin
            cosine_reg0 <= 36'sb110111101101001110100111101011000;
            sine_reg0   <= 36'sb100000110001000100110111100011010000;
        end
        12861: begin
            cosine_reg0 <= 36'sb110111110011010111000101110100010;
            sine_reg0   <= 36'sb100000110001001111110100001011110001;
        end
        12862: begin
            cosine_reg0 <= 36'sb110111111001011111100001110011111;
            sine_reg0   <= 36'sb100000110001011010110010000001010101;
        end
        12863: begin
            cosine_reg0 <= 36'sb110111111111100111111011101001100;
            sine_reg0   <= 36'sb100000110001100101110001000011111101;
        end
        12864: begin
            cosine_reg0 <= 36'sb111000000101110000010011010101000;
            sine_reg0   <= 36'sb100000110001110000110001010011101000;
        end
        12865: begin
            cosine_reg0 <= 36'sb111000001011111000101000110110000;
            sine_reg0   <= 36'sb100000110001111011110010110000010101;
        end
        12866: begin
            cosine_reg0 <= 36'sb111000010010000000111100001100100;
            sine_reg0   <= 36'sb100000110010000110110101011010000100;
        end
        12867: begin
            cosine_reg0 <= 36'sb111000011000001001001101011000001;
            sine_reg0   <= 36'sb100000110010010001111001010000110101;
        end
        12868: begin
            cosine_reg0 <= 36'sb111000011110010001011100011000101;
            sine_reg0   <= 36'sb100000110010011100111110010100100111;
        end
        12869: begin
            cosine_reg0 <= 36'sb111000100100011001101001001101110;
            sine_reg0   <= 36'sb100000110010101000000100100101011010;
        end
        12870: begin
            cosine_reg0 <= 36'sb111000101010100001110011110111010;
            sine_reg0   <= 36'sb100000110010110011001100000011001101;
        end
        12871: begin
            cosine_reg0 <= 36'sb111000110000101001111100010101000;
            sine_reg0   <= 36'sb100000110010111110010100101110000000;
        end
        12872: begin
            cosine_reg0 <= 36'sb111000110110110010000010100110110;
            sine_reg0   <= 36'sb100000110011001001011110100101110010;
        end
        12873: begin
            cosine_reg0 <= 36'sb111000111100111010000110101100001;
            sine_reg0   <= 36'sb100000110011010100101001101010100100;
        end
        12874: begin
            cosine_reg0 <= 36'sb111001000011000010001000100101000;
            sine_reg0   <= 36'sb100000110011011111110101111100010100;
        end
        12875: begin
            cosine_reg0 <= 36'sb111001001001001010001000010001001;
            sine_reg0   <= 36'sb100000110011101011000011011011000010;
        end
        12876: begin
            cosine_reg0 <= 36'sb111001001111010010000101110000010;
            sine_reg0   <= 36'sb100000110011110110010010000110101110;
        end
        12877: begin
            cosine_reg0 <= 36'sb111001010101011010000001000010001;
            sine_reg0   <= 36'sb100000110100000001100001111111010111;
        end
        12878: begin
            cosine_reg0 <= 36'sb111001011011100001111010000110101;
            sine_reg0   <= 36'sb100000110100001100110011000100111110;
        end
        12879: begin
            cosine_reg0 <= 36'sb111001100001101001110000111101011;
            sine_reg0   <= 36'sb100000110100011000000101010111100000;
        end
        12880: begin
            cosine_reg0 <= 36'sb111001100111110001100101100110001;
            sine_reg0   <= 36'sb100000110100100011011000110110111111;
        end
        12881: begin
            cosine_reg0 <= 36'sb111001101101111001011000000000110;
            sine_reg0   <= 36'sb100000110100101110101101100011011001;
        end
        12882: begin
            cosine_reg0 <= 36'sb111001110100000001001000001101000;
            sine_reg0   <= 36'sb100000110100111010000011011100101110;
        end
        12883: begin
            cosine_reg0 <= 36'sb111001111010001000110110001010100;
            sine_reg0   <= 36'sb100000110101000101011010100010111110;
        end
        12884: begin
            cosine_reg0 <= 36'sb111010000000010000100001111001001;
            sine_reg0   <= 36'sb100000110101010000110010110110001001;
        end
        12885: begin
            cosine_reg0 <= 36'sb111010000110011000001011011000110;
            sine_reg0   <= 36'sb100000110101011100001100010110001101;
        end
        12886: begin
            cosine_reg0 <= 36'sb111010001100011111110010101000111;
            sine_reg0   <= 36'sb100000110101100111100111000011001010;
        end
        12887: begin
            cosine_reg0 <= 36'sb111010010010100111010111101001100;
            sine_reg0   <= 36'sb100000110101110011000010111101000001;
        end
        12888: begin
            cosine_reg0 <= 36'sb111010011000101110111010011010011;
            sine_reg0   <= 36'sb100000110101111110100000000011101111;
        end
        12889: begin
            cosine_reg0 <= 36'sb111010011110110110011010111011000;
            sine_reg0   <= 36'sb100000110110001001111110010111010110;
        end
        12890: begin
            cosine_reg0 <= 36'sb111010100100111101111001001011100;
            sine_reg0   <= 36'sb100000110110010101011101110111110101;
        end
        12891: begin
            cosine_reg0 <= 36'sb111010101011000101010101001011011;
            sine_reg0   <= 36'sb100000110110100000111110100101001011;
        end
        12892: begin
            cosine_reg0 <= 36'sb111010110001001100101110111010100;
            sine_reg0   <= 36'sb100000110110101100100000011111010111;
        end
        12893: begin
            cosine_reg0 <= 36'sb111010110111010100000110011000101;
            sine_reg0   <= 36'sb100000110110111000000011100110011010;
        end
        12894: begin
            cosine_reg0 <= 36'sb111010111101011011011011100101100;
            sine_reg0   <= 36'sb100000110111000011100111111010010011;
        end
        12895: begin
            cosine_reg0 <= 36'sb111011000011100010101110100000111;
            sine_reg0   <= 36'sb100000110111001111001101011011000000;
        end
        12896: begin
            cosine_reg0 <= 36'sb111011001001101001111111001010100;
            sine_reg0   <= 36'sb100000110111011010110100001000100011;
        end
        12897: begin
            cosine_reg0 <= 36'sb111011001111110001001101100010010;
            sine_reg0   <= 36'sb100000110111100110011100000010111011;
        end
        12898: begin
            cosine_reg0 <= 36'sb111011010101111000011001100111110;
            sine_reg0   <= 36'sb100000110111110010000101001010000110;
        end
        12899: begin
            cosine_reg0 <= 36'sb111011011011111111100011011010111;
            sine_reg0   <= 36'sb100000110111111101101111011110000101;
        end
        12900: begin
            cosine_reg0 <= 36'sb111011100010000110101010111011011;
            sine_reg0   <= 36'sb100000111000001001011010111110111000;
        end
        12901: begin
            cosine_reg0 <= 36'sb111011101000001101110000001001000;
            sine_reg0   <= 36'sb100000111000010101000111101100011100;
        end
        12902: begin
            cosine_reg0 <= 36'sb111011101110010100110011000011011;
            sine_reg0   <= 36'sb100000111000100000110101100110110100;
        end
        12903: begin
            cosine_reg0 <= 36'sb111011110100011011110011101010100;
            sine_reg0   <= 36'sb100000111000101100100100101101111101;
        end
        12904: begin
            cosine_reg0 <= 36'sb111011111010100010110001111110000;
            sine_reg0   <= 36'sb100000111000111000010101000001110111;
        end
        12905: begin
            cosine_reg0 <= 36'sb111100000000101001101101111101101;
            sine_reg0   <= 36'sb100000111001000100000110100010100010;
        end
        12906: begin
            cosine_reg0 <= 36'sb111100000110110000100111101001010;
            sine_reg0   <= 36'sb100000111001001111111001001111111110;
        end
        12907: begin
            cosine_reg0 <= 36'sb111100001100110111011111000000100;
            sine_reg0   <= 36'sb100000111001011011101101001010001001;
        end
        12908: begin
            cosine_reg0 <= 36'sb111100010010111110010100000011010;
            sine_reg0   <= 36'sb100000111001100111100010010001000100;
        end
        12909: begin
            cosine_reg0 <= 36'sb111100011001000101000110110001010;
            sine_reg0   <= 36'sb100000111001110011011000100100101111;
        end
        12910: begin
            cosine_reg0 <= 36'sb111100011111001011110111001010001;
            sine_reg0   <= 36'sb100000111001111111010000000101001000;
        end
        12911: begin
            cosine_reg0 <= 36'sb111100100101010010100101001101111;
            sine_reg0   <= 36'sb100000111010001011001000110010001111;
        end
        12912: begin
            cosine_reg0 <= 36'sb111100101011011001010000111100001;
            sine_reg0   <= 36'sb100000111010010111000010101100000011;
        end
        12913: begin
            cosine_reg0 <= 36'sb111100110001011111111010010100101;
            sine_reg0   <= 36'sb100000111010100010111101110010100101;
        end
        12914: begin
            cosine_reg0 <= 36'sb111100110111100110100001010111001;
            sine_reg0   <= 36'sb100000111010101110111010000101110100;
        end
        12915: begin
            cosine_reg0 <= 36'sb111100111101101101000110000011100;
            sine_reg0   <= 36'sb100000111010111010110111100101101111;
        end
        12916: begin
            cosine_reg0 <= 36'sb111101000011110011101000011001100;
            sine_reg0   <= 36'sb100000111011000110110110010010010110;
        end
        12917: begin
            cosine_reg0 <= 36'sb111101001001111010001000011000110;
            sine_reg0   <= 36'sb100000111011010010110110001011101000;
        end
        12918: begin
            cosine_reg0 <= 36'sb111101010000000000100110000001001;
            sine_reg0   <= 36'sb100000111011011110110111010001100101;
        end
        12919: begin
            cosine_reg0 <= 36'sb111101010110000111000001010010011;
            sine_reg0   <= 36'sb100000111011101010111001100100001101;
        end
        12920: begin
            cosine_reg0 <= 36'sb111101011100001101011010001100011;
            sine_reg0   <= 36'sb100000111011110110111101000011011111;
        end
        12921: begin
            cosine_reg0 <= 36'sb111101100010010011110000101110101;
            sine_reg0   <= 36'sb100000111100000011000001101111011010;
        end
        12922: begin
            cosine_reg0 <= 36'sb111101101000011010000100111001001;
            sine_reg0   <= 36'sb100000111100001111000111100111111110;
        end
        12923: begin
            cosine_reg0 <= 36'sb111101101110100000010110101011100;
            sine_reg0   <= 36'sb100000111100011011001110101101001011;
        end
        12924: begin
            cosine_reg0 <= 36'sb111101110100100110100110000101101;
            sine_reg0   <= 36'sb100000111100100111010110111111000000;
        end
        12925: begin
            cosine_reg0 <= 36'sb111101111010101100110011000111001;
            sine_reg0   <= 36'sb100000111100110011100000011101011101;
        end
        12926: begin
            cosine_reg0 <= 36'sb111110000000110010111101101111111;
            sine_reg0   <= 36'sb100000111100111111101011001000100001;
        end
        12927: begin
            cosine_reg0 <= 36'sb111110000110111001000101111111110;
            sine_reg0   <= 36'sb100000111101001011110111000000001011;
        end
        12928: begin
            cosine_reg0 <= 36'sb111110001100111111001011110110010;
            sine_reg0   <= 36'sb100000111101011000000100000100011100;
        end
        12929: begin
            cosine_reg0 <= 36'sb111110010011000101001111010011010;
            sine_reg0   <= 36'sb100000111101100100010010010101010011;
        end
        12930: begin
            cosine_reg0 <= 36'sb111110011001001011010000010110101;
            sine_reg0   <= 36'sb100000111101110000100001110010101111;
        end
        12931: begin
            cosine_reg0 <= 36'sb111110011111010001001111000000000;
            sine_reg0   <= 36'sb100000111101111100110010011100110000;
        end
        12932: begin
            cosine_reg0 <= 36'sb111110100101010111001011001111010;
            sine_reg0   <= 36'sb100000111110001001000100010011010101;
        end
        12933: begin
            cosine_reg0 <= 36'sb111110101011011101000101000100000;
            sine_reg0   <= 36'sb100000111110010101010111010110011111;
        end
        12934: begin
            cosine_reg0 <= 36'sb111110110001100010111100011110001;
            sine_reg0   <= 36'sb100000111110100001101011100110001011;
        end
        12935: begin
            cosine_reg0 <= 36'sb111110110111101000110001011101011;
            sine_reg0   <= 36'sb100000111110101110000001000010011011;
        end
        12936: begin
            cosine_reg0 <= 36'sb111110111101101110100100000001100;
            sine_reg0   <= 36'sb100000111110111010010111101011001101;
        end
        12937: begin
            cosine_reg0 <= 36'sb111111000011110100010100001010010;
            sine_reg0   <= 36'sb100000111111000110101111100000100001;
        end
        12938: begin
            cosine_reg0 <= 36'sb111111001001111010000001110111011;
            sine_reg0   <= 36'sb100000111111010011001000100010010111;
        end
        12939: begin
            cosine_reg0 <= 36'sb111111001111111111101101001000110;
            sine_reg0   <= 36'sb100000111111011111100010110000101110;
        end
        12940: begin
            cosine_reg0 <= 36'sb111111010110000101010101111110000;
            sine_reg0   <= 36'sb100000111111101011111110001011100101;
        end
        12941: begin
            cosine_reg0 <= 36'sb111111011100001010111100010110111;
            sine_reg0   <= 36'sb100000111111111000011010110010111100;
        end
        12942: begin
            cosine_reg0 <= 36'sb111111100010010000100000010011011;
            sine_reg0   <= 36'sb100001000000000100111000100110110011;
        end
        12943: begin
            cosine_reg0 <= 36'sb111111101000010110000001110011000;
            sine_reg0   <= 36'sb100001000000010001010111100111001001;
        end
        12944: begin
            cosine_reg0 <= 36'sb111111101110011011100000110101110;
            sine_reg0   <= 36'sb100001000000011101110111110011111110;
        end
        12945: begin
            cosine_reg0 <= 36'sb111111110100100000111101011011001;
            sine_reg0   <= 36'sb100001000000101010011001001101010001;
        end
        12946: begin
            cosine_reg0 <= 36'sb111111111010100110010111100011001;
            sine_reg0   <= 36'sb100001000000110110111011110011000010;
        end
        12947: begin
            cosine_reg0 <= 36'sb1000000000000101011101111001101011;
            sine_reg0   <= 36'sb100001000001000011011111100101001111;
        end
        12948: begin
            cosine_reg0 <= 36'sb1000000000110110001000100011001110;
            sine_reg0   <= 36'sb100001000001010000000100100011111010;
        end
        12949: begin
            cosine_reg0 <= 36'sb1000000001100110110010111000111111;
            sine_reg0   <= 36'sb100001000001011100101010101111000001;
        end
        12950: begin
            cosine_reg0 <= 36'sb1000000010010111011100111010111101;
            sine_reg0   <= 36'sb100001000001101001010010000110100011;
        end
        12951: begin
            cosine_reg0 <= 36'sb1000000011001000000110101001000101;
            sine_reg0   <= 36'sb100001000001110101111010101010100001;
        end
        12952: begin
            cosine_reg0 <= 36'sb1000000011111000110000000011010111;
            sine_reg0   <= 36'sb100001000010000010100100011010111010;
        end
        12953: begin
            cosine_reg0 <= 36'sb1000000100101001011001001001110000;
            sine_reg0   <= 36'sb100001000010001111001111010111101101;
        end
        12954: begin
            cosine_reg0 <= 36'sb1000000101011010000001111100001110;
            sine_reg0   <= 36'sb100001000010011011111011100000111001;
        end
        12955: begin
            cosine_reg0 <= 36'sb1000000110001010101010011010101111;
            sine_reg0   <= 36'sb100001000010101000101000110110011111;
        end
        12956: begin
            cosine_reg0 <= 36'sb1000000110111011010010100101010010;
            sine_reg0   <= 36'sb100001000010110101010111011000011110;
        end
        12957: begin
            cosine_reg0 <= 36'sb1000000111101011111010011011110101;
            sine_reg0   <= 36'sb100001000011000010000111000110110101;
        end
        12958: begin
            cosine_reg0 <= 36'sb1000001000011100100001111110010101;
            sine_reg0   <= 36'sb100001000011001110111000000001100100;
        end
        12959: begin
            cosine_reg0 <= 36'sb1000001001001101001001001100110001;
            sine_reg0   <= 36'sb100001000011011011101010001000101011;
        end
        12960: begin
            cosine_reg0 <= 36'sb1000001001111101110000000111000111;
            sine_reg0   <= 36'sb100001000011101000011101011100001000;
        end
        12961: begin
            cosine_reg0 <= 36'sb1000001010101110010110101101010101;
            sine_reg0   <= 36'sb100001000011110101010001111011111011;
        end
        12962: begin
            cosine_reg0 <= 36'sb1000001011011110111100111111011001;
            sine_reg0   <= 36'sb100001000100000010000111101000000101;
        end
        12963: begin
            cosine_reg0 <= 36'sb1000001100001111100010111101010010;
            sine_reg0   <= 36'sb100001000100001110111110100000100100;
        end
        12964: begin
            cosine_reg0 <= 36'sb1000001101000000001000100110111101;
            sine_reg0   <= 36'sb100001000100011011110110100101010111;
        end
        12965: begin
            cosine_reg0 <= 36'sb1000001101110000101101111100011001;
            sine_reg0   <= 36'sb100001000100101000101111110110011111;
        end
        12966: begin
            cosine_reg0 <= 36'sb1000001110100001010010111101100011;
            sine_reg0   <= 36'sb100001000100110101101010010011111011;
        end
        12967: begin
            cosine_reg0 <= 36'sb1000001111010001110111101010011011;
            sine_reg0   <= 36'sb100001000101000010100101111101101011;
        end
        12968: begin
            cosine_reg0 <= 36'sb1000010000000010011100000010111101;
            sine_reg0   <= 36'sb100001000101001111100010110011101101;
        end
        12969: begin
            cosine_reg0 <= 36'sb1000010000110011000000000111001001;
            sine_reg0   <= 36'sb100001000101011100100000110110000001;
        end
        12970: begin
            cosine_reg0 <= 36'sb1000010001100011100011110110111011;
            sine_reg0   <= 36'sb100001000101101001100000000100101000;
        end
        12971: begin
            cosine_reg0 <= 36'sb1000010010010100000111010010010100;
            sine_reg0   <= 36'sb100001000101110110100000011111100000;
        end
        12972: begin
            cosine_reg0 <= 36'sb1000010011000100101010011001001111;
            sine_reg0   <= 36'sb100001000110000011100010000110101001;
        end
        12973: begin
            cosine_reg0 <= 36'sb1000010011110101001101001011101100;
            sine_reg0   <= 36'sb100001000110010000100100111010000010;
        end
        12974: begin
            cosine_reg0 <= 36'sb1000010100100101101111101001101001;
            sine_reg0   <= 36'sb100001000110011101101000111001101011;
        end
        12975: begin
            cosine_reg0 <= 36'sb1000010101010110010001110011000100;
            sine_reg0   <= 36'sb100001000110101010101110000101100011;
        end
        12976: begin
            cosine_reg0 <= 36'sb1000010110000110110011100111111011;
            sine_reg0   <= 36'sb100001000110110111110100011101101010;
        end
        12977: begin
            cosine_reg0 <= 36'sb1000010110110111010101001000001100;
            sine_reg0   <= 36'sb100001000111000100111100000010000000;
        end
        12978: begin
            cosine_reg0 <= 36'sb1000010111100111110110010011110110;
            sine_reg0   <= 36'sb100001000111010010000100110010100011;
        end
        12979: begin
            cosine_reg0 <= 36'sb1000011000011000010111001010110101;
            sine_reg0   <= 36'sb100001000111011111001110101111010100;
        end
        12980: begin
            cosine_reg0 <= 36'sb1000011001001000110111101101001010;
            sine_reg0   <= 36'sb100001000111101100011001111000010010;
        end
        12981: begin
            cosine_reg0 <= 36'sb1000011001111001010111111010110001;
            sine_reg0   <= 36'sb100001000111111001100110001101011100;
        end
        12982: begin
            cosine_reg0 <= 36'sb1000011010101001110111110011101000;
            sine_reg0   <= 36'sb100001001000000110110011101110110010;
        end
        12983: begin
            cosine_reg0 <= 36'sb1000011011011010010111010111101111;
            sine_reg0   <= 36'sb100001001000010100000010011100010011;
        end
        12984: begin
            cosine_reg0 <= 36'sb1000011100001010110110100111000011;
            sine_reg0   <= 36'sb100001001000100001010010010101111111;
        end
        12985: begin
            cosine_reg0 <= 36'sb1000011100111011010101100001100010;
            sine_reg0   <= 36'sb100001001000101110100011011011110101;
        end
        12986: begin
            cosine_reg0 <= 36'sb1000011101101011110100000111001010;
            sine_reg0   <= 36'sb100001001000111011110101101101110101;
        end
        12987: begin
            cosine_reg0 <= 36'sb1000011110011100010010010111111001;
            sine_reg0   <= 36'sb100001001001001001001001001011111111;
        end
        12988: begin
            cosine_reg0 <= 36'sb1000011111001100110000010011101111;
            sine_reg0   <= 36'sb100001001001010110011101110110010001;
        end
        12989: begin
            cosine_reg0 <= 36'sb1000011111111101001101111010101000;
            sine_reg0   <= 36'sb100001001001100011110011101100101011;
        end
        12990: begin
            cosine_reg0 <= 36'sb1000100000101101101011001100100010;
            sine_reg0   <= 36'sb100001001001110001001010101111001101;
        end
        12991: begin
            cosine_reg0 <= 36'sb1000100001011110001000001001011101;
            sine_reg0   <= 36'sb100001001001111110100010111101110111;
        end
        12992: begin
            cosine_reg0 <= 36'sb1000100010001110100100110001010110;
            sine_reg0   <= 36'sb100001001010001011111100011000100111;
        end
        12993: begin
            cosine_reg0 <= 36'sb1000100010111111000001000100001011;
            sine_reg0   <= 36'sb100001001010011001010110111111011101;
        end
        12994: begin
            cosine_reg0 <= 36'sb1000100011101111011101000001111011;
            sine_reg0   <= 36'sb100001001010100110110010110010011001;
        end
        12995: begin
            cosine_reg0 <= 36'sb1000100100011111111000101010100011;
            sine_reg0   <= 36'sb100001001010110100001111110001011010;
        end
        12996: begin
            cosine_reg0 <= 36'sb1000100101010000010011111110000001;
            sine_reg0   <= 36'sb100001001011000001101101111100100000;
        end
        12997: begin
            cosine_reg0 <= 36'sb1000100110000000101110111100010100;
            sine_reg0   <= 36'sb100001001011001111001101010011101010;
        end
        12998: begin
            cosine_reg0 <= 36'sb1000100110110001001001100101011011;
            sine_reg0   <= 36'sb100001001011011100101101110110110111;
        end
        12999: begin
            cosine_reg0 <= 36'sb1000100111100001100011111001010010;
            sine_reg0   <= 36'sb100001001011101010001111100110001000;
        end
        13000: begin
            cosine_reg0 <= 36'sb1000101000010001111101110111111001;
            sine_reg0   <= 36'sb100001001011110111110010100001011011;
        end
        13001: begin
            cosine_reg0 <= 36'sb1000101001000010010111100001001100;
            sine_reg0   <= 36'sb100001001100000101010110101000110000;
        end
        13002: begin
            cosine_reg0 <= 36'sb1000101001110010110000110101001100;
            sine_reg0   <= 36'sb100001001100010010111011111100000110;
        end
        13003: begin
            cosine_reg0 <= 36'sb1000101010100011001001110011110100;
            sine_reg0   <= 36'sb100001001100100000100010011011011110;
        end
        13004: begin
            cosine_reg0 <= 36'sb1000101011010011100010011101000101;
            sine_reg0   <= 36'sb100001001100101110001010000110110110;
        end
        13005: begin
            cosine_reg0 <= 36'sb1000101100000011111010110000111011;
            sine_reg0   <= 36'sb100001001100111011110010111110001110;
        end
        13006: begin
            cosine_reg0 <= 36'sb1000101100110100010010101111010101;
            sine_reg0   <= 36'sb100001001101001001011101000001100101;
        end
        13007: begin
            cosine_reg0 <= 36'sb1000101101100100101010011000010010;
            sine_reg0   <= 36'sb100001001101010111001000010000111011;
        end
        13008: begin
            cosine_reg0 <= 36'sb1000101110010101000001101011101111;
            sine_reg0   <= 36'sb100001001101100100110100101100010000;
        end
        13009: begin
            cosine_reg0 <= 36'sb1000101111000101011000101001101010;
            sine_reg0   <= 36'sb100001001101110010100010010011100010;
        end
        13010: begin
            cosine_reg0 <= 36'sb1000101111110101101111010010000001;
            sine_reg0   <= 36'sb100001001110000000010001000110110010;
        end
        13011: begin
            cosine_reg0 <= 36'sb1000110000100110000101100100110011;
            sine_reg0   <= 36'sb100001001110001110000001000101111111;
        end
        13012: begin
            cosine_reg0 <= 36'sb1000110001010110011011100001111110;
            sine_reg0   <= 36'sb100001001110011011110010010001000111;
        end
        13013: begin
            cosine_reg0 <= 36'sb1000110010000110110001001001100000;
            sine_reg0   <= 36'sb100001001110101001100100101000001100;
        end
        13014: begin
            cosine_reg0 <= 36'sb1000110010110111000110011011010111;
            sine_reg0   <= 36'sb100001001110110111011000001011001100;
        end
        13015: begin
            cosine_reg0 <= 36'sb1000110011100111011011010111100001;
            sine_reg0   <= 36'sb100001001111000101001100111010000110;
        end
        13016: begin
            cosine_reg0 <= 36'sb1000110100010111101111111101111101;
            sine_reg0   <= 36'sb100001001111010011000010110100111010;
        end
        13017: begin
            cosine_reg0 <= 36'sb1000110101001000000100001110101000;
            sine_reg0   <= 36'sb100001001111100000111001111011101000;
        end
        13018: begin
            cosine_reg0 <= 36'sb1000110101111000011000001001100000;
            sine_reg0   <= 36'sb100001001111101110110010001110001111;
        end
        13019: begin
            cosine_reg0 <= 36'sb1000110110101000101011101110100101;
            sine_reg0   <= 36'sb100001001111111100101011101100101111;
        end
        13020: begin
            cosine_reg0 <= 36'sb1000110111011000111110111101110011;
            sine_reg0   <= 36'sb100001010000001010100110010111000110;
        end
        13021: begin
            cosine_reg0 <= 36'sb1000111000001001010001110111001001;
            sine_reg0   <= 36'sb100001010000011000100010001101010101;
        end
        13022: begin
            cosine_reg0 <= 36'sb1000111000111001100100011010100110;
            sine_reg0   <= 36'sb100001010000100110011111001111011011;
        end
        13023: begin
            cosine_reg0 <= 36'sb1000111001101001110110101000000110;
            sine_reg0   <= 36'sb100001010000110100011101011101010111;
        end
        13024: begin
            cosine_reg0 <= 36'sb1000111010011010001000011111101001;
            sine_reg0   <= 36'sb100001010001000010011100110111001001;
        end
        13025: begin
            cosine_reg0 <= 36'sb1000111011001010011010000001001101;
            sine_reg0   <= 36'sb100001010001010000011101011100110000;
        end
        13026: begin
            cosine_reg0 <= 36'sb1000111011111010101011001100101111;
            sine_reg0   <= 36'sb100001010001011110011111001110001101;
        end
        13027: begin
            cosine_reg0 <= 36'sb1000111100101010111100000010001111;
            sine_reg0   <= 36'sb100001010001101100100010001011011101;
        end
        13028: begin
            cosine_reg0 <= 36'sb1000111101011011001100100001101001;
            sine_reg0   <= 36'sb100001010001111010100110010100100001;
        end
        13029: begin
            cosine_reg0 <= 36'sb1000111110001011011100101010111100;
            sine_reg0   <= 36'sb100001010010001000101011101001011000;
        end
        13030: begin
            cosine_reg0 <= 36'sb1000111110111011101100011110000111;
            sine_reg0   <= 36'sb100001010010010110110010001010000001;
        end
        13031: begin
            cosine_reg0 <= 36'sb1000111111101011111011111011000111;
            sine_reg0   <= 36'sb100001010010100100111001110110011101;
        end
        13032: begin
            cosine_reg0 <= 36'sb1001000000011100001011000001111011;
            sine_reg0   <= 36'sb100001010010110011000010101110101010;
        end
        13033: begin
            cosine_reg0 <= 36'sb1001000001001100011001110010100000;
            sine_reg0   <= 36'sb100001010011000001001100110010101000;
        end
        13034: begin
            cosine_reg0 <= 36'sb1001000001111100101000001100110101;
            sine_reg0   <= 36'sb100001010011001111011000000010010111;
        end
        13035: begin
            cosine_reg0 <= 36'sb1001000010101100110110010000111000;
            sine_reg0   <= 36'sb100001010011011101100100011101110101;
        end
        13036: begin
            cosine_reg0 <= 36'sb1001000011011101000011111110100111;
            sine_reg0   <= 36'sb100001010011101011110010000101000011;
        end
        13037: begin
            cosine_reg0 <= 36'sb1001000100001101010001010110000001;
            sine_reg0   <= 36'sb100001010011111010000000110111111111;
        end
        13038: begin
            cosine_reg0 <= 36'sb1001000100111101011110010111000011;
            sine_reg0   <= 36'sb100001010100001000010000110110101001;
        end
        13039: begin
            cosine_reg0 <= 36'sb1001000101101101101011000001101011;
            sine_reg0   <= 36'sb100001010100010110100010000001000010;
        end
        13040: begin
            cosine_reg0 <= 36'sb1001000110011101110111010101111000;
            sine_reg0   <= 36'sb100001010100100100110100010111000111;
        end
        13041: begin
            cosine_reg0 <= 36'sb1001000111001110000011010011101000;
            sine_reg0   <= 36'sb100001010100110011000111111000111001;
        end
        13042: begin
            cosine_reg0 <= 36'sb1001000111111110001110111010111001;
            sine_reg0   <= 36'sb100001010101000001011100100110010111;
        end
        13043: begin
            cosine_reg0 <= 36'sb1001001000101110011010001011101001;
            sine_reg0   <= 36'sb100001010101001111110010011111100000;
        end
        13044: begin
            cosine_reg0 <= 36'sb1001001001011110100101000101110110;
            sine_reg0   <= 36'sb100001010101011110001001100100010100;
        end
        13045: begin
            cosine_reg0 <= 36'sb1001001010001110101111101001011111;
            sine_reg0   <= 36'sb100001010101101100100001110100110011;
        end
        13046: begin
            cosine_reg0 <= 36'sb1001001010111110111001110110100001;
            sine_reg0   <= 36'sb100001010101111010111011010000111011;
        end
        13047: begin
            cosine_reg0 <= 36'sb1001001011101111000011101100111011;
            sine_reg0   <= 36'sb100001010110001001010101111000101101;
        end
        13048: begin
            cosine_reg0 <= 36'sb1001001100011111001101001100101010;
            sine_reg0   <= 36'sb100001010110010111110001101100000111;
        end
        13049: begin
            cosine_reg0 <= 36'sb1001001101001111010110010101101110;
            sine_reg0   <= 36'sb100001010110100110001110101011001010;
        end
        13050: begin
            cosine_reg0 <= 36'sb1001001101111111011111001000000100;
            sine_reg0   <= 36'sb100001010110110100101100110101110100;
        end
        13051: begin
            cosine_reg0 <= 36'sb1001001110101111100111100011101010;
            sine_reg0   <= 36'sb100001010111000011001100001100000101;
        end
        13052: begin
            cosine_reg0 <= 36'sb1001001111011111101111101000011110;
            sine_reg0   <= 36'sb100001010111010001101100101101111100;
        end
        13053: begin
            cosine_reg0 <= 36'sb1001010000001111110111010110011111;
            sine_reg0   <= 36'sb100001010111100000001110011011011010;
        end
        13054: begin
            cosine_reg0 <= 36'sb1001010000111111111110101101101011;
            sine_reg0   <= 36'sb100001010111101110110001010100011100;
        end
        13055: begin
            cosine_reg0 <= 36'sb1001010001110000000101101101111111;
            sine_reg0   <= 36'sb100001010111111101010101011001000100;
        end
        13056: begin
            cosine_reg0 <= 36'sb1001010010100000001100010111011010;
            sine_reg0   <= 36'sb100001011000001011111010101001001111;
        end
        13057: begin
            cosine_reg0 <= 36'sb1001010011010000010010101001111011;
            sine_reg0   <= 36'sb100001011000011010100001000100111111;
        end
        13058: begin
            cosine_reg0 <= 36'sb1001010100000000011000100101011111;
            sine_reg0   <= 36'sb100001011000101001001000101100010001;
        end
        13059: begin
            cosine_reg0 <= 36'sb1001010100110000011110001010000100;
            sine_reg0   <= 36'sb100001011000110111110001011111000110;
        end
        13060: begin
            cosine_reg0 <= 36'sb1001010101100000100011010111101001;
            sine_reg0   <= 36'sb100001011001000110011011011101011101;
        end
        13061: begin
            cosine_reg0 <= 36'sb1001010110010000101000001110001011;
            sine_reg0   <= 36'sb100001011001010101000110100111010101;
        end
        13062: begin
            cosine_reg0 <= 36'sb1001010111000000101100101101101010;
            sine_reg0   <= 36'sb100001011001100011110010111100101110;
        end
        13063: begin
            cosine_reg0 <= 36'sb1001010111110000110000110110000010;
            sine_reg0   <= 36'sb100001011001110010100000011101101000;
        end
        13064: begin
            cosine_reg0 <= 36'sb1001011000100000110100100111010010;
            sine_reg0   <= 36'sb100001011010000001001111001010000001;
        end
        13065: begin
            cosine_reg0 <= 36'sb1001011001010000111000000001011001;
            sine_reg0   <= 36'sb100001011010001111111111000001111001;
        end
        13066: begin
            cosine_reg0 <= 36'sb1001011010000000111011000100010100;
            sine_reg0   <= 36'sb100001011010011110110000000101001111;
        end
        13067: begin
            cosine_reg0 <= 36'sb1001011010110000111101110000000010;
            sine_reg0   <= 36'sb100001011010101101100010010100000100;
        end
        13068: begin
            cosine_reg0 <= 36'sb1001011011100001000000000100100001;
            sine_reg0   <= 36'sb100001011010111100010101101110010110;
        end
        13069: begin
            cosine_reg0 <= 36'sb1001011100010001000010000001101110;
            sine_reg0   <= 36'sb100001011011001011001010010100000101;
        end
        13070: begin
            cosine_reg0 <= 36'sb1001011101000001000011100111101001;
            sine_reg0   <= 36'sb100001011011011010000000000101010000;
        end
        13071: begin
            cosine_reg0 <= 36'sb1001011101110001000100110110001110;
            sine_reg0   <= 36'sb100001011011101000110111000001110111;
        end
        13072: begin
            cosine_reg0 <= 36'sb1001011110100001000101101101011101;
            sine_reg0   <= 36'sb100001011011110111101111001001111001;
        end
        13073: begin
            cosine_reg0 <= 36'sb1001011111010001000110001101010100;
            sine_reg0   <= 36'sb100001011100000110101000011101010110;
        end
        13074: begin
            cosine_reg0 <= 36'sb1001100000000001000110010101110000;
            sine_reg0   <= 36'sb100001011100010101100010111100001101;
        end
        13075: begin
            cosine_reg0 <= 36'sb1001100000110001000110000110110000;
            sine_reg0   <= 36'sb100001011100100100011110100110011101;
        end
        13076: begin
            cosine_reg0 <= 36'sb1001100001100001000101100000010001;
            sine_reg0   <= 36'sb100001011100110011011011011100000110;
        end
        13077: begin
            cosine_reg0 <= 36'sb1001100010010001000100100010010011;
            sine_reg0   <= 36'sb100001011101000010011001011101000111;
        end
        13078: begin
            cosine_reg0 <= 36'sb1001100011000001000011001100110011;
            sine_reg0   <= 36'sb100001011101010001011000101001011111;
        end
        13079: begin
            cosine_reg0 <= 36'sb1001100011110001000001011111110000;
            sine_reg0   <= 36'sb100001011101100000011001000001001111;
        end
        13080: begin
            cosine_reg0 <= 36'sb1001100100100000111111011011000111;
            sine_reg0   <= 36'sb100001011101101111011010100100010110;
        end
        13081: begin
            cosine_reg0 <= 36'sb1001100101010000111100111110110110;
            sine_reg0   <= 36'sb100001011101111110011101010010110010;
        end
        13082: begin
            cosine_reg0 <= 36'sb1001100110000000111010001010111101;
            sine_reg0   <= 36'sb100001011110001101100001001100100100;
        end
        13083: begin
            cosine_reg0 <= 36'sb1001100110110000110110111111011000;
            sine_reg0   <= 36'sb100001011110011100100110010001101010;
        end
        13084: begin
            cosine_reg0 <= 36'sb1001100111100000110011011100000111;
            sine_reg0   <= 36'sb100001011110101011101100100010000101;
        end
        13085: begin
            cosine_reg0 <= 36'sb1001101000010000101111100001000111;
            sine_reg0   <= 36'sb100001011110111010110011111101110011;
        end
        13086: begin
            cosine_reg0 <= 36'sb1001101001000000101011001110010110;
            sine_reg0   <= 36'sb100001011111001001111100100100110100;
        end
        13087: begin
            cosine_reg0 <= 36'sb1001101001110000100110100011110011;
            sine_reg0   <= 36'sb100001011111011001000110010111001000;
        end
        13088: begin
            cosine_reg0 <= 36'sb1001101010100000100001100001011100;
            sine_reg0   <= 36'sb100001011111101000010001010100101110;
        end
        13089: begin
            cosine_reg0 <= 36'sb1001101011010000011100000111001110;
            sine_reg0   <= 36'sb100001011111110111011101011101100101;
        end
        13090: begin
            cosine_reg0 <= 36'sb1001101100000000010110010101001001;
            sine_reg0   <= 36'sb100001100000000110101010110001101100;
        end
        13091: begin
            cosine_reg0 <= 36'sb1001101100110000010000001011001010;
            sine_reg0   <= 36'sb100001100000010101111001010001000100;
        end
        13092: begin
            cosine_reg0 <= 36'sb1001101101100000001001101001001111;
            sine_reg0   <= 36'sb100001100000100101001000111011101011;
        end
        13093: begin
            cosine_reg0 <= 36'sb1001101110010000000010101111010111;
            sine_reg0   <= 36'sb100001100000110100011001110001100001;
        end
        13094: begin
            cosine_reg0 <= 36'sb1001101110111111111011011101011111;
            sine_reg0   <= 36'sb100001100001000011101011110010100110;
        end
        13095: begin
            cosine_reg0 <= 36'sb1001101111101111110011110011100110;
            sine_reg0   <= 36'sb100001100001010010111110111110111000;
        end
        13096: begin
            cosine_reg0 <= 36'sb1001110000011111101011110001101010;
            sine_reg0   <= 36'sb100001100001100010010011010110011000;
        end
        13097: begin
            cosine_reg0 <= 36'sb1001110001001111100011010111101001;
            sine_reg0   <= 36'sb100001100001110001101000111001000100;
        end
        13098: begin
            cosine_reg0 <= 36'sb1001110001111111011010100101100010;
            sine_reg0   <= 36'sb100001100010000000111111100110111100;
        end
        13099: begin
            cosine_reg0 <= 36'sb1001110010101111010001011011010010;
            sine_reg0   <= 36'sb100001100010010000010111011111111111;
        end
        13100: begin
            cosine_reg0 <= 36'sb1001110011011111000111111000110111;
            sine_reg0   <= 36'sb100001100010011111110000100100001101;
        end
        13101: begin
            cosine_reg0 <= 36'sb1001110100001110111101111110010000;
            sine_reg0   <= 36'sb100001100010101111001010110011100110;
        end
        13102: begin
            cosine_reg0 <= 36'sb1001110100111110110011101011011100;
            sine_reg0   <= 36'sb100001100010111110100110001110001000;
        end
        13103: begin
            cosine_reg0 <= 36'sb1001110101101110101001000000010111;
            sine_reg0   <= 36'sb100001100011001110000010110011110011;
        end
        13104: begin
            cosine_reg0 <= 36'sb1001110110011110011101111101000000;
            sine_reg0   <= 36'sb100001100011011101100000100100100110;
        end
        13105: begin
            cosine_reg0 <= 36'sb1001110111001110010010100001010110;
            sine_reg0   <= 36'sb100001100011101100111111100000100010;
        end
        13106: begin
            cosine_reg0 <= 36'sb1001110111111110000110101101010110;
            sine_reg0   <= 36'sb100001100011111100011111100111100100;
        end
        13107: begin
            cosine_reg0 <= 36'sb1001111000101101111010100000111111;
            sine_reg0   <= 36'sb100001100100001100000000111001101101;
        end
        13108: begin
            cosine_reg0 <= 36'sb1001111001011101101101111100001111;
            sine_reg0   <= 36'sb100001100100011011100011010110111100;
        end
        13109: begin
            cosine_reg0 <= 36'sb1001111010001101100000111111000100;
            sine_reg0   <= 36'sb100001100100101011000110111111010001;
        end
        13110: begin
            cosine_reg0 <= 36'sb1001111010111101010011101001011100;
            sine_reg0   <= 36'sb100001100100111010101011110010101011;
        end
        13111: begin
            cosine_reg0 <= 36'sb1001111011101101000101111011010101;
            sine_reg0   <= 36'sb100001100101001010010001110001001000;
        end
        13112: begin
            cosine_reg0 <= 36'sb1001111100011100110111110100101110;
            sine_reg0   <= 36'sb100001100101011001111000111010101010;
        end
        13113: begin
            cosine_reg0 <= 36'sb1001111101001100101001010101100100;
            sine_reg0   <= 36'sb100001100101101001100001001111001110;
        end
        13114: begin
            cosine_reg0 <= 36'sb1001111101111100011010011101110110;
            sine_reg0   <= 36'sb100001100101111001001010101110110101;
        end
        13115: begin
            cosine_reg0 <= 36'sb1001111110101100001011001101100010;
            sine_reg0   <= 36'sb100001100110001000110101011001011101;
        end
        13116: begin
            cosine_reg0 <= 36'sb1001111111011011111011100100100110;
            sine_reg0   <= 36'sb100001100110011000100001001111000111;
        end
        13117: begin
            cosine_reg0 <= 36'sb1010000000001011101011100011000000;
            sine_reg0   <= 36'sb100001100110101000001110001111110010;
        end
        13118: begin
            cosine_reg0 <= 36'sb1010000000111011011011001000101111;
            sine_reg0   <= 36'sb100001100110110111111100011011011100;
        end
        13119: begin
            cosine_reg0 <= 36'sb1010000001101011001010010101110001;
            sine_reg0   <= 36'sb100001100111000111101011110010000110;
        end
        13120: begin
            cosine_reg0 <= 36'sb1010000010011010111001001010000011;
            sine_reg0   <= 36'sb100001100111010111011100010011101111;
        end
        13121: begin
            cosine_reg0 <= 36'sb1010000011001010100111100101100100;
            sine_reg0   <= 36'sb100001100111100111001110000000010110;
        end
        13122: begin
            cosine_reg0 <= 36'sb1010000011111010010101101000010010;
            sine_reg0   <= 36'sb100001100111110111000000110111111010;
        end
        13123: begin
            cosine_reg0 <= 36'sb1010000100101010000011010010001011;
            sine_reg0   <= 36'sb100001101000000110110100111010011011;
        end
        13124: begin
            cosine_reg0 <= 36'sb1010000101011001110000100011001101;
            sine_reg0   <= 36'sb100001101000010110101010000111111001;
        end
        13125: begin
            cosine_reg0 <= 36'sb1010000110001001011101011011011000;
            sine_reg0   <= 36'sb100001101000100110100000100000010011;
        end
        13126: begin
            cosine_reg0 <= 36'sb1010000110111001001001111010100111;
            sine_reg0   <= 36'sb100001101000110110011000000011100111;
        end
        13127: begin
            cosine_reg0 <= 36'sb1010000111101000110110000000111011;
            sine_reg0   <= 36'sb100001101001000110010000110001110111;
        end
        13128: begin
            cosine_reg0 <= 36'sb1010001000011000100001101110010001;
            sine_reg0   <= 36'sb100001101001010110001010101011000000;
        end
        13129: begin
            cosine_reg0 <= 36'sb1010001001001000001101000010100111;
            sine_reg0   <= 36'sb100001101001100110000101101111000010;
        end
        13130: begin
            cosine_reg0 <= 36'sb1010001001110111110111111101111011;
            sine_reg0   <= 36'sb100001101001110110000001111101111101;
        end
        13131: begin
            cosine_reg0 <= 36'sb1010001010100111100010100000001100;
            sine_reg0   <= 36'sb100001101010000101111111010111110001;
        end
        13132: begin
            cosine_reg0 <= 36'sb1010001011010111001100101001010111;
            sine_reg0   <= 36'sb100001101010010101111101111100011011;
        end
        13133: begin
            cosine_reg0 <= 36'sb1010001100000110110110011001011011;
            sine_reg0   <= 36'sb100001101010100101111101101011111101;
        end
        13134: begin
            cosine_reg0 <= 36'sb1010001100110110011111110000010111;
            sine_reg0   <= 36'sb100001101010110101111110100110010101;
        end
        13135: begin
            cosine_reg0 <= 36'sb1010001101100110001000101110000111;
            sine_reg0   <= 36'sb100001101011000110000000101011100010;
        end
        13136: begin
            cosine_reg0 <= 36'sb1010001110010101110001010010101011;
            sine_reg0   <= 36'sb100001101011010110000011111011100100;
        end
        13137: begin
            cosine_reg0 <= 36'sb1010001111000101011001011110000000;
            sine_reg0   <= 36'sb100001101011100110001000010110011011;
        end
        13138: begin
            cosine_reg0 <= 36'sb1010001111110101000001010000000101;
            sine_reg0   <= 36'sb100001101011110110001101111100000110;
        end
        13139: begin
            cosine_reg0 <= 36'sb1010010000100100101000101000110111;
            sine_reg0   <= 36'sb100001101100000110010100101100100011;
        end
        13140: begin
            cosine_reg0 <= 36'sb1010010001010100001111101000010110;
            sine_reg0   <= 36'sb100001101100010110011100100111110011;
        end
        13141: begin
            cosine_reg0 <= 36'sb1010010010000011110110001110011110;
            sine_reg0   <= 36'sb100001101100100110100101101101110101;
        end
        13142: begin
            cosine_reg0 <= 36'sb1010010010110011011100011011001111;
            sine_reg0   <= 36'sb100001101100110110101111111110101001;
        end
        13143: begin
            cosine_reg0 <= 36'sb1010010011100011000010001110100111;
            sine_reg0   <= 36'sb100001101101000110111011011010001101;
        end
        13144: begin
            cosine_reg0 <= 36'sb1010010100010010100111101000100011;
            sine_reg0   <= 36'sb100001101101010111001000000000100000;
        end
        13145: begin
            cosine_reg0 <= 36'sb1010010101000010001100101001000010;
            sine_reg0   <= 36'sb100001101101100111010101110001100100;
        end
        13146: begin
            cosine_reg0 <= 36'sb1010010101110001110001010000000010;
            sine_reg0   <= 36'sb100001101101110111100100101101010110;
        end
        13147: begin
            cosine_reg0 <= 36'sb1010010110100001010101011101100001;
            sine_reg0   <= 36'sb100001101110000111110100110011110110;
        end
        13148: begin
            cosine_reg0 <= 36'sb1010010111010000111001010001011101;
            sine_reg0   <= 36'sb100001101110011000000110000101000100;
        end
        13149: begin
            cosine_reg0 <= 36'sb1010011000000000011100101011110101;
            sine_reg0   <= 36'sb100001101110101000011000100000111111;
        end
        13150: begin
            cosine_reg0 <= 36'sb1010011000101111111111101100100110;
            sine_reg0   <= 36'sb100001101110111000101100000111100110;
        end
        13151: begin
            cosine_reg0 <= 36'sb1010011001011111100010010011110000;
            sine_reg0   <= 36'sb100001101111001001000000111000111000;
        end
        13152: begin
            cosine_reg0 <= 36'sb1010011010001111000100100001001111;
            sine_reg0   <= 36'sb100001101111011001010110110100110110;
        end
        13153: begin
            cosine_reg0 <= 36'sb1010011010111110100110010101000010;
            sine_reg0   <= 36'sb100001101111101001101101111011011110;
        end
        13154: begin
            cosine_reg0 <= 36'sb1010011011101110000111101111001000;
            sine_reg0   <= 36'sb100001101111111010000110001100110000;
        end
        13155: begin
            cosine_reg0 <= 36'sb1010011100011101101000101111011110;
            sine_reg0   <= 36'sb100001110000001010011111101000101011;
        end
        13156: begin
            cosine_reg0 <= 36'sb1010011101001101001001010110000010;
            sine_reg0   <= 36'sb100001110000011010111010001111001110;
        end
        13157: begin
            cosine_reg0 <= 36'sb1010011101111100101001100010110100;
            sine_reg0   <= 36'sb100001110000101011010110000000011001;
        end
        13158: begin
            cosine_reg0 <= 36'sb1010011110101100001001010101110000;
            sine_reg0   <= 36'sb100001110000111011110010111100001100;
        end
        13159: begin
            cosine_reg0 <= 36'sb1010011111011011101000101110110110;
            sine_reg0   <= 36'sb100001110001001100010001000010100101;
        end
        13160: begin
            cosine_reg0 <= 36'sb1010100000001011000111101110000011;
            sine_reg0   <= 36'sb100001110001011100110000010011100011;
        end
        13161: begin
            cosine_reg0 <= 36'sb1010100000111010100110010011010101;
            sine_reg0   <= 36'sb100001110001101101010000101111001000;
        end
        13162: begin
            cosine_reg0 <= 36'sb1010100001101010000100011110101011;
            sine_reg0   <= 36'sb100001110001111101110010010101010001;
        end
        13163: begin
            cosine_reg0 <= 36'sb1010100010011001100010010000000011;
            sine_reg0   <= 36'sb100001110010001110010101000101111110;
        end
        13164: begin
            cosine_reg0 <= 36'sb1010100011001000111111100111011011;
            sine_reg0   <= 36'sb100001110010011110111001000001001110;
        end
        13165: begin
            cosine_reg0 <= 36'sb1010100011111000011100100100110001;
            sine_reg0   <= 36'sb100001110010101111011110000111000001;
        end
        13166: begin
            cosine_reg0 <= 36'sb1010100100100111111001001000000011;
            sine_reg0   <= 36'sb100001110011000000000100010111010110;
        end
        13167: begin
            cosine_reg0 <= 36'sb1010100101010111010101010001010000;
            sine_reg0   <= 36'sb100001110011010000101011110010001101;
        end
        13168: begin
            cosine_reg0 <= 36'sb1010100110000110110001000000010110;
            sine_reg0   <= 36'sb100001110011100001010100010111100101;
        end
        13169: begin
            cosine_reg0 <= 36'sb1010100110110110001100010101010010;
            sine_reg0   <= 36'sb100001110011110001111110000111011101;
        end
        13170: begin
            cosine_reg0 <= 36'sb1010100111100101100111010000000011;
            sine_reg0   <= 36'sb100001110100000010101001000001110100;
        end
        13171: begin
            cosine_reg0 <= 36'sb1010101000010101000001110000101000;
            sine_reg0   <= 36'sb100001110100010011010101000110101010;
        end
        13172: begin
            cosine_reg0 <= 36'sb1010101001000100011011110110111110;
            sine_reg0   <= 36'sb100001110100100100000010010101111111;
        end
        13173: begin
            cosine_reg0 <= 36'sb1010101001110011110101100011000011;
            sine_reg0   <= 36'sb100001110100110100110000101111110001;
        end
        13174: begin
            cosine_reg0 <= 36'sb1010101010100011001110110100110110;
            sine_reg0   <= 36'sb100001110101000101100000010100000000;
        end
        13175: begin
            cosine_reg0 <= 36'sb1010101011010010100111101100010101;
            sine_reg0   <= 36'sb100001110101010110010001000010101011;
        end
        13176: begin
            cosine_reg0 <= 36'sb1010101100000010000000001001011110;
            sine_reg0   <= 36'sb100001110101100111000010111011110011;
        end
        13177: begin
            cosine_reg0 <= 36'sb1010101100110001011000001100001111;
            sine_reg0   <= 36'sb100001110101110111110101111111010101;
        end
        13178: begin
            cosine_reg0 <= 36'sb1010101101100000101111110100100111;
            sine_reg0   <= 36'sb100001110110001000101010001101010010;
        end
        13179: begin
            cosine_reg0 <= 36'sb1010101110010000000111000010100011;
            sine_reg0   <= 36'sb100001110110011001011111100101101000;
        end
        13180: begin
            cosine_reg0 <= 36'sb1010101110111111011101110110000010;
            sine_reg0   <= 36'sb100001110110101010010110001000010111;
        end
        13181: begin
            cosine_reg0 <= 36'sb1010101111101110110100001111000010;
            sine_reg0   <= 36'sb100001110110111011001101110101011111;
        end
        13182: begin
            cosine_reg0 <= 36'sb1010110000011110001010001101100001;
            sine_reg0   <= 36'sb100001110111001100000110101100111111;
        end
        13183: begin
            cosine_reg0 <= 36'sb1010110001001101011111110001011101;
            sine_reg0   <= 36'sb100001110111011101000000101110110110;
        end
        13184: begin
            cosine_reg0 <= 36'sb1010110001111100110100111010110101;
            sine_reg0   <= 36'sb100001110111101101111011111011000011;
        end
        13185: begin
            cosine_reg0 <= 36'sb1010110010101100001001101001100110;
            sine_reg0   <= 36'sb100001110111111110111000010001100111;
        end
        13186: begin
            cosine_reg0 <= 36'sb1010110011011011011101111101101111;
            sine_reg0   <= 36'sb100001111000001111110101110010011111;
        end
        13187: begin
            cosine_reg0 <= 36'sb1010110100001010110001110111001110;
            sine_reg0   <= 36'sb100001111000100000110100011101101100;
        end
        13188: begin
            cosine_reg0 <= 36'sb1010110100111010000101010110000010;
            sine_reg0   <= 36'sb100001111000110001110100010011001101;
        end
        13189: begin
            cosine_reg0 <= 36'sb1010110101101001011000011010000111;
            sine_reg0   <= 36'sb100001111001000010110101010011000001;
        end
        13190: begin
            cosine_reg0 <= 36'sb1010110110011000101011000011011101;
            sine_reg0   <= 36'sb100001111001010011110111011101000111;
        end
        13191: begin
            cosine_reg0 <= 36'sb1010110111000111111101010010000010;
            sine_reg0   <= 36'sb100001111001100100111010110001100000;
        end
        13192: begin
            cosine_reg0 <= 36'sb1010110111110111001111000101110011;
            sine_reg0   <= 36'sb100001111001110101111111010000001010;
        end
        13193: begin
            cosine_reg0 <= 36'sb1010111000100110100000011110110000;
            sine_reg0   <= 36'sb100001111010000111000100111001000100;
        end
        13194: begin
            cosine_reg0 <= 36'sb1010111001010101110001011100110110;
            sine_reg0   <= 36'sb100001111010011000001011101100001111;
        end
        13195: begin
            cosine_reg0 <= 36'sb1010111010000101000010000000000011;
            sine_reg0   <= 36'sb100001111010101001010011101001101000;
        end
        13196: begin
            cosine_reg0 <= 36'sb1010111010110100010010001000010110;
            sine_reg0   <= 36'sb100001111010111010011100110001010001;
        end
        13197: begin
            cosine_reg0 <= 36'sb1010111011100011100001110101101100;
            sine_reg0   <= 36'sb100001111011001011100111000011000111;
        end
        13198: begin
            cosine_reg0 <= 36'sb1010111100010010110001001000000100;
            sine_reg0   <= 36'sb100001111011011100110010011111001010;
        end
        13199: begin
            cosine_reg0 <= 36'sb1010111101000001111111111111011101;
            sine_reg0   <= 36'sb100001111011101101111111000101011010;
        end
        13200: begin
            cosine_reg0 <= 36'sb1010111101110001001110011011110011;
            sine_reg0   <= 36'sb100001111011111111001100110101110111;
        end
        13201: begin
            cosine_reg0 <= 36'sb1010111110100000011100011101000111;
            sine_reg0   <= 36'sb100001111100010000011011110000011110;
        end
        13202: begin
            cosine_reg0 <= 36'sb1010111111001111101010000011010100;
            sine_reg0   <= 36'sb100001111100100001101011110101010000;
        end
        13203: begin
            cosine_reg0 <= 36'sb1010111111111110110111001110011011;
            sine_reg0   <= 36'sb100001111100110010111101000100001100;
        end
        13204: begin
            cosine_reg0 <= 36'sb1011000000101110000011111110011001;
            sine_reg0   <= 36'sb100001111101000100001111011101010010;
        end
        13205: begin
            cosine_reg0 <= 36'sb1011000001011101010000010011001100;
            sine_reg0   <= 36'sb100001111101010101100011000000100000;
        end
        13206: begin
            cosine_reg0 <= 36'sb1011000010001100011100001100110010;
            sine_reg0   <= 36'sb100001111101100110110111101101110110;
        end
        13207: begin
            cosine_reg0 <= 36'sb1011000010111011100111101011001001;
            sine_reg0   <= 36'sb100001111101111000001101100101010011;
        end
        13208: begin
            cosine_reg0 <= 36'sb1011000011101010110010101110010001;
            sine_reg0   <= 36'sb100001111110001001100100100110110111;
        end
        13209: begin
            cosine_reg0 <= 36'sb1011000100011001111101010110000110;
            sine_reg0   <= 36'sb100001111110011010111100110010100001;
        end
        13210: begin
            cosine_reg0 <= 36'sb1011000101001001000111100010100111;
            sine_reg0   <= 36'sb100001111110101100010110001000010000;
        end
        13211: begin
            cosine_reg0 <= 36'sb1011000101111000010001010011110011;
            sine_reg0   <= 36'sb100001111110111101110000101000000100;
        end
        13212: begin
            cosine_reg0 <= 36'sb1011000110100111011010101001100111;
            sine_reg0   <= 36'sb100001111111001111001100010001111100;
        end
        13213: begin
            cosine_reg0 <= 36'sb1011000111010110100011100100000010;
            sine_reg0   <= 36'sb100001111111100000101001000101110111;
        end
        13214: begin
            cosine_reg0 <= 36'sb1011001000000101101100000011000001;
            sine_reg0   <= 36'sb100001111111110010000111000011110101;
        end
        13215: begin
            cosine_reg0 <= 36'sb1011001000110100110100000110100100;
            sine_reg0   <= 36'sb100010000000000011100110001011110101;
        end
        13216: begin
            cosine_reg0 <= 36'sb1011001001100011111011101110101000;
            sine_reg0   <= 36'sb100010000000010101000110011101110110;
        end
        13217: begin
            cosine_reg0 <= 36'sb1011001010010011000010111011001011;
            sine_reg0   <= 36'sb100010000000100110100111111001110111;
        end
        13218: begin
            cosine_reg0 <= 36'sb1011001011000010001001101100001011;
            sine_reg0   <= 36'sb100010000000111000001010011111111001;
        end
        13219: begin
            cosine_reg0 <= 36'sb1011001011110001010000000001100111;
            sine_reg0   <= 36'sb100010000001001001101110001111111001;
        end
        13220: begin
            cosine_reg0 <= 36'sb1011001100100000010101111011011110;
            sine_reg0   <= 36'sb100010000001011011010011001001111001;
        end
        13221: begin
            cosine_reg0 <= 36'sb1011001101001111011011011001101100;
            sine_reg0   <= 36'sb100010000001101100111001001101110110;
        end
        13222: begin
            cosine_reg0 <= 36'sb1011001101111110100000011100010001;
            sine_reg0   <= 36'sb100010000001111110100000011011110000;
        end
        13223: begin
            cosine_reg0 <= 36'sb1011001110101101100101000011001010;
            sine_reg0   <= 36'sb100010000010010000001000110011100111;
        end
        13224: begin
            cosine_reg0 <= 36'sb1011001111011100101001001110010101;
            sine_reg0   <= 36'sb100010000010100001110010010101011010;
        end
        13225: begin
            cosine_reg0 <= 36'sb1011010000001011101100111101110010;
            sine_reg0   <= 36'sb100010000010110011011101000001001000;
        end
        13226: begin
            cosine_reg0 <= 36'sb1011010000111010110000010001011101;
            sine_reg0   <= 36'sb100010000011000101001000110110110000;
        end
        13227: begin
            cosine_reg0 <= 36'sb1011010001101001110011001001010110;
            sine_reg0   <= 36'sb100010000011010110110101110110010011;
        end
        13228: begin
            cosine_reg0 <= 36'sb1011010010011000110101100101011010;
            sine_reg0   <= 36'sb100010000011101000100011111111101110;
        end
        13229: begin
            cosine_reg0 <= 36'sb1011010011000111110111100101101000;
            sine_reg0   <= 36'sb100010000011111010010011010011000010;
        end
        13230: begin
            cosine_reg0 <= 36'sb1011010011110110111001001001111110;
            sine_reg0   <= 36'sb100010000100001100000011110000001110;
        end
        13231: begin
            cosine_reg0 <= 36'sb1011010100100101111010010010011001;
            sine_reg0   <= 36'sb100010000100011101110101010111010000;
        end
        13232: begin
            cosine_reg0 <= 36'sb1011010101010100111010111110111001;
            sine_reg0   <= 36'sb100010000100101111101000001000001001;
        end
        13233: begin
            cosine_reg0 <= 36'sb1011010110000011111011001111011010;
            sine_reg0   <= 36'sb100010000101000001011100000010111000;
        end
        13234: begin
            cosine_reg0 <= 36'sb1011010110110010111011000011111101;
            sine_reg0   <= 36'sb100010000101010011010001000111011100;
        end
        13235: begin
            cosine_reg0 <= 36'sb1011010111100001111010011100011110;
            sine_reg0   <= 36'sb100010000101100101000111010101110100;
        end
        13236: begin
            cosine_reg0 <= 36'sb1011011000010000111001011000111100;
            sine_reg0   <= 36'sb100010000101110110111110101110000000;
        end
        13237: begin
            cosine_reg0 <= 36'sb1011011000111111110111111001010101;
            sine_reg0   <= 36'sb100010000110001000110111001111111111;
        end
        13238: begin
            cosine_reg0 <= 36'sb1011011001101110110101111101101000;
            sine_reg0   <= 36'sb100010000110011010110000111011110000;
        end
        13239: begin
            cosine_reg0 <= 36'sb1011011010011101110011100101110001;
            sine_reg0   <= 36'sb100010000110101100101011110001010010;
        end
        13240: begin
            cosine_reg0 <= 36'sb1011011011001100110000110001110001;
            sine_reg0   <= 36'sb100010000110111110100111110000100110;
        end
        13241: begin
            cosine_reg0 <= 36'sb1011011011111011101101100001100100;
            sine_reg0   <= 36'sb100010000111010000100100111001101001;
        end
        13242: begin
            cosine_reg0 <= 36'sb1011011100101010101001110101001010;
            sine_reg0   <= 36'sb100010000111100010100011001100011100;
        end
        13243: begin
            cosine_reg0 <= 36'sb1011011101011001100101101100011111;
            sine_reg0   <= 36'sb100010000111110100100010101000111110;
        end
        13244: begin
            cosine_reg0 <= 36'sb1011011110001000100001000111100011;
            sine_reg0   <= 36'sb100010001000000110100011001111001110;
        end
        13245: begin
            cosine_reg0 <= 36'sb1011011110110111011100000110010100;
            sine_reg0   <= 36'sb100010001000011000100100111111001100;
        end
        13246: begin
            cosine_reg0 <= 36'sb1011011111100110010110101000101111;
            sine_reg0   <= 36'sb100010001000101010100111111000110110;
        end
        13247: begin
            cosine_reg0 <= 36'sb1011100000010101010000101110110011;
            sine_reg0   <= 36'sb100010001000111100101011111100001100;
        end
        13248: begin
            cosine_reg0 <= 36'sb1011100001000100001010011000011111;
            sine_reg0   <= 36'sb100010001001001110110001001001001110;
        end
        13249: begin
            cosine_reg0 <= 36'sb1011100001110011000011100101110000;
            sine_reg0   <= 36'sb100010001001100000110111011111111010;
        end
        13250: begin
            cosine_reg0 <= 36'sb1011100010100001111100010110100100;
            sine_reg0   <= 36'sb100010001001110010111111000000010000;
        end
        13251: begin
            cosine_reg0 <= 36'sb1011100011010000110100101010111010;
            sine_reg0   <= 36'sb100010001010000101000111101010001111;
        end
        13252: begin
            cosine_reg0 <= 36'sb1011100011111111101100100010110001;
            sine_reg0   <= 36'sb100010001010010111010001011101110111;
        end
        13253: begin
            cosine_reg0 <= 36'sb1011100100101110100011111110000101;
            sine_reg0   <= 36'sb100010001010101001011100011011000111;
        end
        13254: begin
            cosine_reg0 <= 36'sb1011100101011101011010111100110101;
            sine_reg0   <= 36'sb100010001010111011101000100001111110;
        end
        13255: begin
            cosine_reg0 <= 36'sb1011100110001100010001011111000001;
            sine_reg0   <= 36'sb100010001011001101110101110010011011;
        end
        13256: begin
            cosine_reg0 <= 36'sb1011100110111011000111100100100100;
            sine_reg0   <= 36'sb100010001011100000000100001100011110;
        end
        13257: begin
            cosine_reg0 <= 36'sb1011100111101001111101001101011111;
            sine_reg0   <= 36'sb100010001011110010010011110000000110;
        end
        13258: begin
            cosine_reg0 <= 36'sb1011101000011000110010011001101111;
            sine_reg0   <= 36'sb100010001100000100100100011101010011;
        end
        13259: begin
            cosine_reg0 <= 36'sb1011101001000111100111001001010010;
            sine_reg0   <= 36'sb100010001100010110110110010100000011;
        end
        13260: begin
            cosine_reg0 <= 36'sb1011101001110110011011011100000111;
            sine_reg0   <= 36'sb100010001100101001001001010100010110;
        end
        13261: begin
            cosine_reg0 <= 36'sb1011101010100101001111010010001011;
            sine_reg0   <= 36'sb100010001100111011011101011110001011;
        end
        13262: begin
            cosine_reg0 <= 36'sb1011101011010100000010101011011101;
            sine_reg0   <= 36'sb100010001101001101110010110001100010;
        end
        13263: begin
            cosine_reg0 <= 36'sb1011101100000010110101100111111100;
            sine_reg0   <= 36'sb100010001101100000001001001110011001;
        end
        13264: begin
            cosine_reg0 <= 36'sb1011101100110001101000000111100100;
            sine_reg0   <= 36'sb100010001101110010100000110100110001;
        end
        13265: begin
            cosine_reg0 <= 36'sb1011101101100000011010001010010101;
            sine_reg0   <= 36'sb100010001110000100111001100100101000;
        end
        13266: begin
            cosine_reg0 <= 36'sb1011101110001111001011110000001101;
            sine_reg0   <= 36'sb100010001110010111010011011101111101;
        end
        13267: begin
            cosine_reg0 <= 36'sb1011101110111101111100111001001001;
            sine_reg0   <= 36'sb100010001110101001101110100000110001;
        end
        13268: begin
            cosine_reg0 <= 36'sb1011101111101100101101100101001001;
            sine_reg0   <= 36'sb100010001110111100001010101101000010;
        end
        13269: begin
            cosine_reg0 <= 36'sb1011110000011011011101110100001010;
            sine_reg0   <= 36'sb100010001111001110101000000010101111;
        end
        13270: begin
            cosine_reg0 <= 36'sb1011110001001010001101100110001010;
            sine_reg0   <= 36'sb100010001111100001000110100001111000;
        end
        13271: begin
            cosine_reg0 <= 36'sb1011110001111000111100111011001000;
            sine_reg0   <= 36'sb100010001111110011100110001010011101;
        end
        13272: begin
            cosine_reg0 <= 36'sb1011110010100111101011110011000010;
            sine_reg0   <= 36'sb100010010000000110000110111100011100;
        end
        13273: begin
            cosine_reg0 <= 36'sb1011110011010110011010001101110110;
            sine_reg0   <= 36'sb100010010000011000101000110111110100;
        end
        13274: begin
            cosine_reg0 <= 36'sb1011110100000101001000001011100010;
            sine_reg0   <= 36'sb100010010000101011001011111100100101;
        end
        13275: begin
            cosine_reg0 <= 36'sb1011110100110011110101101100000101;
            sine_reg0   <= 36'sb100010010000111101110000001010101111;
        end
        13276: begin
            cosine_reg0 <= 36'sb1011110101100010100010101111011100;
            sine_reg0   <= 36'sb100010010001010000010101100010010000;
        end
        13277: begin
            cosine_reg0 <= 36'sb1011110110010001001111010101100110;
            sine_reg0   <= 36'sb100010010001100010111100000011001001;
        end
        13278: begin
            cosine_reg0 <= 36'sb1011110110111111111011011110100001;
            sine_reg0   <= 36'sb100010010001110101100011101101010111;
        end
        13279: begin
            cosine_reg0 <= 36'sb1011110111101110100111001010001100;
            sine_reg0   <= 36'sb100010010010001000001100100000111010;
        end
        13280: begin
            cosine_reg0 <= 36'sb1011111000011101010010011000100011;
            sine_reg0   <= 36'sb100010010010011010110110011101110011;
        end
        13281: begin
            cosine_reg0 <= 36'sb1011111001001011111101001001100111;
            sine_reg0   <= 36'sb100010010010101101100001100011111111;
        end
        13282: begin
            cosine_reg0 <= 36'sb1011111001111010100111011101010100;
            sine_reg0   <= 36'sb100010010011000000001101110011011111;
        end
        13283: begin
            cosine_reg0 <= 36'sb1011111010101001010001010011101001;
            sine_reg0   <= 36'sb100010010011010010111011001100010001;
        end
        13284: begin
            cosine_reg0 <= 36'sb1011111011010111111010101100100101;
            sine_reg0   <= 36'sb100010010011100101101001101110010100;
        end
        13285: begin
            cosine_reg0 <= 36'sb1011111100000110100011101000000101;
            sine_reg0   <= 36'sb100010010011111000011001011001101001;
        end
        13286: begin
            cosine_reg0 <= 36'sb1011111100110101001100000110001000;
            sine_reg0   <= 36'sb100010010100001011001010001110001111;
        end
        13287: begin
            cosine_reg0 <= 36'sb1011111101100011110100000110101011;
            sine_reg0   <= 36'sb100010010100011101111100001100000011;
        end
        13288: begin
            cosine_reg0 <= 36'sb1011111110010010011011101001101110;
            sine_reg0   <= 36'sb100010010100110000101111010011000111;
        end
        13289: begin
            cosine_reg0 <= 36'sb1011111111000001000010101111001110;
            sine_reg0   <= 36'sb100010010101000011100011100011011001;
        end
        13290: begin
            cosine_reg0 <= 36'sb1011111111101111101001010111001001;
            sine_reg0   <= 36'sb100010010101010110011000111100111001;
        end
        13291: begin
            cosine_reg0 <= 36'sb1100000000011110001111100001011110;
            sine_reg0   <= 36'sb100010010101101001001111011111100101;
        end
        13292: begin
            cosine_reg0 <= 36'sb1100000001001100110101001110001011;
            sine_reg0   <= 36'sb100010010101111100000111001011011101;
        end
        13293: begin
            cosine_reg0 <= 36'sb1100000001111011011010011101001110;
            sine_reg0   <= 36'sb100010010110001111000000000000100001;
        end
        13294: begin
            cosine_reg0 <= 36'sb1100000010101001111111001110100101;
            sine_reg0   <= 36'sb100010010110100001111001111110101111;
        end
        13295: begin
            cosine_reg0 <= 36'sb1100000011011000100011100010001111;
            sine_reg0   <= 36'sb100010010110110100110101000110000110;
        end
        13296: begin
            cosine_reg0 <= 36'sb1100000100000111000111011000001001;
            sine_reg0   <= 36'sb100010010111000111110001010110100111;
        end
        13297: begin
            cosine_reg0 <= 36'sb1100000100110101101010110000010011;
            sine_reg0   <= 36'sb100010010111011010101110110000010001;
        end
        13298: begin
            cosine_reg0 <= 36'sb1100000101100100001101101010101001;
            sine_reg0   <= 36'sb100010010111101101101101010011000001;
        end
        13299: begin
            cosine_reg0 <= 36'sb1100000110010010110000000111001011;
            sine_reg0   <= 36'sb100010011000000000101100111110111001;
        end
        13300: begin
            cosine_reg0 <= 36'sb1100000111000001010010000101110110;
            sine_reg0   <= 36'sb100010011000010011101101110011110111;
        end
        13301: begin
            cosine_reg0 <= 36'sb1100000111101111110011100110101001;
            sine_reg0   <= 36'sb100010011000100110101111110001111011;
        end
        13302: begin
            cosine_reg0 <= 36'sb1100001000011110010100101001100010;
            sine_reg0   <= 36'sb100010011000111001110010111001000011;
        end
        13303: begin
            cosine_reg0 <= 36'sb1100001001001100110101001110011111;
            sine_reg0   <= 36'sb100010011001001100110111001001001111;
        end
        13304: begin
            cosine_reg0 <= 36'sb1100001001111011010101010101011110;
            sine_reg0   <= 36'sb100010011001011111111100100010011110;
        end
        13305: begin
            cosine_reg0 <= 36'sb1100001010101001110100111110011110;
            sine_reg0   <= 36'sb100010011001110011000011000100110000;
        end
        13306: begin
            cosine_reg0 <= 36'sb1100001011011000010100001001011101;
            sine_reg0   <= 36'sb100010011010000110001010110000000011;
        end
        13307: begin
            cosine_reg0 <= 36'sb1100001100000110110010110110011000;
            sine_reg0   <= 36'sb100010011010011001010011100100011000;
        end
        13308: begin
            cosine_reg0 <= 36'sb1100001100110101010001000101001111;
            sine_reg0   <= 36'sb100010011010101100011101100001101101;
        end
        13309: begin
            cosine_reg0 <= 36'sb1100001101100011101110110101111111;
            sine_reg0   <= 36'sb100010011010111111101000101000000001;
        end
        13310: begin
            cosine_reg0 <= 36'sb1100001110010010001100001000100111;
            sine_reg0   <= 36'sb100010011011010010110100110111010100;
        end
        13311: begin
            cosine_reg0 <= 36'sb1100001111000000101000111101000100;
            sine_reg0   <= 36'sb100010011011100110000010001111100110;
        end
        13312: begin
            cosine_reg0 <= 36'sb1100001111101111000101010011010101;
            sine_reg0   <= 36'sb100010011011111001010000110000110100;
        end
        13313: begin
            cosine_reg0 <= 36'sb1100010000011101100001001011011001;
            sine_reg0   <= 36'sb100010011100001100100000011010111111;
        end
        13314: begin
            cosine_reg0 <= 36'sb1100010001001011111100100101001101;
            sine_reg0   <= 36'sb100010011100011111110001001110000110;
        end
        13315: begin
            cosine_reg0 <= 36'sb1100010001111010010111100000110000;
            sine_reg0   <= 36'sb100010011100110011000011001010001001;
        end
        13316: begin
            cosine_reg0 <= 36'sb1100010010101000110001111101111111;
            sine_reg0   <= 36'sb100010011101000110010110001111000101;
        end
        13317: begin
            cosine_reg0 <= 36'sb1100010011010111001011111100111010;
            sine_reg0   <= 36'sb100010011101011001101010011100111011;
        end
        13318: begin
            cosine_reg0 <= 36'sb1100010100000101100101011101011110;
            sine_reg0   <= 36'sb100010011101101100111111110011101010;
        end
        13319: begin
            cosine_reg0 <= 36'sb1100010100110011111110011111101001;
            sine_reg0   <= 36'sb100010011110000000010110010011010001;
        end
        13320: begin
            cosine_reg0 <= 36'sb1100010101100010010111000011011010;
            sine_reg0   <= 36'sb100010011110010011101101111011110000;
        end
        13321: begin
            cosine_reg0 <= 36'sb1100010110010000101111001000101111;
            sine_reg0   <= 36'sb100010011110100111000110101101000101;
        end
        13322: begin
            cosine_reg0 <= 36'sb1100010110111111000110101111100110;
            sine_reg0   <= 36'sb100010011110111010100000100111010000;
        end
        13323: begin
            cosine_reg0 <= 36'sb1100010111101101011101110111111110;
            sine_reg0   <= 36'sb100010011111001101111011101010010000;
        end
        13324: begin
            cosine_reg0 <= 36'sb1100011000011011110100100001110100;
            sine_reg0   <= 36'sb100010011111100001010111110110000100;
        end
        13325: begin
            cosine_reg0 <= 36'sb1100011001001010001010101101000110;
            sine_reg0   <= 36'sb100010011111110100110101001010101100;
        end
        13326: begin
            cosine_reg0 <= 36'sb1100011001111000100000011001110100;
            sine_reg0   <= 36'sb100010100000001000010011101000000111;
        end
        13327: begin
            cosine_reg0 <= 36'sb1100011010100110110101100111111011;
            sine_reg0   <= 36'sb100010100000011011110011001110010100;
        end
        13328: begin
            cosine_reg0 <= 36'sb1100011011010101001010010111011001;
            sine_reg0   <= 36'sb100010100000101111010011111101010011;
        end
        13329: begin
            cosine_reg0 <= 36'sb1100011100000011011110101000001100;
            sine_reg0   <= 36'sb100010100001000010110101110101000010;
        end
        13330: begin
            cosine_reg0 <= 36'sb1100011100110001110010011010010100;
            sine_reg0   <= 36'sb100010100001010110011000110101100001;
        end
        13331: begin
            cosine_reg0 <= 36'sb1100011101100000000101101101101110;
            sine_reg0   <= 36'sb100010100001101001111100111110101111;
        end
        13332: begin
            cosine_reg0 <= 36'sb1100011110001110011000100010010111;
            sine_reg0   <= 36'sb100010100001111101100010010000101011;
        end
        13333: begin
            cosine_reg0 <= 36'sb1100011110111100101010111000010000;
            sine_reg0   <= 36'sb100010100010010001001000101011010101;
        end
        13334: begin
            cosine_reg0 <= 36'sb1100011111101010111100101111010101;
            sine_reg0   <= 36'sb100010100010100100110000001110101100;
        end
        13335: begin
            cosine_reg0 <= 36'sb1100100000011001001110000111100101;
            sine_reg0   <= 36'sb100010100010111000011000111010110000;
        end
        13336: begin
            cosine_reg0 <= 36'sb1100100001000111011111000000111110;
            sine_reg0   <= 36'sb100010100011001100000010101111011110;
        end
        13337: begin
            cosine_reg0 <= 36'sb1100100001110101101111011011011110;
            sine_reg0   <= 36'sb100010100011011111101101101100110111;
        end
        13338: begin
            cosine_reg0 <= 36'sb1100100010100011111111010111000100;
            sine_reg0   <= 36'sb100010100011110011011001110010111010;
        end
        13339: begin
            cosine_reg0 <= 36'sb1100100011010010001110110011101101;
            sine_reg0   <= 36'sb100010100100000111000111000001100110;
        end
        13340: begin
            cosine_reg0 <= 36'sb1100100100000000011101110001011001;
            sine_reg0   <= 36'sb100010100100011010110101011000111010;
        end
        13341: begin
            cosine_reg0 <= 36'sb1100100100101110101100010000000101;
            sine_reg0   <= 36'sb100010100100101110100100111000110110;
        end
        13342: begin
            cosine_reg0 <= 36'sb1100100101011100111010001111101111;
            sine_reg0   <= 36'sb100010100101000010010101100001011000;
        end
        13343: begin
            cosine_reg0 <= 36'sb1100100110001011000111110000010110;
            sine_reg0   <= 36'sb100010100101010110000111010010100001;
        end
        13344: begin
            cosine_reg0 <= 36'sb1100100110111001010100110001110111;
            sine_reg0   <= 36'sb100010100101101001111010001100001110;
        end
        13345: begin
            cosine_reg0 <= 36'sb1100100111100111100001010100010010;
            sine_reg0   <= 36'sb100010100101111101101110001110100001;
        end
        13346: begin
            cosine_reg0 <= 36'sb1100101000010101101101010111100100;
            sine_reg0   <= 36'sb100010100110010001100011011001010111;
        end
        13347: begin
            cosine_reg0 <= 36'sb1100101001000011111000111011101011;
            sine_reg0   <= 36'sb100010100110100101011001101100110000;
        end
        13348: begin
            cosine_reg0 <= 36'sb1100101001110010000100000000100111;
            sine_reg0   <= 36'sb100010100110111001010001001000101011;
        end
        13349: begin
            cosine_reg0 <= 36'sb1100101010100000001110100110010100;
            sine_reg0   <= 36'sb100010100111001101001001101101001000;
        end
        13350: begin
            cosine_reg0 <= 36'sb1100101011001110011000101100110001;
            sine_reg0   <= 36'sb100010100111100001000011011010000101;
        end
        13351: begin
            cosine_reg0 <= 36'sb1100101011111100100010010011111101;
            sine_reg0   <= 36'sb100010100111110100111110001111100010;
        end
        13352: begin
            cosine_reg0 <= 36'sb1100101100101010101011011011110101;
            sine_reg0   <= 36'sb100010101000001000111010001101011111;
        end
        13353: begin
            cosine_reg0 <= 36'sb1100101101011000110100000100011000;
            sine_reg0   <= 36'sb100010101000011100110111010011111010;
        end
        13354: begin
            cosine_reg0 <= 36'sb1100101110000110111100001101100100;
            sine_reg0   <= 36'sb100010101000110000110101100010110010;
        end
        13355: begin
            cosine_reg0 <= 36'sb1100101110110101000011110111011000;
            sine_reg0   <= 36'sb100010101001000100110100111010000111;
        end
        13356: begin
            cosine_reg0 <= 36'sb1100101111100011001011000001110001;
            sine_reg0   <= 36'sb100010101001011000110101011001111000;
        end
        13357: begin
            cosine_reg0 <= 36'sb1100110000010001010001101100101101;
            sine_reg0   <= 36'sb100010101001101100110111000010000101;
        end
        13358: begin
            cosine_reg0 <= 36'sb1100110000111111010111111000001100;
            sine_reg0   <= 36'sb100010101010000000111001110010101100;
        end
        13359: begin
            cosine_reg0 <= 36'sb1100110001101101011101100100001011;
            sine_reg0   <= 36'sb100010101010010100111101101011101101;
        end
        13360: begin
            cosine_reg0 <= 36'sb1100110010011011100010110000101000;
            sine_reg0   <= 36'sb100010101010101001000010101101000111;
        end
        13361: begin
            cosine_reg0 <= 36'sb1100110011001001100111011101100010;
            sine_reg0   <= 36'sb100010101010111101001000110110111001;
        end
        13362: begin
            cosine_reg0 <= 36'sb1100110011110111101011101010110110;
            sine_reg0   <= 36'sb100010101011010001010000001001000010;
        end
        13363: begin
            cosine_reg0 <= 36'sb1100110100100101101111011000100100;
            sine_reg0   <= 36'sb100010101011100101011000100011100010;
        end
        13364: begin
            cosine_reg0 <= 36'sb1100110101010011110010100110101001;
            sine_reg0   <= 36'sb100010101011111001100010000110011000;
        end
        13365: begin
            cosine_reg0 <= 36'sb1100110110000001110101010101000011;
            sine_reg0   <= 36'sb100010101100001101101100110001100011;
        end
        13366: begin
            cosine_reg0 <= 36'sb1100110110101111110111100011110001;
            sine_reg0   <= 36'sb100010101100100001111000100101000010;
        end
        13367: begin
            cosine_reg0 <= 36'sb1100110111011101111001010010110001;
            sine_reg0   <= 36'sb100010101100110110000101100000110101;
        end
        13368: begin
            cosine_reg0 <= 36'sb1100111000001011111010100010000001;
            sine_reg0   <= 36'sb100010101101001010010011100100111011;
        end
        13369: begin
            cosine_reg0 <= 36'sb1100111000111001111011010001100000;
            sine_reg0   <= 36'sb100010101101011110100010110001010010;
        end
        13370: begin
            cosine_reg0 <= 36'sb1100111001100111111011100001001011;
            sine_reg0   <= 36'sb100010101101110010110011000101111011;
        end
        13371: begin
            cosine_reg0 <= 36'sb1100111010010101111011010001000001;
            sine_reg0   <= 36'sb100010101110000111000100100010110100;
        end
        13372: begin
            cosine_reg0 <= 36'sb1100111011000011111010100001000001;
            sine_reg0   <= 36'sb100010101110011011010111000111111101;
        end
        13373: begin
            cosine_reg0 <= 36'sb1100111011110001111001010001000111;
            sine_reg0   <= 36'sb100010101110101111101010110101010101;
        end
        13374: begin
            cosine_reg0 <= 36'sb1100111100011111110111100001010011;
            sine_reg0   <= 36'sb100010101111000011111111101010111011;
        end
        13375: begin
            cosine_reg0 <= 36'sb1100111101001101110101010001100011;
            sine_reg0   <= 36'sb100010101111011000010101101000101110;
        end
        13376: begin
            cosine_reg0 <= 36'sb1100111101111011110010100001110101;
            sine_reg0   <= 36'sb100010101111101100101100101110101101;
        end
        13377: begin
            cosine_reg0 <= 36'sb1100111110101001101111010010000111;
            sine_reg0   <= 36'sb100010110000000001000100111100111001;
        end
        13378: begin
            cosine_reg0 <= 36'sb1100111111010111101011100010010111;
            sine_reg0   <= 36'sb100010110000010101011110010011001111;
        end
        13379: begin
            cosine_reg0 <= 36'sb1101000000000101100111010010100100;
            sine_reg0   <= 36'sb100010110000101001111000110001101111;
        end
        13380: begin
            cosine_reg0 <= 36'sb1101000000110011100010100010101100;
            sine_reg0   <= 36'sb100010110000111110010100011000011001;
        end
        13381: begin
            cosine_reg0 <= 36'sb1101000001100001011101010010101110;
            sine_reg0   <= 36'sb100010110001010010110001000111001011;
        end
        13382: begin
            cosine_reg0 <= 36'sb1101000010001111010111100010100110;
            sine_reg0   <= 36'sb100010110001100111001110111110000110;
        end
        13383: begin
            cosine_reg0 <= 36'sb1101000010111101010001010010010100;
            sine_reg0   <= 36'sb100010110001111011101101111101000111;
        end
        13384: begin
            cosine_reg0 <= 36'sb1101000011101011001010100001110110;
            sine_reg0   <= 36'sb100010110010010000001110000100001110;
        end
        13385: begin
            cosine_reg0 <= 36'sb1101000100011001000011010001001010;
            sine_reg0   <= 36'sb100010110010100100101111010011011011;
        end
        13386: begin
            cosine_reg0 <= 36'sb1101000101000110111011100000001111;
            sine_reg0   <= 36'sb100010110010111001010001101010101100;
        end
        13387: begin
            cosine_reg0 <= 36'sb1101000101110100110011001111000001;
            sine_reg0   <= 36'sb100010110011001101110101001010000001;
        end
        13388: begin
            cosine_reg0 <= 36'sb1101000110100010101010011101100001;
            sine_reg0   <= 36'sb100010110011100010011001110001011001;
        end
        13389: begin
            cosine_reg0 <= 36'sb1101000111010000100001001011101100;
            sine_reg0   <= 36'sb100010110011110110111111100000110100;
        end
        13390: begin
            cosine_reg0 <= 36'sb1101000111111110010111011001011111;
            sine_reg0   <= 36'sb100010110100001011100110011000010000;
        end
        13391: begin
            cosine_reg0 <= 36'sb1101001000101100001101000110111011;
            sine_reg0   <= 36'sb100010110100100000001110010111101100;
        end
        13392: begin
            cosine_reg0 <= 36'sb1101001001011010000010010011111011;
            sine_reg0   <= 36'sb100010110100110100110111011111001001;
        end
        13393: begin
            cosine_reg0 <= 36'sb1101001010000111110111000000100000;
            sine_reg0   <= 36'sb100010110101001001100001101110100100;
        end
        13394: begin
            cosine_reg0 <= 36'sb1101001010110101101011001100100111;
            sine_reg0   <= 36'sb100010110101011110001101000101111110;
        end
        13395: begin
            cosine_reg0 <= 36'sb1101001011100011011110111000001111;
            sine_reg0   <= 36'sb100010110101110010111001100101010101;
        end
        13396: begin
            cosine_reg0 <= 36'sb1101001100010001010010000011010100;
            sine_reg0   <= 36'sb100010110110000111100111001100101001;
        end
        13397: begin
            cosine_reg0 <= 36'sb1101001100111111000100101101110111;
            sine_reg0   <= 36'sb100010110110011100010101111011111001;
        end
        13398: begin
            cosine_reg0 <= 36'sb1101001101101100110110110111110101;
            sine_reg0   <= 36'sb100010110110110001000101110011000100;
        end
        13399: begin
            cosine_reg0 <= 36'sb1101001110011010101000100001001100;
            sine_reg0   <= 36'sb100010110111000101110110110010001001;
        end
        13400: begin
            cosine_reg0 <= 36'sb1101001111001000011001101001111011;
            sine_reg0   <= 36'sb100010110111011010101000111001000111;
        end
        13401: begin
            cosine_reg0 <= 36'sb1101001111110110001010010010000000;
            sine_reg0   <= 36'sb100010110111101111011100000111111111;
        end
        13402: begin
            cosine_reg0 <= 36'sb1101010000100011111010011001011000;
            sine_reg0   <= 36'sb100010111000000100010000011110101110;
        end
        13403: begin
            cosine_reg0 <= 36'sb1101010001010001101010000000000011;
            sine_reg0   <= 36'sb100010111000011001000101111101010100;
        end
        13404: begin
            cosine_reg0 <= 36'sb1101010001111111011001000101111110;
            sine_reg0   <= 36'sb100010111000101101111100100011110001;
        end
        13405: begin
            cosine_reg0 <= 36'sb1101010010101101000111101011001000;
            sine_reg0   <= 36'sb100010111001000010110100010010000011;
        end
        13406: begin
            cosine_reg0 <= 36'sb1101010011011010110101101111011111;
            sine_reg0   <= 36'sb100010111001010111101101001000001001;
        end
        13407: begin
            cosine_reg0 <= 36'sb1101010100001000100011010011000010;
            sine_reg0   <= 36'sb100010111001101100100111000110000100;
        end
        13408: begin
            cosine_reg0 <= 36'sb1101010100110110010000010101101101;
            sine_reg0   <= 36'sb100010111010000001100010001011110001;
        end
        13409: begin
            cosine_reg0 <= 36'sb1101010101100011111100110111100001;
            sine_reg0   <= 36'sb100010111010010110011110011001010001;
        end
        13410: begin
            cosine_reg0 <= 36'sb1101010110010001101000111000011010;
            sine_reg0   <= 36'sb100010111010101011011011101110100010;
        end
        13411: begin
            cosine_reg0 <= 36'sb1101010110111111010100011000010111;
            sine_reg0   <= 36'sb100010111011000000011010001011100100;
        end
        13412: begin
            cosine_reg0 <= 36'sb1101010111101100111111010111010111;
            sine_reg0   <= 36'sb100010111011010101011001110000010110;
        end
        13413: begin
            cosine_reg0 <= 36'sb1101011000011010101001110101011000;
            sine_reg0   <= 36'sb100010111011101010011010011100110111;
        end
        13414: begin
            cosine_reg0 <= 36'sb1101011001001000010011110010010111;
            sine_reg0   <= 36'sb100010111011111111011100010001000101;
        end
        13415: begin
            cosine_reg0 <= 36'sb1101011001110101111101001110010011;
            sine_reg0   <= 36'sb100010111100010100011111001101000010;
        end
        13416: begin
            cosine_reg0 <= 36'sb1101011010100011100110001001001011;
            sine_reg0   <= 36'sb100010111100101001100011010000101010;
        end
        13417: begin
            cosine_reg0 <= 36'sb1101011011010001001110100010111101;
            sine_reg0   <= 36'sb100010111100111110101000011011111111;
        end
        13418: begin
            cosine_reg0 <= 36'sb1101011011111110110110011011100110;
            sine_reg0   <= 36'sb100010111101010011101110101110111111;
        end
        13419: begin
            cosine_reg0 <= 36'sb1101011100101100011101110011000101;
            sine_reg0   <= 36'sb100010111101101000110110001001101000;
        end
        13420: begin
            cosine_reg0 <= 36'sb1101011101011010000100101001011001;
            sine_reg0   <= 36'sb100010111101111101111110101011111011;
        end
        13421: begin
            cosine_reg0 <= 36'sb1101011110000111101010111110011111;
            sine_reg0   <= 36'sb100010111110010011001000010101110111;
        end
        13422: begin
            cosine_reg0 <= 36'sb1101011110110101010000110010010110;
            sine_reg0   <= 36'sb100010111110101000010011000111011010;
        end
        13423: begin
            cosine_reg0 <= 36'sb1101011111100010110110000100111100;
            sine_reg0   <= 36'sb100010111110111101011111000000100100;
        end
        13424: begin
            cosine_reg0 <= 36'sb1101100000010000011010110110001111;
            sine_reg0   <= 36'sb100010111111010010101100000001010100;
        end
        13425: begin
            cosine_reg0 <= 36'sb1101100000111101111111000110001110;
            sine_reg0   <= 36'sb100010111111100111111010001001101010;
        end
        13426: begin
            cosine_reg0 <= 36'sb1101100001101011100010110100110111;
            sine_reg0   <= 36'sb100010111111111101001001011001100011;
        end
        13427: begin
            cosine_reg0 <= 36'sb1101100010011001000110000010001000;
            sine_reg0   <= 36'sb100011000000010010011001110001000001;
        end
        13428: begin
            cosine_reg0 <= 36'sb1101100011000110101000101101111111;
            sine_reg0   <= 36'sb100011000000100111101011010000000001;
        end
        13429: begin
            cosine_reg0 <= 36'sb1101100011110100001010111000011010;
            sine_reg0   <= 36'sb100011000000111100111101110110100011;
        end
        13430: begin
            cosine_reg0 <= 36'sb1101100100100001101100100001011000;
            sine_reg0   <= 36'sb100011000001010010010001100100100111;
        end
        13431: begin
            cosine_reg0 <= 36'sb1101100101001111001101101000111000;
            sine_reg0   <= 36'sb100011000001100111100110011010001010;
        end
        13432: begin
            cosine_reg0 <= 36'sb1101100101111100101110001110110110;
            sine_reg0   <= 36'sb100011000001111100111100010111001101;
        end
        13433: begin
            cosine_reg0 <= 36'sb1101100110101010001110010011010010;
            sine_reg0   <= 36'sb100011000010010010010011011011101111;
        end
        13434: begin
            cosine_reg0 <= 36'sb1101100111010111101101110110001010;
            sine_reg0   <= 36'sb100011000010100111101011100111101111;
        end
        13435: begin
            cosine_reg0 <= 36'sb1101101000000101001100110111011011;
            sine_reg0   <= 36'sb100011000010111101000100111011001100;
        end
        13436: begin
            cosine_reg0 <= 36'sb1101101000110010101011010111000101;
            sine_reg0   <= 36'sb100011000011010010011111010110000100;
        end
        13437: begin
            cosine_reg0 <= 36'sb1101101001100000001001010101000101;
            sine_reg0   <= 36'sb100011000011100111111010111000011001;
        end
        13438: begin
            cosine_reg0 <= 36'sb1101101010001101100110110001011010;
            sine_reg0   <= 36'sb100011000011111101010111100010001000;
        end
        13439: begin
            cosine_reg0 <= 36'sb1101101010111011000011101100000011;
            sine_reg0   <= 36'sb100011000100010010110101010011010000;
        end
        13440: begin
            cosine_reg0 <= 36'sb1101101011101000100000000100111100;
            sine_reg0   <= 36'sb100011000100101000010100001011110010;
        end
        13441: begin
            cosine_reg0 <= 36'sb1101101100010101111011111100000100;
            sine_reg0   <= 36'sb100011000100111101110100001011101011;
        end
        13442: begin
            cosine_reg0 <= 36'sb1101101101000011010111010001011011;
            sine_reg0   <= 36'sb100011000101010011010101010010111100;
        end
        13443: begin
            cosine_reg0 <= 36'sb1101101101110000110010000100111101;
            sine_reg0   <= 36'sb100011000101101000110111100001100011;
        end
        13444: begin
            cosine_reg0 <= 36'sb1101101110011110001100010110101010;
            sine_reg0   <= 36'sb100011000101111110011010110111100000;
        end
        13445: begin
            cosine_reg0 <= 36'sb1101101111001011100110000110011111;
            sine_reg0   <= 36'sb100011000110010011111111010100110010;
        end
        13446: begin
            cosine_reg0 <= 36'sb1101101111111000111111010100011011;
            sine_reg0   <= 36'sb100011000110101001100100111001010111;
        end
        13447: begin
            cosine_reg0 <= 36'sb1101110000100110011000000000011011;
            sine_reg0   <= 36'sb100011000110111111001011100101010000;
        end
        13448: begin
            cosine_reg0 <= 36'sb1101110001010011110000001010011111;
            sine_reg0   <= 36'sb100011000111010100110011011000011010;
        end
        13449: begin
            cosine_reg0 <= 36'sb1101110010000001000111110010100101;
            sine_reg0   <= 36'sb100011000111101010011100010010110111;
        end
        13450: begin
            cosine_reg0 <= 36'sb1101110010101110011110111000101010;
            sine_reg0   <= 36'sb100011001000000000000110010100100100;
        end
        13451: begin
            cosine_reg0 <= 36'sb1101110011011011110101011100101101;
            sine_reg0   <= 36'sb100011001000010101110001011101100000;
        end
        13452: begin
            cosine_reg0 <= 36'sb1101110100001001001011011110101100;
            sine_reg0   <= 36'sb100011001000101011011101101101101100;
        end
        13453: begin
            cosine_reg0 <= 36'sb1101110100110110100000111110100110;
            sine_reg0   <= 36'sb100011001001000001001011000101000101;
        end
        13454: begin
            cosine_reg0 <= 36'sb1101110101100011110101111100011000;
            sine_reg0   <= 36'sb100011001001010110111001100011101100;
        end
        13455: begin
            cosine_reg0 <= 36'sb1101110110010001001010011000000010;
            sine_reg0   <= 36'sb100011001001101100101001001001011111;
        end
        13456: begin
            cosine_reg0 <= 36'sb1101110110111110011110010001100000;
            sine_reg0   <= 36'sb100011001010000010011001110110011110;
        end
        13457: begin
            cosine_reg0 <= 36'sb1101110111101011110001101000110010;
            sine_reg0   <= 36'sb100011001010011000001011101010101000;
        end
        13458: begin
            cosine_reg0 <= 36'sb1101111000011001000100011101110110;
            sine_reg0   <= 36'sb100011001010101101111110100101111011;
        end
        13459: begin
            cosine_reg0 <= 36'sb1101111001000110010110110000101010;
            sine_reg0   <= 36'sb100011001011000011110010101000011000;
        end
        13460: begin
            cosine_reg0 <= 36'sb1101111001110011101000100001001100;
            sine_reg0   <= 36'sb100011001011011001100111110001111100;
        end
        13461: begin
            cosine_reg0 <= 36'sb1101111010100000111001101111011010;
            sine_reg0   <= 36'sb100011001011101111011110000010101000;
        end
        13462: begin
            cosine_reg0 <= 36'sb1101111011001110001010011011010100;
            sine_reg0   <= 36'sb100011001100000101010101011010011011;
        end
        13463: begin
            cosine_reg0 <= 36'sb1101111011111011011010100100110110;
            sine_reg0   <= 36'sb100011001100011011001101111001010011;
        end
        13464: begin
            cosine_reg0 <= 36'sb1101111100101000101010001100000000;
            sine_reg0   <= 36'sb100011001100110001000111011111010000;
        end
        13465: begin
            cosine_reg0 <= 36'sb1101111101010101111001010000101111;
            sine_reg0   <= 36'sb100011001101000111000010001100010001;
        end
        13466: begin
            cosine_reg0 <= 36'sb1101111110000011000111110011000001;
            sine_reg0   <= 36'sb100011001101011100111110000000010110;
        end
        13467: begin
            cosine_reg0 <= 36'sb1101111110110000010101110010110110;
            sine_reg0   <= 36'sb100011001101110010111010111011011100;
        end
        13468: begin
            cosine_reg0 <= 36'sb1101111111011101100011010000001011;
            sine_reg0   <= 36'sb100011001110001000111000111101100100;
        end
        13469: begin
            cosine_reg0 <= 36'sb1110000000001010110000001010111111;
            sine_reg0   <= 36'sb100011001110011110111000000110101101;
        end
        13470: begin
            cosine_reg0 <= 36'sb1110000000110111111100100011001111;
            sine_reg0   <= 36'sb100011001110110100111000010110110101;
        end
        13471: begin
            cosine_reg0 <= 36'sb1110000001100101001000011000111011;
            sine_reg0   <= 36'sb100011001111001010111001101101111100;
        end
        13472: begin
            cosine_reg0 <= 36'sb1110000010010010010011101100000000;
            sine_reg0   <= 36'sb100011001111100000111100001100000010;
        end
        13473: begin
            cosine_reg0 <= 36'sb1110000010111111011110011100011100;
            sine_reg0   <= 36'sb100011001111110110111111110001000100;
        end
        13474: begin
            cosine_reg0 <= 36'sb1110000011101100101000101010001110;
            sine_reg0   <= 36'sb100011010000001101000100011101000011;
        end
        13475: begin
            cosine_reg0 <= 36'sb1110000100011001110010010101010101;
            sine_reg0   <= 36'sb100011010000100011001010001111111110;
        end
        13476: begin
            cosine_reg0 <= 36'sb1110000101000110111011011101101101;
            sine_reg0   <= 36'sb100011010000111001010001001001110011;
        end
        13477: begin
            cosine_reg0 <= 36'sb1110000101110100000100000011010110;
            sine_reg0   <= 36'sb100011010001001111011001001010100010;
        end
        13478: begin
            cosine_reg0 <= 36'sb1110000110100001001100000110001111;
            sine_reg0   <= 36'sb100011010001100101100010010010001001;
        end
        13479: begin
            cosine_reg0 <= 36'sb1110000111001110010011100110010100;
            sine_reg0   <= 36'sb100011010001111011101100100000101001;
        end
        13480: begin
            cosine_reg0 <= 36'sb1110000111111011011010100011100100;
            sine_reg0   <= 36'sb100011010010010001110111110110000001;
        end
        13481: begin
            cosine_reg0 <= 36'sb1110001000101000100000111101111111;
            sine_reg0   <= 36'sb100011010010101000000100010010001110;
        end
        13482: begin
            cosine_reg0 <= 36'sb1110001001010101100110110101100001;
            sine_reg0   <= 36'sb100011010010111110010001110101010001;
        end
        13483: begin
            cosine_reg0 <= 36'sb1110001010000010101100001010001001;
            sine_reg0   <= 36'sb100011010011010100100000011111001001;
        end
        13484: begin
            cosine_reg0 <= 36'sb1110001010101111110000111011110110;
            sine_reg0   <= 36'sb100011010011101010110000001111110101;
        end
        13485: begin
            cosine_reg0 <= 36'sb1110001011011100110101001010100101;
            sine_reg0   <= 36'sb100011010100000001000001000111010100;
        end
        13486: begin
            cosine_reg0 <= 36'sb1110001100001001111000110110010110;
            sine_reg0   <= 36'sb100011010100010111010011000101100100;
        end
        13487: begin
            cosine_reg0 <= 36'sb1110001100110110111011111111000101;
            sine_reg0   <= 36'sb100011010100101101100110001010100110;
        end
        13488: begin
            cosine_reg0 <= 36'sb1110001101100011111110100100110010;
            sine_reg0   <= 36'sb100011010101000011111010010110011001;
        end
        13489: begin
            cosine_reg0 <= 36'sb1110001110010001000000100111011011;
            sine_reg0   <= 36'sb100011010101011010001111101000111011;
        end
        13490: begin
            cosine_reg0 <= 36'sb1110001110111110000010000110111110;
            sine_reg0   <= 36'sb100011010101110000100110000010001011;
        end
        13491: begin
            cosine_reg0 <= 36'sb1110001111101011000011000011011001;
            sine_reg0   <= 36'sb100011010110000110111101100010001010;
        end
        13492: begin
            cosine_reg0 <= 36'sb1110010000011000000011011100101011;
            sine_reg0   <= 36'sb100011010110011101010110001000110101;
        end
        13493: begin
            cosine_reg0 <= 36'sb1110010001000101000011010010110001;
            sine_reg0   <= 36'sb100011010110110011101111110110001100;
        end
        13494: begin
            cosine_reg0 <= 36'sb1110010001110010000010100101101011;
            sine_reg0   <= 36'sb100011010111001010001010101010001111;
        end
        13495: begin
            cosine_reg0 <= 36'sb1110010010011111000001010101010110;
            sine_reg0   <= 36'sb100011010111100000100110100100111100;
        end
        13496: begin
            cosine_reg0 <= 36'sb1110010011001011111111100001110000;
            sine_reg0   <= 36'sb100011010111110111000011100110010010;
        end
        13497: begin
            cosine_reg0 <= 36'sb1110010011111000111101001010111001;
            sine_reg0   <= 36'sb100011011000001101100001101110010010;
        end
        13498: begin
            cosine_reg0 <= 36'sb1110010100100101111010010000101101;
            sine_reg0   <= 36'sb100011011000100100000000111100111000;
        end
        13499: begin
            cosine_reg0 <= 36'sb1110010101010010110110110011001100;
            sine_reg0   <= 36'sb100011011000111010100001010010000110;
        end
        13500: begin
            cosine_reg0 <= 36'sb1110010101111111110010110010010100;
            sine_reg0   <= 36'sb100011011001010001000010101101111010;
        end
        13501: begin
            cosine_reg0 <= 36'sb1110010110101100101110001110000010;
            sine_reg0   <= 36'sb100011011001100111100101010000010011;
        end
        13502: begin
            cosine_reg0 <= 36'sb1110010111011001101001000110010110;
            sine_reg0   <= 36'sb100011011001111110001000111001010000;
        end
        13503: begin
            cosine_reg0 <= 36'sb1110011000000110100011011011001101;
            sine_reg0   <= 36'sb100011011010010100101101101000110001;
        end
        13504: begin
            cosine_reg0 <= 36'sb1110011000110011011101001100100110;
            sine_reg0   <= 36'sb100011011010101011010011011110110100;
        end
        13505: begin
            cosine_reg0 <= 36'sb1110011001100000010110011010011111;
            sine_reg0   <= 36'sb100011011011000001111010011011011001;
        end
        13506: begin
            cosine_reg0 <= 36'sb1110011010001101001111000100110110;
            sine_reg0   <= 36'sb100011011011011000100010011110011110;
        end
        13507: begin
            cosine_reg0 <= 36'sb1110011010111010000111001011101010;
            sine_reg0   <= 36'sb100011011011101111001011101000000100;
        end
        13508: begin
            cosine_reg0 <= 36'sb1110011011100110111110101110111000;
            sine_reg0   <= 36'sb100011011100000101110101111000001001;
        end
        13509: begin
            cosine_reg0 <= 36'sb1110011100010011110101101110100000;
            sine_reg0   <= 36'sb100011011100011100100001001110101011;
        end
        13510: begin
            cosine_reg0 <= 36'sb1110011101000000101100001010011111;
            sine_reg0   <= 36'sb100011011100110011001101101011101100;
        end
        13511: begin
            cosine_reg0 <= 36'sb1110011101101101100010000010110011;
            sine_reg0   <= 36'sb100011011101001001111011001111001000;
        end
        13512: begin
            cosine_reg0 <= 36'sb1110011110011010010111010111011100;
            sine_reg0   <= 36'sb100011011101100000101001111001000000;
        end
        13513: begin
            cosine_reg0 <= 36'sb1110011111000111001100001000010110;
            sine_reg0   <= 36'sb100011011101110111011001101001010011;
        end
        13514: begin
            cosine_reg0 <= 36'sb1110011111110100000000010101100010;
            sine_reg0   <= 36'sb100011011110001110001010100000000000;
        end
        13515: begin
            cosine_reg0 <= 36'sb1110100000100000110011111110111011;
            sine_reg0   <= 36'sb100011011110100100111100011101000101;
        end
        13516: begin
            cosine_reg0 <= 36'sb1110100001001101100111000100100010;
            sine_reg0   <= 36'sb100011011110111011101111100000100011;
        end
        13517: begin
            cosine_reg0 <= 36'sb1110100001111010011001100110010100;
            sine_reg0   <= 36'sb100011011111010010100011101010011000;
        end
        13518: begin
            cosine_reg0 <= 36'sb1110100010100111001011100100010000;
            sine_reg0   <= 36'sb100011011111101001011000111010100011;
        end
        13519: begin
            cosine_reg0 <= 36'sb1110100011010011111100111110010011;
            sine_reg0   <= 36'sb100011100000000000001111010001000011;
        end
        13520: begin
            cosine_reg0 <= 36'sb1110100100000000101101110100011101;
            sine_reg0   <= 36'sb100011100000010111000110101101111000;
        end
        13521: begin
            cosine_reg0 <= 36'sb1110100100101101011110000110101011;
            sine_reg0   <= 36'sb100011100000101101111111010001000001;
        end
        13522: begin
            cosine_reg0 <= 36'sb1110100101011010001101110100111011;
            sine_reg0   <= 36'sb100011100001000100111000111010011100;
        end
        13523: begin
            cosine_reg0 <= 36'sb1110100110000110111100111111001100;
            sine_reg0   <= 36'sb100011100001011011110011101010001001;
        end
        13524: begin
            cosine_reg0 <= 36'sb1110100110110011101011100101011101;
            sine_reg0   <= 36'sb100011100001110010101111100000001000;
        end
        13525: begin
            cosine_reg0 <= 36'sb1110100111100000011001100111101011;
            sine_reg0   <= 36'sb100011100010001001101100011100010110;
        end
        13526: begin
            cosine_reg0 <= 36'sb1110101000001101000111000101110101;
            sine_reg0   <= 36'sb100011100010100000101010011110110100;
        end
        13527: begin
            cosine_reg0 <= 36'sb1110101000111001110011111111111001;
            sine_reg0   <= 36'sb100011100010110111101001100111100000;
        end
        13528: begin
            cosine_reg0 <= 36'sb1110101001100110100000010101110101;
            sine_reg0   <= 36'sb100011100011001110101001110110011001;
        end
        13529: begin
            cosine_reg0 <= 36'sb1110101010010011001100000111100111;
            sine_reg0   <= 36'sb100011100011100101101011001011011111;
        end
        13530: begin
            cosine_reg0 <= 36'sb1110101010111111110111010101001111;
            sine_reg0   <= 36'sb100011100011111100101101100110110001;
        end
        13531: begin
            cosine_reg0 <= 36'sb1110101011101100100001111110101001;
            sine_reg0   <= 36'sb100011100100010011110001001000001101;
        end
        13532: begin
            cosine_reg0 <= 36'sb1110101100011001001100000011110101;
            sine_reg0   <= 36'sb100011100100101010110101101111110100;
        end
        13533: begin
            cosine_reg0 <= 36'sb1110101101000101110101100100110001;
            sine_reg0   <= 36'sb100011100101000001111011011101100011;
        end
        13534: begin
            cosine_reg0 <= 36'sb1110101101110010011110100001011010;
            sine_reg0   <= 36'sb100011100101011001000010010001011011;
        end
        13535: begin
            cosine_reg0 <= 36'sb1110101110011111000110111001110000;
            sine_reg0   <= 36'sb100011100101110000001010001011011010;
        end
        13536: begin
            cosine_reg0 <= 36'sb1110101111001011101110101101110000;
            sine_reg0   <= 36'sb100011100110000111010011001011011111;
        end
        13537: begin
            cosine_reg0 <= 36'sb1110101111111000010101111101011001;
            sine_reg0   <= 36'sb100011100110011110011101010001101001;
        end
        13538: begin
            cosine_reg0 <= 36'sb1110110000100100111100101000101010;
            sine_reg0   <= 36'sb100011100110110101101000011101111001;
        end
        13539: begin
            cosine_reg0 <= 36'sb1110110001010001100010101111011111;
            sine_reg0   <= 36'sb100011100111001100110100110000001011;
        end
        13540: begin
            cosine_reg0 <= 36'sb1110110001111110001000010001111000;
            sine_reg0   <= 36'sb100011100111100100000010001000100001;
        end
        13541: begin
            cosine_reg0 <= 36'sb1110110010101010101101001111110011;
            sine_reg0   <= 36'sb100011100111111011010000100110111000;
        end
        13542: begin
            cosine_reg0 <= 36'sb1110110011010111010001101001001111;
            sine_reg0   <= 36'sb100011101000010010100000001011010001;
        end
        13543: begin
            cosine_reg0 <= 36'sb1110110100000011110101011110001000;
            sine_reg0   <= 36'sb100011101000101001110000110101101001;
        end
        13544: begin
            cosine_reg0 <= 36'sb1110110100110000011000101110011111;
            sine_reg0   <= 36'sb100011101001000001000010100110000001;
        end
        13545: begin
            cosine_reg0 <= 36'sb1110110101011100111011011010010000;
            sine_reg0   <= 36'sb100011101001011000010101011100010111;
        end
        13546: begin
            cosine_reg0 <= 36'sb1110110110001001011101100001011011;
            sine_reg0   <= 36'sb100011101001101111101001011000101011;
        end
        13547: begin
            cosine_reg0 <= 36'sb1110110110110101111111000011111110;
            sine_reg0   <= 36'sb100011101010000110111110011010111011;
        end
        13548: begin
            cosine_reg0 <= 36'sb1110110111100010100000000001110110;
            sine_reg0   <= 36'sb100011101010011110010100100011000110;
        end
        13549: begin
            cosine_reg0 <= 36'sb1110111000001111000000011011000010;
            sine_reg0   <= 36'sb100011101010110101101011110001001100;
        end
        13550: begin
            cosine_reg0 <= 36'sb1110111000111011100000001111100001;
            sine_reg0   <= 36'sb100011101011001101000100000101001100;
        end
        13551: begin
            cosine_reg0 <= 36'sb1110111001100111111111011111010001;
            sine_reg0   <= 36'sb100011101011100100011101011111000101;
        end
        13552: begin
            cosine_reg0 <= 36'sb1110111010010100011110001010010000;
            sine_reg0   <= 36'sb100011101011111011110111111110110110;
        end
        13553: begin
            cosine_reg0 <= 36'sb1110111011000000111100010000011100;
            sine_reg0   <= 36'sb100011101100010011010011100100011110;
        end
        13554: begin
            cosine_reg0 <= 36'sb1110111011101101011001110001110011;
            sine_reg0   <= 36'sb100011101100101010110000001111111100;
        end
        13555: begin
            cosine_reg0 <= 36'sb1110111100011001110110101110010101;
            sine_reg0   <= 36'sb100011101101000010001110000001010000;
        end
        13556: begin
            cosine_reg0 <= 36'sb1110111101000110010011000101111111;
            sine_reg0   <= 36'sb100011101101011001101100111000010111;
        end
        13557: begin
            cosine_reg0 <= 36'sb1110111101110010101110111000101111;
            sine_reg0   <= 36'sb100011101101110001001100110101010011;
        end
        13558: begin
            cosine_reg0 <= 36'sb1110111110011111001010000110100100;
            sine_reg0   <= 36'sb100011101110001000101101111000000001;
        end
        13559: begin
            cosine_reg0 <= 36'sb1110111111001011100100101111011011;
            sine_reg0   <= 36'sb100011101110100000010000000000100000;
        end
        13560: begin
            cosine_reg0 <= 36'sb1110111111110111111110110011010101;
            sine_reg0   <= 36'sb100011101110110111110011001110110000;
        end
        13561: begin
            cosine_reg0 <= 36'sb1111000000100100011000010010001110;
            sine_reg0   <= 36'sb100011101111001111010111100010110001;
        end
        13562: begin
            cosine_reg0 <= 36'sb1111000001010000110001001100000100;
            sine_reg0   <= 36'sb100011101111100110111100111100100000;
        end
        13563: begin
            cosine_reg0 <= 36'sb1111000001111101001001100000110111;
            sine_reg0   <= 36'sb100011101111111110100011011011111101;
        end
        13564: begin
            cosine_reg0 <= 36'sb1111000010101001100001010000100100;
            sine_reg0   <= 36'sb100011110000010110001011000001000111;
        end
        13565: begin
            cosine_reg0 <= 36'sb1111000011010101111000011011001011;
            sine_reg0   <= 36'sb100011110000101101110011101011111101;
        end
        13566: begin
            cosine_reg0 <= 36'sb1111000100000010001111000000101000;
            sine_reg0   <= 36'sb100011110001000101011101011100011111;
        end
        13567: begin
            cosine_reg0 <= 36'sb1111000100101110100101000000111010;
            sine_reg0   <= 36'sb100011110001011101001000010010101011;
        end
        13568: begin
            cosine_reg0 <= 36'sb1111000101011010111010011100000000;
            sine_reg0   <= 36'sb100011110001110100110100001110100001;
        end
        13569: begin
            cosine_reg0 <= 36'sb1111000110000111001111010001111000;
            sine_reg0   <= 36'sb100011110010001100100001001111111111;
        end
        13570: begin
            cosine_reg0 <= 36'sb1111000110110011100011100010100001;
            sine_reg0   <= 36'sb100011110010100100001111010111000101;
        end
        13571: begin
            cosine_reg0 <= 36'sb1111000111011111110111001101110111;
            sine_reg0   <= 36'sb100011110010111011111110100011110001;
        end
        13572: begin
            cosine_reg0 <= 36'sb1111001000001100001010010011111011;
            sine_reg0   <= 36'sb100011110011010011101110110110000011;
        end
        13573: begin
            cosine_reg0 <= 36'sb1111001000111000011100110100101010;
            sine_reg0   <= 36'sb100011110011101011100000001101111011;
        end
        13574: begin
            cosine_reg0 <= 36'sb1111001001100100101110110000000010;
            sine_reg0   <= 36'sb100011110100000011010010101011010110;
        end
        13575: begin
            cosine_reg0 <= 36'sb1111001010010001000000000110000001;
            sine_reg0   <= 36'sb100011110100011011000110001110010100;
        end
        13576: begin
            cosine_reg0 <= 36'sb1111001010111101010000110110100111;
            sine_reg0   <= 36'sb100011110100110010111010110110110100;
        end
        13577: begin
            cosine_reg0 <= 36'sb1111001011101001100001000001110001;
            sine_reg0   <= 36'sb100011110101001010110000100100110110;
        end
        13578: begin
            cosine_reg0 <= 36'sb1111001100010101110000100111011110;
            sine_reg0   <= 36'sb100011110101100010100111011000011000;
        end
        13579: begin
            cosine_reg0 <= 36'sb1111001101000001111111100111101011;
            sine_reg0   <= 36'sb100011110101111010011111010001011001;
        end
        13580: begin
            cosine_reg0 <= 36'sb1111001101101110001110000010010111;
            sine_reg0   <= 36'sb100011110110010010011000001111111001;
        end
        13581: begin
            cosine_reg0 <= 36'sb1111001110011010011011110111100001;
            sine_reg0   <= 36'sb100011110110101010010010010011110110;
        end
        13582: begin
            cosine_reg0 <= 36'sb1111001111000110101001000111000111;
            sine_reg0   <= 36'sb100011110111000010001101011101010000;
        end
        13583: begin
            cosine_reg0 <= 36'sb1111001111110010110101110001000111;
            sine_reg0   <= 36'sb100011110111011010001001101100000110;
        end
        13584: begin
            cosine_reg0 <= 36'sb1111010000011111000001110101011111;
            sine_reg0   <= 36'sb100011110111110010000111000000010111;
        end
        13585: begin
            cosine_reg0 <= 36'sb1111010001001011001101010100001101;
            sine_reg0   <= 36'sb100011111000001010000101011010000001;
        end
        13586: begin
            cosine_reg0 <= 36'sb1111010001110111011000001101010001;
            sine_reg0   <= 36'sb100011111000100010000100111001000100;
        end
        13587: begin
            cosine_reg0 <= 36'sb1111010010100011100010100000100111;
            sine_reg0   <= 36'sb100011111000111010000101011101011111;
        end
        13588: begin
            cosine_reg0 <= 36'sb1111010011001111101100001110010000;
            sine_reg0   <= 36'sb100011111001010010000111000111010010;
        end
        13589: begin
            cosine_reg0 <= 36'sb1111010011111011110101010110001000;
            sine_reg0   <= 36'sb100011111001101010001001110110011010;
        end
        13590: begin
            cosine_reg0 <= 36'sb1111010100100111111101111000001110;
            sine_reg0   <= 36'sb100011111010000010001101101010111000;
        end
        13591: begin
            cosine_reg0 <= 36'sb1111010101010100000101110100100001;
            sine_reg0   <= 36'sb100011111010011010010010100100101010;
        end
        13592: begin
            cosine_reg0 <= 36'sb1111010110000000001101001010111110;
            sine_reg0   <= 36'sb100011111010110010011000100011101111;
        end
        13593: begin
            cosine_reg0 <= 36'sb1111010110101100010011111011100100;
            sine_reg0   <= 36'sb100011111011001010011111101000000111;
        end
        13594: begin
            cosine_reg0 <= 36'sb1111010111011000011010000110010010;
            sine_reg0   <= 36'sb100011111011100010100111110001110000;
        end
        13595: begin
            cosine_reg0 <= 36'sb1111011000000100011111101011000101;
            sine_reg0   <= 36'sb100011111011111010110001000000101010;
        end
        13596: begin
            cosine_reg0 <= 36'sb1111011000110000100100101001111100;
            sine_reg0   <= 36'sb100011111100010010111011010100110100;
        end
        13597: begin
            cosine_reg0 <= 36'sb1111011001011100101001000010110101;
            sine_reg0   <= 36'sb100011111100101011000110101110001100;
        end
        13598: begin
            cosine_reg0 <= 36'sb1111011010001000101100110101101111;
            sine_reg0   <= 36'sb100011111101000011010011001100110010;
        end
        13599: begin
            cosine_reg0 <= 36'sb1111011010110100110000000010101000;
            sine_reg0   <= 36'sb100011111101011011100000110000100101;
        end
        13600: begin
            cosine_reg0 <= 36'sb1111011011100000110010101001011101;
            sine_reg0   <= 36'sb100011111101110011101111011001100100;
        end
        13601: begin
            cosine_reg0 <= 36'sb1111011100001100110100101010001111;
            sine_reg0   <= 36'sb100011111110001011111111000111101110;
        end
        13602: begin
            cosine_reg0 <= 36'sb1111011100111000110110000100111001;
            sine_reg0   <= 36'sb100011111110100100001111111011000010;
        end
        13603: begin
            cosine_reg0 <= 36'sb1111011101100100110110111001011100;
            sine_reg0   <= 36'sb100011111110111100100001110011011111;
        end
        13604: begin
            cosine_reg0 <= 36'sb1111011110010000110111000111110101;
            sine_reg0   <= 36'sb100011111111010100110100110001000100;
        end
        13605: begin
            cosine_reg0 <= 36'sb1111011110111100110110110000000011;
            sine_reg0   <= 36'sb100011111111101101001000110011110001;
        end
        13606: begin
            cosine_reg0 <= 36'sb1111011111101000110101110010000100;
            sine_reg0   <= 36'sb100100000000000101011101111011100100;
        end
        13607: begin
            cosine_reg0 <= 36'sb1111100000010100110100001101110110;
            sine_reg0   <= 36'sb100100000000011101110100001000011100;
        end
        13608: begin
            cosine_reg0 <= 36'sb1111100001000000110010000011011000;
            sine_reg0   <= 36'sb100100000000110110001011011010011000;
        end
        13609: begin
            cosine_reg0 <= 36'sb1111100001101100101111010010100111;
            sine_reg0   <= 36'sb100100000001001110100011110001011001;
        end
        13610: begin
            cosine_reg0 <= 36'sb1111100010011000101011111011100010;
            sine_reg0   <= 36'sb100100000001100110111101001101011011;
        end
        13611: begin
            cosine_reg0 <= 36'sb1111100011000100100111111110001000;
            sine_reg0   <= 36'sb100100000001111111010111101110011111;
        end
        13612: begin
            cosine_reg0 <= 36'sb1111100011110000100011011010010111;
            sine_reg0   <= 36'sb100100000010010111110011010100100100;
        end
        13613: begin
            cosine_reg0 <= 36'sb1111100100011100011110010000001101;
            sine_reg0   <= 36'sb100100000010110000001111111111101001;
        end
        13614: begin
            cosine_reg0 <= 36'sb1111100101001000011000011111101000;
            sine_reg0   <= 36'sb100100000011001000101101101111101101;
        end
        13615: begin
            cosine_reg0 <= 36'sb1111100101110100010010001000100111;
            sine_reg0   <= 36'sb100100000011100001001100100100101110;
        end
        13616: begin
            cosine_reg0 <= 36'sb1111100110100000001011001011000111;
            sine_reg0   <= 36'sb100100000011111001101100011110101100;
        end
        13617: begin
            cosine_reg0 <= 36'sb1111100111001100000011100111001001;
            sine_reg0   <= 36'sb100100000100010010001101011101100110;
        end
        13618: begin
            cosine_reg0 <= 36'sb1111100111110111111011011100101000;
            sine_reg0   <= 36'sb100100000100101010101111100001011011;
        end
        13619: begin
            cosine_reg0 <= 36'sb1111101000100011110010101011100101;
            sine_reg0   <= 36'sb100100000101000011010010101010001011;
        end
        13620: begin
            cosine_reg0 <= 36'sb1111101001001111101001010011111101;
            sine_reg0   <= 36'sb100100000101011011110110110111110011;
        end
        13621: begin
            cosine_reg0 <= 36'sb1111101001111011011111010101101110;
            sine_reg0   <= 36'sb100100000101110100011100001010010011;
        end
        13622: begin
            cosine_reg0 <= 36'sb1111101010100111010100110000110111;
            sine_reg0   <= 36'sb100100000110001101000010100001101011;
        end
        13623: begin
            cosine_reg0 <= 36'sb1111101011010011001001100101010111;
            sine_reg0   <= 36'sb100100000110100101101001111101111001;
        end
        13624: begin
            cosine_reg0 <= 36'sb1111101011111110111101110011001010;
            sine_reg0   <= 36'sb100100000110111110010010011110111101;
        end
        13625: begin
            cosine_reg0 <= 36'sb1111101100101010110001011010010001;
            sine_reg0   <= 36'sb100100000111010110111100000100110100;
        end
        13626: begin
            cosine_reg0 <= 36'sb1111101101010110100100011010101001;
            sine_reg0   <= 36'sb100100000111101111100110101111011111;
        end
        13627: begin
            cosine_reg0 <= 36'sb1111101110000010010110110100010000;
            sine_reg0   <= 36'sb100100001000001000010010011110111101;
        end
        13628: begin
            cosine_reg0 <= 36'sb1111101110101110001000100111000100;
            sine_reg0   <= 36'sb100100001000100000111111010011001100;
        end
        13629: begin
            cosine_reg0 <= 36'sb1111101111011001111001110011000101;
            sine_reg0   <= 36'sb100100001000111001101101001100001100;
        end
        13630: begin
            cosine_reg0 <= 36'sb1111110000000101101010011000010000;
            sine_reg0   <= 36'sb100100001001010010011100001001111011;
        end
        13631: begin
            cosine_reg0 <= 36'sb1111110000110001011010010110100100;
            sine_reg0   <= 36'sb100100001001101011001100001100011001;
        end
        13632: begin
            cosine_reg0 <= 36'sb1111110001011101001001101101111111;
            sine_reg0   <= 36'sb100100001010000011111101010011100101;
        end
        13633: begin
            cosine_reg0 <= 36'sb1111110010001000111000011110011111;
            sine_reg0   <= 36'sb100100001010011100101111011111011101;
        end
        13634: begin
            cosine_reg0 <= 36'sb1111110010110100100110101000000010;
            sine_reg0   <= 36'sb100100001010110101100010110000000010;
        end
        13635: begin
            cosine_reg0 <= 36'sb1111110011100000010100001010100111;
            sine_reg0   <= 36'sb100100001011001110010111000101010001;
        end
        13636: begin
            cosine_reg0 <= 36'sb1111110100001100000001000110001101;
            sine_reg0   <= 36'sb100100001011100111001100011111001010;
        end
        13637: begin
            cosine_reg0 <= 36'sb1111110100110111101101011010110001;
            sine_reg0   <= 36'sb100100001100000000000010111101101100;
        end
        13638: begin
            cosine_reg0 <= 36'sb1111110101100011011001001000010010;
            sine_reg0   <= 36'sb100100001100011000111010100000110110;
        end
        13639: begin
            cosine_reg0 <= 36'sb1111110110001111000100001110101110;
            sine_reg0   <= 36'sb100100001100110001110011001000100111;
        end
        13640: begin
            cosine_reg0 <= 36'sb1111110110111010101110101110000100;
            sine_reg0   <= 36'sb100100001101001010101100110100111110;
        end
        13641: begin
            cosine_reg0 <= 36'sb1111110111100110011000100110010010;
            sine_reg0   <= 36'sb100100001101100011100111100101111010;
        end
        13642: begin
            cosine_reg0 <= 36'sb1111111000010010000001110111010101;
            sine_reg0   <= 36'sb100100001101111100100011011011011010;
        end
        13643: begin
            cosine_reg0 <= 36'sb1111111000111101101010100001001101;
            sine_reg0   <= 36'sb100100001110010101100000010101011101;
        end
        13644: begin
            cosine_reg0 <= 36'sb1111111001101001010010100011111000;
            sine_reg0   <= 36'sb100100001110101110011110010100000011;
        end
        13645: begin
            cosine_reg0 <= 36'sb1111111010010100111001111111010100;
            sine_reg0   <= 36'sb100100001111000111011101010111001010;
        end
        13646: begin
            cosine_reg0 <= 36'sb1111111011000000100000110011011111;
            sine_reg0   <= 36'sb100100001111100000011101011110110001;
        end
        13647: begin
            cosine_reg0 <= 36'sb1111111011101100000111000000011000;
            sine_reg0   <= 36'sb100100001111111001011110101010110111;
        end
        13648: begin
            cosine_reg0 <= 36'sb1111111100010111101100100101111100;
            sine_reg0   <= 36'sb100100010000010010100000111011011100;
        end
        13649: begin
            cosine_reg0 <= 36'sb1111111101000011010001100100001100;
            sine_reg0   <= 36'sb100100010000101011100100010000011110;
        end
        13650: begin
            cosine_reg0 <= 36'sb1111111101101110110101111011000011;
            sine_reg0   <= 36'sb100100010001000100101000101001111101;
        end
        13651: begin
            cosine_reg0 <= 36'sb1111111110011010011001101010100010;
            sine_reg0   <= 36'sb100100010001011101101110000111110111;
        end
        13652: begin
            cosine_reg0 <= 36'sb1111111111000101111100110010100110;
            sine_reg0   <= 36'sb100100010001110110110100101010001011;
        end
        13653: begin
            cosine_reg0 <= 36'sb1111111111110001011111010011001110;
            sine_reg0   <= 36'sb100100010010001111111100010000111001;
        end
        13654: begin
            cosine_reg0 <= 36'sb10000000000011101000001001100011000;
            sine_reg0   <= 36'sb100100010010101001000100111100000000;
        end
        13655: begin
            cosine_reg0 <= 36'sb10000000001001000100010011110000010;
            sine_reg0   <= 36'sb100100010011000010001110101011011110;
        end
        13656: begin
            cosine_reg0 <= 36'sb10000000001110100000011001000001010;
            sine_reg0   <= 36'sb100100010011011011011001011111010011;
        end
        13657: begin
            cosine_reg0 <= 36'sb10000000010011111100011001010110000;
            sine_reg0   <= 36'sb100100010011110100100101010111011110;
        end
        13658: begin
            cosine_reg0 <= 36'sb10000000011001011000010100101110001;
            sine_reg0   <= 36'sb100100010100001101110010010011111101;
        end
        13659: begin
            cosine_reg0 <= 36'sb10000000011110110100001011001001011;
            sine_reg0   <= 36'sb100100010100100111000000010100110000;
        end
        13660: begin
            cosine_reg0 <= 36'sb10000000100100001111111100100111101;
            sine_reg0   <= 36'sb100100010101000000001111011001110101;
        end
        13661: begin
            cosine_reg0 <= 36'sb10000000101001101011101001001000101;
            sine_reg0   <= 36'sb100100010101011001011111100011001101;
        end
        13662: begin
            cosine_reg0 <= 36'sb10000000101111000111010000101100010;
            sine_reg0   <= 36'sb100100010101110010110000110000110101;
        end
        13663: begin
            cosine_reg0 <= 36'sb10000000110100100010110011010010010;
            sine_reg0   <= 36'sb100100010110001100000011000010101101;
        end
        13664: begin
            cosine_reg0 <= 36'sb10000000111001111110010000111010011;
            sine_reg0   <= 36'sb100100010110100101010110011000110011;
        end
        13665: begin
            cosine_reg0 <= 36'sb10000000111111011001101001100100011;
            sine_reg0   <= 36'sb100100010110111110101010110011001000;
        end
        13666: begin
            cosine_reg0 <= 36'sb10000001000100110100111101010000001;
            sine_reg0   <= 36'sb100100010111011000000000010001101010;
        end
        13667: begin
            cosine_reg0 <= 36'sb10000001001010010000001011111101011;
            sine_reg0   <= 36'sb100100010111110001010110110100010111;
        end
        13668: begin
            cosine_reg0 <= 36'sb10000001001111101011010101101100000;
            sine_reg0   <= 36'sb100100011000001010101110011011001111;
        end
        13669: begin
            cosine_reg0 <= 36'sb10000001010101000110011010011011110;
            sine_reg0   <= 36'sb100100011000100100000111000110010010;
        end
        13670: begin
            cosine_reg0 <= 36'sb10000001011010100001011010001100011;
            sine_reg0   <= 36'sb100100011000111101100000110101011101;
        end
        13671: begin
            cosine_reg0 <= 36'sb10000001011111111100010100111101101;
            sine_reg0   <= 36'sb100100011001010110111011101000110000;
        end
        13672: begin
            cosine_reg0 <= 36'sb10000001100101010111001010101111011;
            sine_reg0   <= 36'sb100100011001110000010111100000001011;
        end
        13673: begin
            cosine_reg0 <= 36'sb10000001101010110001111011100001011;
            sine_reg0   <= 36'sb100100011010001001110100011011101011;
        end
        13674: begin
            cosine_reg0 <= 36'sb10000001110000001100100111010011100;
            sine_reg0   <= 36'sb100100011010100011010010011011010000;
        end
        13675: begin
            cosine_reg0 <= 36'sb10000001110101100111001110000101011;
            sine_reg0   <= 36'sb100100011010111100110001011110111010;
        end
        13676: begin
            cosine_reg0 <= 36'sb10000001111011000001101111110110111;
            sine_reg0   <= 36'sb100100011011010110010001100110100110;
        end
        13677: begin
            cosine_reg0 <= 36'sb10000010000000011100001100100111111;
            sine_reg0   <= 36'sb100100011011101111110010110010010101;
        end
        13678: begin
            cosine_reg0 <= 36'sb10000010000101110110100100011000001;
            sine_reg0   <= 36'sb100100011100001001010101000010000101;
        end
        13679: begin
            cosine_reg0 <= 36'sb10000010001011010000110111000111011;
            sine_reg0   <= 36'sb100100011100100010111000010101110101;
        end
        13680: begin
            cosine_reg0 <= 36'sb10000010010000101011000100110101011;
            sine_reg0   <= 36'sb100100011100111100011100101101100100;
        end
        13681: begin
            cosine_reg0 <= 36'sb10000010010110000101001101100010000;
            sine_reg0   <= 36'sb100100011101010110000010001001010001;
        end
        13682: begin
            cosine_reg0 <= 36'sb10000010011011011111010001001101000;
            sine_reg0   <= 36'sb100100011101101111101000101000111011;
        end
        13683: begin
            cosine_reg0 <= 36'sb10000010100000111001001111110110010;
            sine_reg0   <= 36'sb100100011110001001010000001100100010;
        end
        13684: begin
            cosine_reg0 <= 36'sb10000010100110010011001001011101011;
            sine_reg0   <= 36'sb100100011110100010111000110100000100;
        end
        13685: begin
            cosine_reg0 <= 36'sb10000010101011101100111110000010010;
            sine_reg0   <= 36'sb100100011110111100100010011111100000;
        end
        13686: begin
            cosine_reg0 <= 36'sb10000010110001000110101101100100110;
            sine_reg0   <= 36'sb100100011111010110001101001110110101;
        end
        13687: begin
            cosine_reg0 <= 36'sb10000010110110100000011000000100100;
            sine_reg0   <= 36'sb100100011111101111111001000010000010;
        end
        13688: begin
            cosine_reg0 <= 36'sb10000010111011111001111101100001100;
            sine_reg0   <= 36'sb100100100000001001100101111001000111;
        end
        13689: begin
            cosine_reg0 <= 36'sb10000011000001010011011101111011011;
            sine_reg0   <= 36'sb100100100000100011010011110100000010;
        end
        13690: begin
            cosine_reg0 <= 36'sb10000011000110101100111001010010000;
            sine_reg0   <= 36'sb100100100000111101000010110010110010;
        end
        13691: begin
            cosine_reg0 <= 36'sb10000011001100000110001111100101001;
            sine_reg0   <= 36'sb100100100001010110110010110101010111;
        end
        13692: begin
            cosine_reg0 <= 36'sb10000011010001011111100000110100100;
            sine_reg0   <= 36'sb100100100001110000100011111011101110;
        end
        13693: begin
            cosine_reg0 <= 36'sb10000011010110111000101101000000000;
            sine_reg0   <= 36'sb100100100010001010010110000101111001;
        end
        13694: begin
            cosine_reg0 <= 36'sb10000011011100010001110100000111011;
            sine_reg0   <= 36'sb100100100010100100001001010011110100;
        end
        13695: begin
            cosine_reg0 <= 36'sb10000011100001101010110110001010100;
            sine_reg0   <= 36'sb100100100010111101111101100101100000;
        end
        13696: begin
            cosine_reg0 <= 36'sb10000011100111000011110011001001000;
            sine_reg0   <= 36'sb100100100011010111110010111010111011;
        end
        13697: begin
            cosine_reg0 <= 36'sb10000011101100011100101011000010111;
            sine_reg0   <= 36'sb100100100011110001101001010100000100;
        end
        13698: begin
            cosine_reg0 <= 36'sb10000011110001110101011101110111110;
            sine_reg0   <= 36'sb100100100100001011100000110000111010;
        end
        13699: begin
            cosine_reg0 <= 36'sb10000011110111001110001011100111100;
            sine_reg0   <= 36'sb100100100100100101011001010001011101;
        end
        13700: begin
            cosine_reg0 <= 36'sb10000011111100100110110100010001110;
            sine_reg0   <= 36'sb100100100100111111010010110101101011;
        end
        13701: begin
            cosine_reg0 <= 36'sb10000100000001111111010111110110101;
            sine_reg0   <= 36'sb100100100101011001001101011101100100;
        end
        13702: begin
            cosine_reg0 <= 36'sb10000100000111010111110110010101101;
            sine_reg0   <= 36'sb100100100101110011001001001001000110;
        end
        13703: begin
            cosine_reg0 <= 36'sb10000100001100110000001111101110101;
            sine_reg0   <= 36'sb100100100110001101000101111000010000;
        end
        13704: begin
            cosine_reg0 <= 36'sb10000100010010001000100100000001100;
            sine_reg0   <= 36'sb100100100110100111000011101011000001;
        end
        13705: begin
            cosine_reg0 <= 36'sb10000100010111100000110011001110000;
            sine_reg0   <= 36'sb100100100111000001000010100001011001;
        end
        13706: begin
            cosine_reg0 <= 36'sb10000100011100111000111101010011111;
            sine_reg0   <= 36'sb100100100111011011000010011011010110;
        end
        13707: begin
            cosine_reg0 <= 36'sb10000100100010010001000010010010111;
            sine_reg0   <= 36'sb100100100111110101000011011000111000;
        end
        13708: begin
            cosine_reg0 <= 36'sb10000100100111101001000010001010111;
            sine_reg0   <= 36'sb100100101000001111000101011001111100;
        end
        13709: begin
            cosine_reg0 <= 36'sb10000100101101000000111100111011110;
            sine_reg0   <= 36'sb100100101000101001001000011110100011;
        end
        13710: begin
            cosine_reg0 <= 36'sb10000100110010011000110010100101001;
            sine_reg0   <= 36'sb100100101001000011001100100110101100;
        end
        13711: begin
            cosine_reg0 <= 36'sb10000100110111110000100011000110110;
            sine_reg0   <= 36'sb100100101001011101010001110010010100;
        end
        13712: begin
            cosine_reg0 <= 36'sb10000100111101001000001110100000101;
            sine_reg0   <= 36'sb100100101001110111011000000001011100;
        end
        13713: begin
            cosine_reg0 <= 36'sb10000101000010011111110100110010100;
            sine_reg0   <= 36'sb100100101010010001011111010100000011;
        end
        13714: begin
            cosine_reg0 <= 36'sb10000101000111110111010101111100001;
            sine_reg0   <= 36'sb100100101010101011100111101010000110;
        end
        13715: begin
            cosine_reg0 <= 36'sb10000101001101001110110001111101001;
            sine_reg0   <= 36'sb100100101011000101110001000011100110;
        end
        13716: begin
            cosine_reg0 <= 36'sb10000101010010100110001000110101101;
            sine_reg0   <= 36'sb100100101011011111111011100000100001;
        end
        13717: begin
            cosine_reg0 <= 36'sb10000101010111111101011010100101001;
            sine_reg0   <= 36'sb100100101011111010000111000000110110;
        end
        13718: begin
            cosine_reg0 <= 36'sb10000101011101010100100111001011101;
            sine_reg0   <= 36'sb100100101100010100010011100100100101;
        end
        13719: begin
            cosine_reg0 <= 36'sb10000101100010101011101110101000110;
            sine_reg0   <= 36'sb100100101100101110100001001011101011;
        end
        13720: begin
            cosine_reg0 <= 36'sb10000101101000000010110000111100011;
            sine_reg0   <= 36'sb100100101101001000101111110110001001;
        end
        13721: begin
            cosine_reg0 <= 36'sb10000101101101011001101110000110011;
            sine_reg0   <= 36'sb100100101101100010111111100011111101;
        end
        13722: begin
            cosine_reg0 <= 36'sb10000101110010110000100110000110011;
            sine_reg0   <= 36'sb100100101101111101010000010101000111;
        end
        13723: begin
            cosine_reg0 <= 36'sb10000101111000000111011000111100011;
            sine_reg0   <= 36'sb100100101110010111100010001001100100;
        end
        13724: begin
            cosine_reg0 <= 36'sb10000101111101011110000110100111111;
            sine_reg0   <= 36'sb100100101110110001110101000001010101;
        end
        13725: begin
            cosine_reg0 <= 36'sb10000110000010110100101111001001000;
            sine_reg0   <= 36'sb100100101111001100001000111100011000;
        end
        13726: begin
            cosine_reg0 <= 36'sb10000110001000001011010010011111010;
            sine_reg0   <= 36'sb100100101111100110011101111010101100;
        end
        13727: begin
            cosine_reg0 <= 36'sb10000110001101100001110000101010101;
            sine_reg0   <= 36'sb100100110000000000110011111100010000;
        end
        13728: begin
            cosine_reg0 <= 36'sb10000110010010111000001001101010111;
            sine_reg0   <= 36'sb100100110000011011001011000001000100;
        end
        13729: begin
            cosine_reg0 <= 36'sb10000110011000001110011101011111110;
            sine_reg0   <= 36'sb100100110000110101100011001001000101;
        end
        13730: begin
            cosine_reg0 <= 36'sb10000110011101100100101100001001000;
            sine_reg0   <= 36'sb100100110001001111111100010100010011;
        end
        13731: begin
            cosine_reg0 <= 36'sb10000110100010111010110101100110100;
            sine_reg0   <= 36'sb100100110001101010010110100010101110;
        end
        13732: begin
            cosine_reg0 <= 36'sb10000110101000010000111001111000000;
            sine_reg0   <= 36'sb100100110010000100110001110100010100;
        end
        13733: begin
            cosine_reg0 <= 36'sb10000110101101100110111000111101011;
            sine_reg0   <= 36'sb100100110010011111001110001001000011;
        end
        13734: begin
            cosine_reg0 <= 36'sb10000110110010111100110010110110011;
            sine_reg0   <= 36'sb100100110010111001101011100000111100;
        end
        13735: begin
            cosine_reg0 <= 36'sb10000110111000010010100111100010110;
            sine_reg0   <= 36'sb100100110011010100001001111011111100;
        end
        13736: begin
            cosine_reg0 <= 36'sb10000110111101101000010111000010010;
            sine_reg0   <= 36'sb100100110011101110101001011010000100;
        end
        13737: begin
            cosine_reg0 <= 36'sb10000111000010111110000001010100111;
            sine_reg0   <= 36'sb100100110100001001001001111011010010;
        end
        13738: begin
            cosine_reg0 <= 36'sb10000111001000010011100110011010010;
            sine_reg0   <= 36'sb100100110100100011101011011111100100;
        end
        13739: begin
            cosine_reg0 <= 36'sb10000111001101101001000110010010001;
            sine_reg0   <= 36'sb100100110100111110001110000110111010;
        end
        13740: begin
            cosine_reg0 <= 36'sb10000111010010111110100000111100011;
            sine_reg0   <= 36'sb100100110101011000110001110001010100;
        end
        13741: begin
            cosine_reg0 <= 36'sb10000111011000010011110110011000111;
            sine_reg0   <= 36'sb100100110101110011010110011110101111;
        end
        13742: begin
            cosine_reg0 <= 36'sb10000111011101101001000110100111011;
            sine_reg0   <= 36'sb100100110110001101111100001111001011;
        end
        13743: begin
            cosine_reg0 <= 36'sb10000111100010111110010001100111100;
            sine_reg0   <= 36'sb100100110110101000100011000010100110;
        end
        13744: begin
            cosine_reg0 <= 36'sb10000111101000010011010111011001010;
            sine_reg0   <= 36'sb100100110111000011001010111001000001;
        end
        13745: begin
            cosine_reg0 <= 36'sb10000111101101101000010111111100011;
            sine_reg0   <= 36'sb100100110111011101110011110010011001;
        end
        13746: begin
            cosine_reg0 <= 36'sb10000111110010111101010011010000101;
            sine_reg0   <= 36'sb100100110111111000011101101110101110;
        end
        13747: begin
            cosine_reg0 <= 36'sb10000111111000010010001001010101110;
            sine_reg0   <= 36'sb100100111000010011001000101101111111;
        end
        13748: begin
            cosine_reg0 <= 36'sb10000111111101100110111010001011101;
            sine_reg0   <= 36'sb100100111000101101110100110000001010;
        end
        13749: begin
            cosine_reg0 <= 36'sb10001000000010111011100101110010001;
            sine_reg0   <= 36'sb100100111001001000100001110101001111;
        end
        13750: begin
            cosine_reg0 <= 36'sb10001000001000010000001100001000111;
            sine_reg0   <= 36'sb100100111001100011001111111101001101;
        end
        13751: begin
            cosine_reg0 <= 36'sb10001000001101100100101101001111101;
            sine_reg0   <= 36'sb100100111001111101111111001000000010;
        end
        13752: begin
            cosine_reg0 <= 36'sb10001000010010111001001001000110100;
            sine_reg0   <= 36'sb100100111010011000101111010101101110;
        end
        13753: begin
            cosine_reg0 <= 36'sb10001000011000001101011111101100111;
            sine_reg0   <= 36'sb100100111010110011100000100110001111;
        end
        13754: begin
            cosine_reg0 <= 36'sb10001000011101100001110001000010111;
            sine_reg0   <= 36'sb100100111011001110010010111001100101;
        end
        13755: begin
            cosine_reg0 <= 36'sb10001000100010110101111101001000001;
            sine_reg0   <= 36'sb100100111011101001000110001111101110;
        end
        13756: begin
            cosine_reg0 <= 36'sb10001000101000001010000011111100100;
            sine_reg0   <= 36'sb100100111100000011111010101000101010;
        end
        13757: begin
            cosine_reg0 <= 36'sb10001000101101011110000101011111110;
            sine_reg0   <= 36'sb100100111100011110110000000100010111;
        end
        13758: begin
            cosine_reg0 <= 36'sb10001000110010110010000001110001110;
            sine_reg0   <= 36'sb100100111100111001100110100010110100;
        end
        13759: begin
            cosine_reg0 <= 36'sb10001000111000000101111000110010001;
            sine_reg0   <= 36'sb100100111101010100011110000100000001;
        end
        13760: begin
            cosine_reg0 <= 36'sb10001000111101011001101010100000110;
            sine_reg0   <= 36'sb100100111101101111010110100111111100;
        end
        13761: begin
            cosine_reg0 <= 36'sb10001001000010101101010110111101100;
            sine_reg0   <= 36'sb100100111110001010010000001110100100;
        end
        13762: begin
            cosine_reg0 <= 36'sb10001001001000000000111110001000001;
            sine_reg0   <= 36'sb100100111110100101001010110111111000;
        end
        13763: begin
            cosine_reg0 <= 36'sb10001001001101010100100000000000011;
            sine_reg0   <= 36'sb100100111111000000000110100011111000;
        end
        13764: begin
            cosine_reg0 <= 36'sb10001001010010100111111100100110001;
            sine_reg0   <= 36'sb100100111111011011000011010010100010;
        end
        13765: begin
            cosine_reg0 <= 36'sb10001001010111111011010011111001000;
            sine_reg0   <= 36'sb100100111111110110000001000011110100;
        end
        13766: begin
            cosine_reg0 <= 36'sb10001001011101001110100101111001000;
            sine_reg0   <= 36'sb100101000000010000111111110111101111;
        end
        13767: begin
            cosine_reg0 <= 36'sb10001001100010100001110010100101111;
            sine_reg0   <= 36'sb100101000000101011111111101110010001;
        end
        13768: begin
            cosine_reg0 <= 36'sb10001001100111110100111001111111011;
            sine_reg0   <= 36'sb100101000001000111000000100111011001;
        end
        13769: begin
            cosine_reg0 <= 36'sb10001001101101000111111100000101010;
            sine_reg0   <= 36'sb100101000001100010000010100011000110;
        end
        13770: begin
            cosine_reg0 <= 36'sb10001001110010011010111000110111011;
            sine_reg0   <= 36'sb100101000001111101000101100001010110;
        end
        13771: begin
            cosine_reg0 <= 36'sb10001001110111101101110000010101101;
            sine_reg0   <= 36'sb100101000010011000001001100010001010;
        end
        13772: begin
            cosine_reg0 <= 36'sb10001001111101000000100010011111100;
            sine_reg0   <= 36'sb100101000010110011001110100101011111;
        end
        13773: begin
            cosine_reg0 <= 36'sb10001010000010010011001111010101001;
            sine_reg0   <= 36'sb100101000011001110010100101011010101;
        end
        13774: begin
            cosine_reg0 <= 36'sb10001010000111100101110110110110001;
            sine_reg0   <= 36'sb100101000011101001011011110011101011;
        end
        13775: begin
            cosine_reg0 <= 36'sb10001010001100111000011001000010011;
            sine_reg0   <= 36'sb100101000100000100100011111110100000;
        end
        13776: begin
            cosine_reg0 <= 36'sb10001010010010001010110101111001100;
            sine_reg0   <= 36'sb100101000100011111101101001011110010;
        end
        13777: begin
            cosine_reg0 <= 36'sb10001010010111011101001101011011100;
            sine_reg0   <= 36'sb100101000100111010110111011011100000;
        end
        13778: begin
            cosine_reg0 <= 36'sb10001010011100101111011111101000001;
            sine_reg0   <= 36'sb100101000101010110000010101101101011;
        end
        13779: begin
            cosine_reg0 <= 36'sb10001010100010000001101100011111001;
            sine_reg0   <= 36'sb100101000101110001001111000010001111;
        end
        13780: begin
            cosine_reg0 <= 36'sb10001010100111010011110100000000010;
            sine_reg0   <= 36'sb100101000110001100011100011001001110;
        end
        13781: begin
            cosine_reg0 <= 36'sb10001010101100100101110110001011100;
            sine_reg0   <= 36'sb100101000110100111101010110010100100;
        end
        13782: begin
            cosine_reg0 <= 36'sb10001010110001110111110011000000011;
            sine_reg0   <= 36'sb100101000111000010111010001110010010;
        end
        13783: begin
            cosine_reg0 <= 36'sb10001010110111001001101010011110111;
            sine_reg0   <= 36'sb100101000111011110001010101100010110;
        end
        13784: begin
            cosine_reg0 <= 36'sb10001010111100011011011100100110110;
            sine_reg0   <= 36'sb100101000111111001011100001100101111;
        end
        13785: begin
            cosine_reg0 <= 36'sb10001011000001101101001001010111111;
            sine_reg0   <= 36'sb100101001000010100101110101111011101;
        end
        13786: begin
            cosine_reg0 <= 36'sb10001011000110111110110000110001111;
            sine_reg0   <= 36'sb100101001000110000000010010100011110;
        end
        13787: begin
            cosine_reg0 <= 36'sb10001011001100010000010010110100101;
            sine_reg0   <= 36'sb100101001001001011010110111011110000;
        end
        13788: begin
            cosine_reg0 <= 36'sb10001011010001100001101111100000000;
            sine_reg0   <= 36'sb100101001001100110101100100101010100;
        end
        13789: begin
            cosine_reg0 <= 36'sb10001011010110110011000110110011110;
            sine_reg0   <= 36'sb100101001010000010000011010001001000;
        end
        13790: begin
            cosine_reg0 <= 36'sb10001011011100000100011000101111100;
            sine_reg0   <= 36'sb100101001010011101011010111111001011;
        end
        13791: begin
            cosine_reg0 <= 36'sb10001011100001010101100101010011011;
            sine_reg0   <= 36'sb100101001010111000110011101111011011;
        end
        13792: begin
            cosine_reg0 <= 36'sb10001011100110100110101100011110111;
            sine_reg0   <= 36'sb100101001011010100001101100001111000;
        end
        13793: begin
            cosine_reg0 <= 36'sb10001011101011110111101110010010000;
            sine_reg0   <= 36'sb100101001011101111101000010110100001;
        end
        13794: begin
            cosine_reg0 <= 36'sb10001011110001001000101010101100011;
            sine_reg0   <= 36'sb100101001100001011000100001101010101;
        end
        13795: begin
            cosine_reg0 <= 36'sb10001011110110011001100001101110000;
            sine_reg0   <= 36'sb100101001100100110100001000110010011;
        end
        13796: begin
            cosine_reg0 <= 36'sb10001011111011101010010011010110100;
            sine_reg0   <= 36'sb100101001101000001111111000001011001;
        end
        13797: begin
            cosine_reg0 <= 36'sb10001100000000111010111111100101110;
            sine_reg0   <= 36'sb100101001101011101011101111110100110;
        end
        13798: begin
            cosine_reg0 <= 36'sb10001100000110001011100110011011100;
            sine_reg0   <= 36'sb100101001101111000111101111101111010;
        end
        13799: begin
            cosine_reg0 <= 36'sb10001100001011011100000111110111100;
            sine_reg0   <= 36'sb100101001110010100011110111111010011;
        end
        13800: begin
            cosine_reg0 <= 36'sb10001100010000101100100011111001110;
            sine_reg0   <= 36'sb100101001110110000000001000010110001;
        end
        13801: begin
            cosine_reg0 <= 36'sb10001100010101111100111010100001111;
            sine_reg0   <= 36'sb100101001111001011100100001000010010;
        end
        13802: begin
            cosine_reg0 <= 36'sb10001100011011001101001011101111110;
            sine_reg0   <= 36'sb100101001111100111001000001111110101;
        end
        13803: begin
            cosine_reg0 <= 36'sb10001100100000011101010111100011001;
            sine_reg0   <= 36'sb100101010000000010101101011001011010;
        end
        13804: begin
            cosine_reg0 <= 36'sb10001100100101101101011101111011110;
            sine_reg0   <= 36'sb100101010000011110010011100100111110;
        end
        13805: begin
            cosine_reg0 <= 36'sb10001100101010111101011110111001100;
            sine_reg0   <= 36'sb100101010000111001111010110010100001;
        end
        13806: begin
            cosine_reg0 <= 36'sb10001100110000001101011010011100010;
            sine_reg0   <= 36'sb100101010001010101100011000010000011;
        end
        13807: begin
            cosine_reg0 <= 36'sb10001100110101011101010000100011101;
            sine_reg0   <= 36'sb100101010001110001001100010011100001;
        end
        13808: begin
            cosine_reg0 <= 36'sb10001100111010101101000001001111100;
            sine_reg0   <= 36'sb100101010010001100110110100110111011;
        end
        13809: begin
            cosine_reg0 <= 36'sb10001100111111111100101100011111110;
            sine_reg0   <= 36'sb100101010010101000100001111100010000;
        end
        13810: begin
            cosine_reg0 <= 36'sb10001101000101001100010010010100000;
            sine_reg0   <= 36'sb100101010011000100001110010011011111;
        end
        13811: begin
            cosine_reg0 <= 36'sb10001101001010011011110010101100010;
            sine_reg0   <= 36'sb100101010011011111111011101100100110;
        end
        13812: begin
            cosine_reg0 <= 36'sb10001101001111101011001101101000001;
            sine_reg0   <= 36'sb100101010011111011101010000111100100;
        end
        13813: begin
            cosine_reg0 <= 36'sb10001101010100111010100011000111100;
            sine_reg0   <= 36'sb100101010100010111011001100100011010;
        end
        13814: begin
            cosine_reg0 <= 36'sb10001101011010001001110011001010001;
            sine_reg0   <= 36'sb100101010100110011001010000011000100;
        end
        13815: begin
            cosine_reg0 <= 36'sb10001101011111011000111101101111111;
            sine_reg0   <= 36'sb100101010101001110111011100011100011;
        end
        13816: begin
            cosine_reg0 <= 36'sb10001101100100101000000010111000100;
            sine_reg0   <= 36'sb100101010101101010101110000101110110;
        end
        13817: begin
            cosine_reg0 <= 36'sb10001101101001110111000010100011111;
            sine_reg0   <= 36'sb100101010110000110100001101001111010;
        end
        13818: begin
            cosine_reg0 <= 36'sb10001101101111000101111100110001101;
            sine_reg0   <= 36'sb100101010110100010010110001111110000;
        end
        13819: begin
            cosine_reg0 <= 36'sb10001101110100010100110001100001110;
            sine_reg0   <= 36'sb100101010110111110001011110111010101;
        end
        13820: begin
            cosine_reg0 <= 36'sb10001101111001100011100000110100000;
            sine_reg0   <= 36'sb100101010111011010000010100000101010;
        end
        13821: begin
            cosine_reg0 <= 36'sb10001101111110110010001010101000000;
            sine_reg0   <= 36'sb100101010111110101111010001011101101;
        end
        13822: begin
            cosine_reg0 <= 36'sb10001110000100000000101110111101110;
            sine_reg0   <= 36'sb100101011000010001110010111000011100;
        end
        13823: begin
            cosine_reg0 <= 36'sb10001110001001001111001101110100111;
            sine_reg0   <= 36'sb100101011000101101101100100110110111;
        end
        13824: begin
            cosine_reg0 <= 36'sb10001110001110011101100111001101011;
            sine_reg0   <= 36'sb100101011001001001100111010110111101;
        end
        13825: begin
            cosine_reg0 <= 36'sb10001110010011101011111011000110111;
            sine_reg0   <= 36'sb100101011001100101100011001000101101;
        end
        13826: begin
            cosine_reg0 <= 36'sb10001110011000111010001001100001011;
            sine_reg0   <= 36'sb100101011010000001011111111100000101;
        end
        13827: begin
            cosine_reg0 <= 36'sb10001110011110001000010010011100011;
            sine_reg0   <= 36'sb100101011010011101011101110001000100;
        end
        13828: begin
            cosine_reg0 <= 36'sb10001110100011010110010101111000000;
            sine_reg0   <= 36'sb100101011010111001011100100111101010;
        end
        13829: begin
            cosine_reg0 <= 36'sb10001110101000100100010011110011110;
            sine_reg0   <= 36'sb100101011011010101011100011111110101;
        end
        13830: begin
            cosine_reg0 <= 36'sb10001110101101110010001100001111101;
            sine_reg0   <= 36'sb100101011011110001011101011001100101;
        end
        13831: begin
            cosine_reg0 <= 36'sb10001110110010111111111111001011011;
            sine_reg0   <= 36'sb100101011100001101011111010100110111;
        end
        13832: begin
            cosine_reg0 <= 36'sb10001110111000001101101100100110111;
            sine_reg0   <= 36'sb100101011100101001100010010001101100;
        end
        13833: begin
            cosine_reg0 <= 36'sb10001110111101011011010100100001101;
            sine_reg0   <= 36'sb100101011101000101100110010000000001;
        end
        13834: begin
            cosine_reg0 <= 36'sb10001111000010101000110110111011111;
            sine_reg0   <= 36'sb100101011101100001101011001111110111;
        end
        13835: begin
            cosine_reg0 <= 36'sb10001111000111110110010011110101000;
            sine_reg0   <= 36'sb100101011101111101110001010001001011;
        end
        13836: begin
            cosine_reg0 <= 36'sb10001111001101000011101011001101000;
            sine_reg0   <= 36'sb100101011110011001111000010011111101;
        end
        13837: begin
            cosine_reg0 <= 36'sb10001111010010010000111101000011110;
            sine_reg0   <= 36'sb100101011110110110000000011000001100;
        end
        13838: begin
            cosine_reg0 <= 36'sb10001111010111011110001001011000111;
            sine_reg0   <= 36'sb100101011111010010001001011101110110;
        end
        13839: begin
            cosine_reg0 <= 36'sb10001111011100101011010000001100011;
            sine_reg0   <= 36'sb100101011111101110010011100100111011;
        end
        13840: begin
            cosine_reg0 <= 36'sb10001111100001111000010001011101111;
            sine_reg0   <= 36'sb100101100000001010011110101101011001;
        end
        13841: begin
            cosine_reg0 <= 36'sb10001111100111000101001101001101001;
            sine_reg0   <= 36'sb100101100000100110101010110111001111;
        end
        13842: begin
            cosine_reg0 <= 36'sb10001111101100010010000011011010001;
            sine_reg0   <= 36'sb100101100001000010111000000010011101;
        end
        13843: begin
            cosine_reg0 <= 36'sb10001111110001011110110100000100101;
            sine_reg0   <= 36'sb100101100001011111000110001111000001;
        end
        13844: begin
            cosine_reg0 <= 36'sb10001111110110101011011111001100010;
            sine_reg0   <= 36'sb100101100001111011010101011100111010;
        end
        13845: begin
            cosine_reg0 <= 36'sb10001111111011111000000100110001000;
            sine_reg0   <= 36'sb100101100010010111100101101100000110;
        end
        13846: begin
            cosine_reg0 <= 36'sb10010000000001000100100100110010101;
            sine_reg0   <= 36'sb100101100010110011110110111100100110;
        end
        13847: begin
            cosine_reg0 <= 36'sb10010000000110010000111111010000111;
            sine_reg0   <= 36'sb100101100011010000001001001110010111;
        end
        13848: begin
            cosine_reg0 <= 36'sb10010000001011011101010100001011101;
            sine_reg0   <= 36'sb100101100011101100011100100001011001;
        end
        13849: begin
            cosine_reg0 <= 36'sb10010000010000101001100011100010100;
            sine_reg0   <= 36'sb100101100100001000110000110101101011;
        end
        13850: begin
            cosine_reg0 <= 36'sb10010000010101110101101101010101101;
            sine_reg0   <= 36'sb100101100100100101000110001011001011;
        end
        13851: begin
            cosine_reg0 <= 36'sb10010000011011000001110001100100100;
            sine_reg0   <= 36'sb100101100101000001011100100001111001;
        end
        13852: begin
            cosine_reg0 <= 36'sb10010000100000001101110000001111000;
            sine_reg0   <= 36'sb100101100101011101110011111001110011;
        end
        13853: begin
            cosine_reg0 <= 36'sb10010000100101011001101001010100111;
            sine_reg0   <= 36'sb100101100101111010001100010010111000;
        end
        13854: begin
            cosine_reg0 <= 36'sb10010000101010100101011100110110001;
            sine_reg0   <= 36'sb100101100110010110100101101101000111;
        end
        13855: begin
            cosine_reg0 <= 36'sb10010000101111110001001010110010011;
            sine_reg0   <= 36'sb100101100110110011000000001000100000;
        end
        13856: begin
            cosine_reg0 <= 36'sb10010000110100111100110011001001100;
            sine_reg0   <= 36'sb100101100111001111011011100101000000;
        end
        13857: begin
            cosine_reg0 <= 36'sb10010000111010001000010101111011011;
            sine_reg0   <= 36'sb100101100111101011111000000010100111;
        end
        13858: begin
            cosine_reg0 <= 36'sb10010000111111010011110011000111101;
            sine_reg0   <= 36'sb100101101000001000010101100001010100;
        end
        13859: begin
            cosine_reg0 <= 36'sb10010001000100011111001010101110000;
            sine_reg0   <= 36'sb100101101000100100110100000001000110;
        end
        13860: begin
            cosine_reg0 <= 36'sb10010001001001101010011100101110101;
            sine_reg0   <= 36'sb100101101001000001010011100001111011;
        end
        13861: begin
            cosine_reg0 <= 36'sb10010001001110110101101001001001000;
            sine_reg0   <= 36'sb100101101001011101110100000011110010;
        end
        13862: begin
            cosine_reg0 <= 36'sb10010001010100000000101111111101000;
            sine_reg0   <= 36'sb100101101001111010010101100110101011;
        end
        13863: begin
            cosine_reg0 <= 36'sb10010001011001001011110001001010100;
            sine_reg0   <= 36'sb100101101010010110111000001010100100;
        end
        13864: begin
            cosine_reg0 <= 36'sb10010001011110010110101100110001010;
            sine_reg0   <= 36'sb100101101010110011011011101111011101;
        end
        13865: begin
            cosine_reg0 <= 36'sb10010001100011100001100010110001001;
            sine_reg0   <= 36'sb100101101011010000000000010101010011;
        end
        13866: begin
            cosine_reg0 <= 36'sb10010001101000101100010011001001110;
            sine_reg0   <= 36'sb100101101011101100100101111100000110;
        end
        13867: begin
            cosine_reg0 <= 36'sb10010001101101110110111101111011001;
            sine_reg0   <= 36'sb100101101100001001001100100011110101;
        end
        13868: begin
            cosine_reg0 <= 36'sb10010001110011000001100011000100111;
            sine_reg0   <= 36'sb100101101100100101110100001100011111;
        end
        13869: begin
            cosine_reg0 <= 36'sb10010001111000001100000010100111000;
            sine_reg0   <= 36'sb100101101101000010011100110110000011;
        end
        13870: begin
            cosine_reg0 <= 36'sb10010001111101010110011100100001001;
            sine_reg0   <= 36'sb100101101101011111000110100000011111;
        end
        13871: begin
            cosine_reg0 <= 36'sb10010010000010100000110000110011001;
            sine_reg0   <= 36'sb100101101101111011110001001011110011;
        end
        13872: begin
            cosine_reg0 <= 36'sb10010010000111101010111111011100110;
            sine_reg0   <= 36'sb100101101110011000011100110111111100;
        end
        13873: begin
            cosine_reg0 <= 36'sb10010010001100110101001000011101110;
            sine_reg0   <= 36'sb100101101110110101001001100100111100;
        end
        13874: begin
            cosine_reg0 <= 36'sb10010010010001111111001011110110001;
            sine_reg0   <= 36'sb100101101111010001110111010010101111;
        end
        13875: begin
            cosine_reg0 <= 36'sb10010010010111001001001001100101101;
            sine_reg0   <= 36'sb100101101111101110100110000001010101;
        end
        13876: begin
            cosine_reg0 <= 36'sb10010010011100010011000001101011111;
            sine_reg0   <= 36'sb100101110000001011010101110000101101;
        end
        13877: begin
            cosine_reg0 <= 36'sb10010010100001011100110100001000111;
            sine_reg0   <= 36'sb100101110000101000000110100000110110;
        end
        13878: begin
            cosine_reg0 <= 36'sb10010010100110100110100000111100010;
            sine_reg0   <= 36'sb100101110001000100111000010001101111;
        end
        13879: begin
            cosine_reg0 <= 36'sb10010010101011110000001000000110000;
            sine_reg0   <= 36'sb100101110001100001101011000011010110;
        end
        13880: begin
            cosine_reg0 <= 36'sb10010010110000111001101001100101110;
            sine_reg0   <= 36'sb100101110001111110011110110101101011;
        end
        13881: begin
            cosine_reg0 <= 36'sb10010010110110000011000101011011100;
            sine_reg0   <= 36'sb100101110010011011010011101000101100;
        end
        13882: begin
            cosine_reg0 <= 36'sb10010010111011001100011011100110110;
            sine_reg0   <= 36'sb100101110010111000001001011100011000;
        end
        13883: begin
            cosine_reg0 <= 36'sb10010011000000010101101100000111101;
            sine_reg0   <= 36'sb100101110011010101000000010000101110;
        end
        13884: begin
            cosine_reg0 <= 36'sb10010011000101011110110110111101101;
            sine_reg0   <= 36'sb100101110011110001111000000101101110;
        end
        13885: begin
            cosine_reg0 <= 36'sb10010011001010100111111100001000111;
            sine_reg0   <= 36'sb100101110100001110110000111011010101;
        end
        13886: begin
            cosine_reg0 <= 36'sb10010011001111110000111011101000111;
            sine_reg0   <= 36'sb100101110100101011101010110001100011;
        end
        13887: begin
            cosine_reg0 <= 36'sb10010011010100111001110101011101101;
            sine_reg0   <= 36'sb100101110101001000100101101000010111;
        end
        13888: begin
            cosine_reg0 <= 36'sb10010011011010000010101001100110111;
            sine_reg0   <= 36'sb100101110101100101100001011111101111;
        end
        13889: begin
            cosine_reg0 <= 36'sb10010011011111001011011000000100011;
            sine_reg0   <= 36'sb100101110110000010011110010111101011;
        end
        13890: begin
            cosine_reg0 <= 36'sb10010011100100010100000000110110000;
            sine_reg0   <= 36'sb100101110110011111011100010000001001;
        end
        13891: begin
            cosine_reg0 <= 36'sb10010011101001011100100011111011011;
            sine_reg0   <= 36'sb100101110110111100011011001001001001;
        end
        13892: begin
            cosine_reg0 <= 36'sb10010011101110100101000001010100101;
            sine_reg0   <= 36'sb100101110111011001011011000010101000;
        end
        13893: begin
            cosine_reg0 <= 36'sb10010011110011101101011001000001010;
            sine_reg0   <= 36'sb100101110111110110011011111100100111;
        end
        13894: begin
            cosine_reg0 <= 36'sb10010011111000110101101011000001010;
            sine_reg0   <= 36'sb100101111000010011011101110111000011;
        end
        13895: begin
            cosine_reg0 <= 36'sb10010011111101111101110111010100011;
            sine_reg0   <= 36'sb100101111000110000100000110001111100;
        end
        13896: begin
            cosine_reg0 <= 36'sb10010100000011000101111101111010011;
            sine_reg0   <= 36'sb100101111001001101100100101101010001;
        end
        13897: begin
            cosine_reg0 <= 36'sb10010100001000001101111110110011000;
            sine_reg0   <= 36'sb100101111001101010101001101001000000;
        end
        13898: begin
            cosine_reg0 <= 36'sb10010100001101010101111001111110010;
            sine_reg0   <= 36'sb100101111010000111101111100101001000;
        end
        13899: begin
            cosine_reg0 <= 36'sb10010100010010011101101111011011110;
            sine_reg0   <= 36'sb100101111010100100110110100001101001;
        end
        13900: begin
            cosine_reg0 <= 36'sb10010100010111100101011111001011011;
            sine_reg0   <= 36'sb100101111011000001111110011110100001;
        end
        13901: begin
            cosine_reg0 <= 36'sb10010100011100101101001001001100111;
            sine_reg0   <= 36'sb100101111011011111000111011011101111;
        end
        13902: begin
            cosine_reg0 <= 36'sb10010100100001110100101101100000001;
            sine_reg0   <= 36'sb100101111011111100010001011001010010;
        end
        13903: begin
            cosine_reg0 <= 36'sb10010100100110111100001100000100111;
            sine_reg0   <= 36'sb100101111100011001011100010111001001;
        end
        13904: begin
            cosine_reg0 <= 36'sb10010100101100000011100100111011000;
            sine_reg0   <= 36'sb100101111100110110101000010101010010;
        end
        13905: begin
            cosine_reg0 <= 36'sb10010100110001001010111000000010010;
            sine_reg0   <= 36'sb100101111101010011110101010011101101;
        end
        13906: begin
            cosine_reg0 <= 36'sb10010100110110010010000101011010011;
            sine_reg0   <= 36'sb100101111101110001000011010010011000;
        end
        13907: begin
            cosine_reg0 <= 36'sb10010100111011011001001101000011010;
            sine_reg0   <= 36'sb100101111110001110010010010001010011;
        end
        13908: begin
            cosine_reg0 <= 36'sb10010101000000100000001110111100101;
            sine_reg0   <= 36'sb100101111110101011100010010000011011;
        end
        13909: begin
            cosine_reg0 <= 36'sb10010101000101100111001011000110100;
            sine_reg0   <= 36'sb100101111111001000110011001111110001;
        end
        13910: begin
            cosine_reg0 <= 36'sb10010101001010101110000001100000011;
            sine_reg0   <= 36'sb100101111111100110000101001111010010;
        end
        13911: begin
            cosine_reg0 <= 36'sb10010101001111110100110010001010001;
            sine_reg0   <= 36'sb100110000000000011011000001110111111;
        end
        13912: begin
            cosine_reg0 <= 36'sb10010101010100111011011101000011110;
            sine_reg0   <= 36'sb100110000000100000101100001110110100;
        end
        13913: begin
            cosine_reg0 <= 36'sb10010101011010000010000010001100111;
            sine_reg0   <= 36'sb100110000000111110000001001110110011;
        end
        13914: begin
            cosine_reg0 <= 36'sb10010101011111001000100001100101011;
            sine_reg0   <= 36'sb100110000001011011010111001110111001;
        end
        13915: begin
            cosine_reg0 <= 36'sb10010101100100001110111011001101000;
            sine_reg0   <= 36'sb100110000001111000101110001111000101;
        end
        13916: begin
            cosine_reg0 <= 36'sb10010101101001010101001111000011101;
            sine_reg0   <= 36'sb100110000010010110000110001111010110;
        end
        13917: begin
            cosine_reg0 <= 36'sb10010101101110011011011101001001000;
            sine_reg0   <= 36'sb100110000010110011011111001111101011;
        end
        13918: begin
            cosine_reg0 <= 36'sb10010101110011100001100101011101000;
            sine_reg0   <= 36'sb100110000011010000111001010000000011;
        end
        13919: begin
            cosine_reg0 <= 36'sb10010101111000100111100111111111010;
            sine_reg0   <= 36'sb100110000011101110010100010000011100;
        end
        13920: begin
            cosine_reg0 <= 36'sb10010101111101101101100100101111110;
            sine_reg0   <= 36'sb100110000100001011110000010000110110;
        end
        13921: begin
            cosine_reg0 <= 36'sb10010110000010110011011011101110010;
            sine_reg0   <= 36'sb100110000100101001001101010001010000;
        end
        13922: begin
            cosine_reg0 <= 36'sb10010110000111111001001100111010100;
            sine_reg0   <= 36'sb100110000101000110101011010001101000;
        end
        13923: begin
            cosine_reg0 <= 36'sb10010110001100111110111000010100010;
            sine_reg0   <= 36'sb100110000101100100001010010001111101;
        end
        13924: begin
            cosine_reg0 <= 36'sb10010110010010000100011101111011100;
            sine_reg0   <= 36'sb100110000110000001101010010010001110;
        end
        13925: begin
            cosine_reg0 <= 36'sb10010110010111001001111101110000000;
            sine_reg0   <= 36'sb100110000110011111001011010010011010;
        end
        13926: begin
            cosine_reg0 <= 36'sb10010110011100001111010111110001011;
            sine_reg0   <= 36'sb100110000110111100101101010010100000;
        end
        13927: begin
            cosine_reg0 <= 36'sb10010110100001010100101011111111101;
            sine_reg0   <= 36'sb100110000111011010010000010010011110;
        end
        13928: begin
            cosine_reg0 <= 36'sb10010110100110011001111010011010011;
            sine_reg0   <= 36'sb100110000111110111110100010010010100;
        end
        13929: begin
            cosine_reg0 <= 36'sb10010110101011011111000011000001101;
            sine_reg0   <= 36'sb100110001000010101011001010010000000;
        end
        13930: begin
            cosine_reg0 <= 36'sb10010110110000100100000101110101000;
            sine_reg0   <= 36'sb100110001000110010111111010001100001;
        end
        13931: begin
            cosine_reg0 <= 36'sb10010110110101101001000010110100100;
            sine_reg0   <= 36'sb100110001001010000100110010000110111;
        end
        13932: begin
            cosine_reg0 <= 36'sb10010110111010101101111001111111110;
            sine_reg0   <= 36'sb100110001001101110001110001111111111;
        end
        13933: begin
            cosine_reg0 <= 36'sb10010110111111110010101011010110110;
            sine_reg0   <= 36'sb100110001010001011110111001110111001;
        end
        13934: begin
            cosine_reg0 <= 36'sb10010111000100110111010110111001000;
            sine_reg0   <= 36'sb100110001010101001100001001101100100;
        end
        13935: begin
            cosine_reg0 <= 36'sb10010111001001111011111100100110101;
            sine_reg0   <= 36'sb100110001011000111001100001011111110;
        end
        13936: begin
            cosine_reg0 <= 36'sb10010111001111000000011100011111010;
            sine_reg0   <= 36'sb100110001011100100111000001010000110;
        end
        13937: begin
            cosine_reg0 <= 36'sb10010111010100000100110110100010101;
            sine_reg0   <= 36'sb100110001100000010100101000111111100;
        end
        13938: begin
            cosine_reg0 <= 36'sb10010111011001001001001010110000110;
            sine_reg0   <= 36'sb100110001100100000010011000101011110;
        end
        13939: begin
            cosine_reg0 <= 36'sb10010111011110001101011001001001011;
            sine_reg0   <= 36'sb100110001100111110000010000010101010;
        end
        13940: begin
            cosine_reg0 <= 36'sb10010111100011010001100001101100001;
            sine_reg0   <= 36'sb100110001101011011110001111111100001;
        end
        13941: begin
            cosine_reg0 <= 36'sb10010111101000010101100100011001000;
            sine_reg0   <= 36'sb100110001101111001100010111100000000;
        end
        13942: begin
            cosine_reg0 <= 36'sb10010111101101011001100001001111110;
            sine_reg0   <= 36'sb100110001110010111010100111000000110;
        end
        13943: begin
            cosine_reg0 <= 36'sb10010111110010011101011000010000001;
            sine_reg0   <= 36'sb100110001110110101000111110011110011;
        end
        13944: begin
            cosine_reg0 <= 36'sb10010111110111100001001001011010000;
            sine_reg0   <= 36'sb100110001111010010111011101111000101;
        end
        13945: begin
            cosine_reg0 <= 36'sb10010111111100100100110100101101010;
            sine_reg0   <= 36'sb100110001111110000110000101001111011;
        end
        13946: begin
            cosine_reg0 <= 36'sb10011000000001101000011010001001100;
            sine_reg0   <= 36'sb100110010000001110100110100100010011;
        end
        13947: begin
            cosine_reg0 <= 36'sb10011000000110101011111001101110101;
            sine_reg0   <= 36'sb100110010000101100011101011110001110;
        end
        13948: begin
            cosine_reg0 <= 36'sb10011000001011101111010011011100100;
            sine_reg0   <= 36'sb100110010001001010010101010111101001;
        end
        13949: begin
            cosine_reg0 <= 36'sb10011000010000110010100111010010111;
            sine_reg0   <= 36'sb100110010001101000001110010000100100;
        end
        13950: begin
            cosine_reg0 <= 36'sb10011000010101110101110101010001100;
            sine_reg0   <= 36'sb100110010010000110001000001000111100;
        end
        13951: begin
            cosine_reg0 <= 36'sb10011000011010111000111101011000010;
            sine_reg0   <= 36'sb100110010010100100000011000000110010;
        end
        13952: begin
            cosine_reg0 <= 36'sb10011000011111111011111111100111000;
            sine_reg0   <= 36'sb100110010011000001111110111000000100;
        end
        13953: begin
            cosine_reg0 <= 36'sb10011000100100111110111011111101011;
            sine_reg0   <= 36'sb100110010011011111111011101110110001;
        end
        13954: begin
            cosine_reg0 <= 36'sb10011000101010000001110010011011011;
            sine_reg0   <= 36'sb100110010011111101111001100100110111;
        end
        13955: begin
            cosine_reg0 <= 36'sb10011000101111000100100011000000101;
            sine_reg0   <= 36'sb100110010100011011111000011010010110;
        end
        13956: begin
            cosine_reg0 <= 36'sb10011000110100000111001101101101000;
            sine_reg0   <= 36'sb100110010100111001111000001111001100;
        end
        13957: begin
            cosine_reg0 <= 36'sb10011000111001001001110010100000011;
            sine_reg0   <= 36'sb100110010101010111111001000011011000;
        end
        13958: begin
            cosine_reg0 <= 36'sb10011000111110001100010001011010100;
            sine_reg0   <= 36'sb100110010101110101111010110110111001;
        end
        13959: begin
            cosine_reg0 <= 36'sb10011001000011001110101010011011010;
            sine_reg0   <= 36'sb100110010110010011111101101001101110;
        end
        13960: begin
            cosine_reg0 <= 36'sb10011001001000010000111101100010010;
            sine_reg0   <= 36'sb100110010110110010000001011011110110;
        end
        13961: begin
            cosine_reg0 <= 36'sb10011001001101010011001010101111011;
            sine_reg0   <= 36'sb100110010111010000000110001101001111;
        end
        13962: begin
            cosine_reg0 <= 36'sb10011001010010010101010010000010101;
            sine_reg0   <= 36'sb100110010111101110001011111101111001;
        end
        13963: begin
            cosine_reg0 <= 36'sb10011001010111010111010011011011101;
            sine_reg0   <= 36'sb100110011000001100010010101101110010;
        end
        13964: begin
            cosine_reg0 <= 36'sb10011001011100011001001110111010001;
            sine_reg0   <= 36'sb100110011000101010011010011100111001;
        end
        13965: begin
            cosine_reg0 <= 36'sb10011001100001011011000100011110001;
            sine_reg0   <= 36'sb100110011001001000100011001011001101;
        end
        13966: begin
            cosine_reg0 <= 36'sb10011001100110011100110100000111010;
            sine_reg0   <= 36'sb100110011001100110101100111000101101;
        end
        13967: begin
            cosine_reg0 <= 36'sb10011001101011011110011101110101011;
            sine_reg0   <= 36'sb100110011010000100110111100101010111;
        end
        13968: begin
            cosine_reg0 <= 36'sb10011001110000100000000001101000011;
            sine_reg0   <= 36'sb100110011010100011000011010001001011;
        end
        13969: begin
            cosine_reg0 <= 36'sb10011001110101100001011111011111111;
            sine_reg0   <= 36'sb100110011011000001001111111100000111;
        end
        13970: begin
            cosine_reg0 <= 36'sb10011001111010100010110111011011111;
            sine_reg0   <= 36'sb100110011011011111011101100110001010;
        end
        13971: begin
            cosine_reg0 <= 36'sb10011001111111100100001001011100001;
            sine_reg0   <= 36'sb100110011011111101101100001111010011;
        end
        13972: begin
            cosine_reg0 <= 36'sb10011010000100100101010101100000011;
            sine_reg0   <= 36'sb100110011100011011111011110111100000;
        end
        13973: begin
            cosine_reg0 <= 36'sb10011010001001100110011011101000100;
            sine_reg0   <= 36'sb100110011100111010001100011110110010;
        end
        13974: begin
            cosine_reg0 <= 36'sb10011010001110100111011011110100010;
            sine_reg0   <= 36'sb100110011101011000011110000101000101;
        end
        13975: begin
            cosine_reg0 <= 36'sb10011010010011101000010110000011100;
            sine_reg0   <= 36'sb100110011101110110110000101010011010;
        end
        13976: begin
            cosine_reg0 <= 36'sb10011010011000101001001010010110000;
            sine_reg0   <= 36'sb100110011110010101000100001110101111;
        end
        13977: begin
            cosine_reg0 <= 36'sb10011010011101101001111000101011100;
            sine_reg0   <= 36'sb100110011110110011011000110010000011;
        end
        13978: begin
            cosine_reg0 <= 36'sb10011010100010101010100001000100000;
            sine_reg0   <= 36'sb100110011111010001101110010100010101;
        end
        13979: begin
            cosine_reg0 <= 36'sb10011010100111101011000011011111000;
            sine_reg0   <= 36'sb100110011111110000000100110101100011;
        end
        13980: begin
            cosine_reg0 <= 36'sb10011010101100101011011111111100101;
            sine_reg0   <= 36'sb100110100000001110011100010101101101;
        end
        13981: begin
            cosine_reg0 <= 36'sb10011010110001101011110110011100101;
            sine_reg0   <= 36'sb100110100000101100110100110100110001;
        end
        13982: begin
            cosine_reg0 <= 36'sb10011010110110101100000110111110101;
            sine_reg0   <= 36'sb100110100001001011001110010010101110;
        end
        13983: begin
            cosine_reg0 <= 36'sb10011010111011101100010001100010100;
            sine_reg0   <= 36'sb100110100001101001101000101111100011;
        end
        13984: begin
            cosine_reg0 <= 36'sb10011011000000101100010110001000001;
            sine_reg0   <= 36'sb100110100010001000000100001011001111;
        end
        13985: begin
            cosine_reg0 <= 36'sb10011011000101101100010100101111010;
            sine_reg0   <= 36'sb100110100010100110100000100101110000;
        end
        13986: begin
            cosine_reg0 <= 36'sb10011011001010101100001101010111110;
            sine_reg0   <= 36'sb100110100011000100111101111111000110;
        end
        13987: begin
            cosine_reg0 <= 36'sb10011011001111101100000000000001011;
            sine_reg0   <= 36'sb100110100011100011011100010111001110;
        end
        13988: begin
            cosine_reg0 <= 36'sb10011011010100101011101100101100000;
            sine_reg0   <= 36'sb100110100100000001111011101110001001;
        end
        13989: begin
            cosine_reg0 <= 36'sb10011011011001101011010011010111011;
            sine_reg0   <= 36'sb100110100100100000011100000011110101;
        end
        13990: begin
            cosine_reg0 <= 36'sb10011011011110101010110100000011010;
            sine_reg0   <= 36'sb100110100100111110111101011000010000;
        end
        13991: begin
            cosine_reg0 <= 36'sb10011011100011101010001110101111100;
            sine_reg0   <= 36'sb100110100101011101011111101011011010;
        end
        13992: begin
            cosine_reg0 <= 36'sb10011011101000101001100011011100000;
            sine_reg0   <= 36'sb100110100101111100000010111101010001;
        end
        13993: begin
            cosine_reg0 <= 36'sb10011011101101101000110010001000011;
            sine_reg0   <= 36'sb100110100110011010100111001101110101;
        end
        13994: begin
            cosine_reg0 <= 36'sb10011011110010100111111010110100101;
            sine_reg0   <= 36'sb100110100110111001001100011101000011;
        end
        13995: begin
            cosine_reg0 <= 36'sb10011011110111100110111101100000100;
            sine_reg0   <= 36'sb100110100111010111110010101010111011;
        end
        13996: begin
            cosine_reg0 <= 36'sb10011011111100100101111010001011110;
            sine_reg0   <= 36'sb100110100111110110011001110111011100;
        end
        13997: begin
            cosine_reg0 <= 36'sb10011100000001100100110000110110001;
            sine_reg0   <= 36'sb100110101000010101000010000010100100;
        end
        13998: begin
            cosine_reg0 <= 36'sb10011100000110100011100001011111101;
            sine_reg0   <= 36'sb100110101000110011101011001100010010;
        end
        13999: begin
            cosine_reg0 <= 36'sb10011100001011100010001100001000000;
            sine_reg0   <= 36'sb100110101001010010010101010100100110;
        end
        14000: begin
            cosine_reg0 <= 36'sb10011100010000100000110000101110111;
            sine_reg0   <= 36'sb100110101001110001000000011011011101;
        end
        14001: begin
            cosine_reg0 <= 36'sb10011100010101011111001111010100011;
            sine_reg0   <= 36'sb100110101010001111101100100000110111;
        end
        14002: begin
            cosine_reg0 <= 36'sb10011100011010011101100111111000000;
            sine_reg0   <= 36'sb100110101010101110011001100100110011;
        end
        14003: begin
            cosine_reg0 <= 36'sb10011100011111011011111010011001110;
            sine_reg0   <= 36'sb100110101011001101000111100111001111;
        end
        14004: begin
            cosine_reg0 <= 36'sb10011100100100011010000110111001011;
            sine_reg0   <= 36'sb100110101011101011110110101000001010;
        end
        14005: begin
            cosine_reg0 <= 36'sb10011100101001011000001101010110101;
            sine_reg0   <= 36'sb100110101100001010100110100111100011;
        end
        14006: begin
            cosine_reg0 <= 36'sb10011100101110010110001101110001011;
            sine_reg0   <= 36'sb100110101100101001010111100101011001;
        end
        14007: begin
            cosine_reg0 <= 36'sb10011100110011010100001000001001100;
            sine_reg0   <= 36'sb100110101101001000001001100001101010;
        end
        14008: begin
            cosine_reg0 <= 36'sb10011100111000010001111100011110101;
            sine_reg0   <= 36'sb100110101101100110111100011100010110;
        end
        14009: begin
            cosine_reg0 <= 36'sb10011100111101001111101010110000110;
            sine_reg0   <= 36'sb100110101110000101110000010101011011;
        end
        14010: begin
            cosine_reg0 <= 36'sb10011101000010001101010010111111100;
            sine_reg0   <= 36'sb100110101110100100100101001100111000;
        end
        14011: begin
            cosine_reg0 <= 36'sb10011101000111001010110101001010111;
            sine_reg0   <= 36'sb100110101111000011011011000010101100;
        end
        14012: begin
            cosine_reg0 <= 36'sb10011101001100001000010001010010101;
            sine_reg0   <= 36'sb100110101111100010010001110110110101;
        end
        14013: begin
            cosine_reg0 <= 36'sb10011101010001000101100111010110011;
            sine_reg0   <= 36'sb100110110000000001001001101001010011;
        end
        14014: begin
            cosine_reg0 <= 36'sb10011101010110000010110111010110010;
            sine_reg0   <= 36'sb100110110000100000000010011010000101;
        end
        14015: begin
            cosine_reg0 <= 36'sb10011101011011000000000001010001110;
            sine_reg0   <= 36'sb100110110000111110111100001001001000;
        end
        14016: begin
            cosine_reg0 <= 36'sb10011101011111111101000101001000111;
            sine_reg0   <= 36'sb100110110001011101110110110110011100;
        end
        14017: begin
            cosine_reg0 <= 36'sb10011101100100111010000010111011100;
            sine_reg0   <= 36'sb100110110001111100110010100010000000;
        end
        14018: begin
            cosine_reg0 <= 36'sb10011101101001110110111010101001010;
            sine_reg0   <= 36'sb100110110010011011101111001011110011;
        end
        14019: begin
            cosine_reg0 <= 36'sb10011101101110110011101100010001111;
            sine_reg0   <= 36'sb100110110010111010101100110011110010;
        end
        14020: begin
            cosine_reg0 <= 36'sb10011101110011110000010111110101100;
            sine_reg0   <= 36'sb100110110011011001101011011001111110;
        end
        14021: begin
            cosine_reg0 <= 36'sb10011101111000101100111101010011101;
            sine_reg0   <= 36'sb100110110011111000101010111110010101;
        end
        14022: begin
            cosine_reg0 <= 36'sb10011101111101101001011100101100010;
            sine_reg0   <= 36'sb100110110100010111101011100000110110;
        end
        14023: begin
            cosine_reg0 <= 36'sb10011110000010100101110101111111001;
            sine_reg0   <= 36'sb100110110100110110101101000001011111;
        end
        14024: begin
            cosine_reg0 <= 36'sb10011110000111100010001001001100000;
            sine_reg0   <= 36'sb100110110101010101101111100000001111;
        end
        14025: begin
            cosine_reg0 <= 36'sb10011110001100011110010110010010110;
            sine_reg0   <= 36'sb100110110101110100110010111101000110;
        end
        14026: begin
            cosine_reg0 <= 36'sb10011110010001011010011101010011001;
            sine_reg0   <= 36'sb100110110110010011110111011000000010;
        end
        14027: begin
            cosine_reg0 <= 36'sb10011110010110010110011110001101000;
            sine_reg0   <= 36'sb100110110110110010111100110001000001;
        end
        14028: begin
            cosine_reg0 <= 36'sb10011110011011010010011001000000010;
            sine_reg0   <= 36'sb100110110111010010000011001000000011;
        end
        14029: begin
            cosine_reg0 <= 36'sb10011110100000001110001101101100100;
            sine_reg0   <= 36'sb100110110111110001001010011101000110;
        end
        14030: begin
            cosine_reg0 <= 36'sb10011110100101001001111100010001110;
            sine_reg0   <= 36'sb100110111000010000010010110000001001;
        end
        14031: begin
            cosine_reg0 <= 36'sb10011110101010000101100100101111101;
            sine_reg0   <= 36'sb100110111000101111011100000001001100;
        end
        14032: begin
            cosine_reg0 <= 36'sb10011110101111000001000111000110001;
            sine_reg0   <= 36'sb100110111001001110100110010000001100;
        end
        14033: begin
            cosine_reg0 <= 36'sb10011110110011111100100011010100111;
            sine_reg0   <= 36'sb100110111001101101110001011101001000;
        end
        14034: begin
            cosine_reg0 <= 36'sb10011110111000110111111001011011110;
            sine_reg0   <= 36'sb100110111010001100111101101000000000;
        end
        14035: begin
            cosine_reg0 <= 36'sb10011110111101110011001001011010110;
            sine_reg0   <= 36'sb100110111010101100001010110000110010;
        end
        14036: begin
            cosine_reg0 <= 36'sb10011111000010101110010011010001011;
            sine_reg0   <= 36'sb100110111011001011011000110111011101;
        end
        14037: begin
            cosine_reg0 <= 36'sb10011111000111101001010110111111101;
            sine_reg0   <= 36'sb100110111011101010100111111100000000;
        end
        14038: begin
            cosine_reg0 <= 36'sb10011111001100100100010100100101010;
            sine_reg0   <= 36'sb100110111100001001110111111110011001;
        end
        14039: begin
            cosine_reg0 <= 36'sb10011111010001011111001100000010000;
            sine_reg0   <= 36'sb100110111100101001001000111110101000;
        end
        14040: begin
            cosine_reg0 <= 36'sb10011111010110011001111101010101111;
            sine_reg0   <= 36'sb100110111101001000011010111100101011;
        end
        14041: begin
            cosine_reg0 <= 36'sb10011111011011010100101000100000100;
            sine_reg0   <= 36'sb100110111101100111101101111000100001;
        end
        14042: begin
            cosine_reg0 <= 36'sb10011111100000001111001101100001110;
            sine_reg0   <= 36'sb100110111110000111000001110010001000;
        end
        14043: begin
            cosine_reg0 <= 36'sb10011111100101001001101100011001100;
            sine_reg0   <= 36'sb100110111110100110010110101001100000;
        end
        14044: begin
            cosine_reg0 <= 36'sb10011111101010000100000101000111100;
            sine_reg0   <= 36'sb100110111111000101101100011110100111;
        end
        14045: begin
            cosine_reg0 <= 36'sb10011111101110111110010111101011100;
            sine_reg0   <= 36'sb100110111111100101000011010001011101;
        end
        14046: begin
            cosine_reg0 <= 36'sb10011111110011111000100100000101011;
            sine_reg0   <= 36'sb100111000000000100011011000001111111;
        end
        14047: begin
            cosine_reg0 <= 36'sb10011111111000110010101010010101000;
            sine_reg0   <= 36'sb100111000000100011110011110000001101;
        end
        14048: begin
            cosine_reg0 <= 36'sb10011111111101101100101010011010001;
            sine_reg0   <= 36'sb100111000001000011001101011100000101;
        end
        14049: begin
            cosine_reg0 <= 36'sb10100000000010100110100100010100100;
            sine_reg0   <= 36'sb100111000001100010101000000101100110;
        end
        14050: begin
            cosine_reg0 <= 36'sb10100000000111100000011000000100000;
            sine_reg0   <= 36'sb100111000010000010000011101100110000;
        end
        14051: begin
            cosine_reg0 <= 36'sb10100000001100011010000101101000011;
            sine_reg0   <= 36'sb100111000010100001100000010001100001;
        end
        14052: begin
            cosine_reg0 <= 36'sb10100000010001010011101101000001101;
            sine_reg0   <= 36'sb100111000011000000111101110011110111;
        end
        14053: begin
            cosine_reg0 <= 36'sb10100000010110001101001110001111010;
            sine_reg0   <= 36'sb100111000011100000011100010011110001;
        end
        14054: begin
            cosine_reg0 <= 36'sb10100000011011000110101001010001011;
            sine_reg0   <= 36'sb100111000011111111111011110001001111;
        end
        14055: begin
            cosine_reg0 <= 36'sb10100000011111111111111110000111101;
            sine_reg0   <= 36'sb100111000100011111011100001100001110;
        end
        14056: begin
            cosine_reg0 <= 36'sb10100000100100111001001100110001111;
            sine_reg0   <= 36'sb100111000100111110111101100100101111;
        end
        14057: begin
            cosine_reg0 <= 36'sb10100000101001110010010101001111111;
            sine_reg0   <= 36'sb100111000101011110011111111010101111;
        end
        14058: begin
            cosine_reg0 <= 36'sb10100000101110101011010111100001100;
            sine_reg0   <= 36'sb100111000101111110000011001110001101;
        end
        14059: begin
            cosine_reg0 <= 36'sb10100000110011100100010011100110100;
            sine_reg0   <= 36'sb100111000110011101100111011111001000;
        end
        14060: begin
            cosine_reg0 <= 36'sb10100000111000011101001001011110110;
            sine_reg0   <= 36'sb100111000110111101001100101101011111;
        end
        14061: begin
            cosine_reg0 <= 36'sb10100000111101010101111001001010001;
            sine_reg0   <= 36'sb100111000111011100110010111001010001;
        end
        14062: begin
            cosine_reg0 <= 36'sb10100001000010001110100010101000010;
            sine_reg0   <= 36'sb100111000111111100011010000010011101;
        end
        14063: begin
            cosine_reg0 <= 36'sb10100001000111000111000101111001001;
            sine_reg0   <= 36'sb100111001000011100000010001001000000;
        end
        14064: begin
            cosine_reg0 <= 36'sb10100001001011111111100010111100011;
            sine_reg0   <= 36'sb100111001000111011101011001100111011;
        end
        14065: begin
            cosine_reg0 <= 36'sb10100001010000110111111001110010000;
            sine_reg0   <= 36'sb100111001001011011010101001110001100;
        end
        14066: begin
            cosine_reg0 <= 36'sb10100001010101110000001010011001101;
            sine_reg0   <= 36'sb100111001001111011000000001100110001;
        end
        14067: begin
            cosine_reg0 <= 36'sb10100001011010101000010100110011010;
            sine_reg0   <= 36'sb100111001010011010101100001000101001;
        end
        14068: begin
            cosine_reg0 <= 36'sb10100001011111100000011000111110100;
            sine_reg0   <= 36'sb100111001010111010011001000001110100;
        end
        14069: begin
            cosine_reg0 <= 36'sb10100001100100011000010110111011011;
            sine_reg0   <= 36'sb100111001011011010000110111000001111;
        end
        14070: begin
            cosine_reg0 <= 36'sb10100001101001010000001110101001101;
            sine_reg0   <= 36'sb100111001011111001110101101011111010;
        end
        14071: begin
            cosine_reg0 <= 36'sb10100001101110001000000000001000111;
            sine_reg0   <= 36'sb100111001100011001100101011100110100;
        end
        14072: begin
            cosine_reg0 <= 36'sb10100001110010111111101011011001010;
            sine_reg0   <= 36'sb100111001100111001010110001010111011;
        end
        14073: begin
            cosine_reg0 <= 36'sb10100001110111110111010000011010011;
            sine_reg0   <= 36'sb100111001101011001000111110110001110;
        end
        14074: begin
            cosine_reg0 <= 36'sb10100001111100101110101111001100000;
            sine_reg0   <= 36'sb100111001101111000111010011110101011;
        end
        14075: begin
            cosine_reg0 <= 36'sb10100010000001100110000111101110001;
            sine_reg0   <= 36'sb100111001110011000101110000100010011;
        end
        14076: begin
            cosine_reg0 <= 36'sb10100010000110011101011010000000100;
            sine_reg0   <= 36'sb100111001110111000100010100111000010;
        end
        14077: begin
            cosine_reg0 <= 36'sb10100010001011010100100110000010111;
            sine_reg0   <= 36'sb100111001111011000011000000110111001;
        end
        14078: begin
            cosine_reg0 <= 36'sb10100010010000001011101011110101000;
            sine_reg0   <= 36'sb100111001111111000001110100011110110;
        end
        14079: begin
            cosine_reg0 <= 36'sb10100010010101000010101011010110111;
            sine_reg0   <= 36'sb100111010000011000000101111101110111;
        end
        14080: begin
            cosine_reg0 <= 36'sb10100010011001111001100100101000010;
            sine_reg0   <= 36'sb100111010000110111111110010100111100;
        end
        14081: begin
            cosine_reg0 <= 36'sb10100010011110110000010111101000111;
            sine_reg0   <= 36'sb100111010001010111110111101001000010;
        end
        14082: begin
            cosine_reg0 <= 36'sb10100010100011100111000100011000100;
            sine_reg0   <= 36'sb100111010001110111110001111010001010;
        end
        14083: begin
            cosine_reg0 <= 36'sb10100010101000011101101010110111001;
            sine_reg0   <= 36'sb100111010010010111101101001000010010;
        end
        14084: begin
            cosine_reg0 <= 36'sb10100010101101010100001011000100100;
            sine_reg0   <= 36'sb100111010010110111101001010011011000;
        end
        14085: begin
            cosine_reg0 <= 36'sb10100010110010001010100101000000011;
            sine_reg0   <= 36'sb100111010011010111100110011011011100;
        end
        14086: begin
            cosine_reg0 <= 36'sb10100010110111000000111000101010100;
            sine_reg0   <= 36'sb100111010011110111100100100000011011;
        end
        14087: begin
            cosine_reg0 <= 36'sb10100010111011110111000110000010111;
            sine_reg0   <= 36'sb100111010100010111100011100010010101;
        end
        14088: begin
            cosine_reg0 <= 36'sb10100011000000101101001101001001010;
            sine_reg0   <= 36'sb100111010100110111100011100001001001;
        end
        14089: begin
            cosine_reg0 <= 36'sb10100011000101100011001101111101011;
            sine_reg0   <= 36'sb100111010101010111100100011100110101;
        end
        14090: begin
            cosine_reg0 <= 36'sb10100011001010011001001000011111001;
            sine_reg0   <= 36'sb100111010101110111100110010101011001;
        end
        14091: begin
            cosine_reg0 <= 36'sb10100011001111001110111100101110010;
            sine_reg0   <= 36'sb100111010110010111101001001010110010;
        end
        14092: begin
            cosine_reg0 <= 36'sb10100011010100000100101010101010101;
            sine_reg0   <= 36'sb100111010110110111101100111101000000;
        end
        14093: begin
            cosine_reg0 <= 36'sb10100011011000111010010010010100001;
            sine_reg0   <= 36'sb100111010111010111110001101100000001;
        end
        14094: begin
            cosine_reg0 <= 36'sb10100011011101101111110011101010011;
            sine_reg0   <= 36'sb100111010111110111110111010111110101;
        end
        14095: begin
            cosine_reg0 <= 36'sb10100011100010100101001110101101010;
            sine_reg0   <= 36'sb100111011000010111111110000000011001;
        end
        14096: begin
            cosine_reg0 <= 36'sb10100011100111011010100011011100101;
            sine_reg0   <= 36'sb100111011000111000000101100101101101;
        end
        14097: begin
            cosine_reg0 <= 36'sb10100011101100001111110001111000011;
            sine_reg0   <= 36'sb100111011001011000001110000111110000;
        end
        14098: begin
            cosine_reg0 <= 36'sb10100011110001000100111010000000010;
            sine_reg0   <= 36'sb100111011001111000010111100110100000;
        end
        14099: begin
            cosine_reg0 <= 36'sb10100011110101111001111011110100000;
            sine_reg0   <= 36'sb100111011010011000100010000001111011;
        end
        14100: begin
            cosine_reg0 <= 36'sb10100011111010101110110111010011011;
            sine_reg0   <= 36'sb100111011010111000101101011010000010;
        end
        14101: begin
            cosine_reg0 <= 36'sb10100011111111100011101100011110011;
            sine_reg0   <= 36'sb100111011011011000111001101110110010;
        end
        14102: begin
            cosine_reg0 <= 36'sb10100100000100011000011011010100111;
            sine_reg0   <= 36'sb100111011011111001000111000000001010;
        end
        14103: begin
            cosine_reg0 <= 36'sb10100100001001001101000011110110011;
            sine_reg0   <= 36'sb100111011100011001010101001110001010;
        end
        14104: begin
            cosine_reg0 <= 36'sb10100100001110000001100110000011000;
            sine_reg0   <= 36'sb100111011100111001100100011000101111;
        end
        14105: begin
            cosine_reg0 <= 36'sb10100100010010110110000001111010010;
            sine_reg0   <= 36'sb100111011101011001110100011111111000;
        end
        14106: begin
            cosine_reg0 <= 36'sb10100100010111101010010111011100010;
            sine_reg0   <= 36'sb100111011101111010000101100011100101;
        end
        14107: begin
            cosine_reg0 <= 36'sb10100100011100011110100110101000110;
            sine_reg0   <= 36'sb100111011110011010010111100011110100;
        end
        14108: begin
            cosine_reg0 <= 36'sb10100100100001010010101111011111011;
            sine_reg0   <= 36'sb100111011110111010101010100000100100;
        end
        14109: begin
            cosine_reg0 <= 36'sb10100100100110000110110010000000001;
            sine_reg0   <= 36'sb100111011111011010111110011001110011;
        end
        14110: begin
            cosine_reg0 <= 36'sb10100100101010111010101110001010101;
            sine_reg0   <= 36'sb100111011111111011010011001111100001;
        end
        14111: begin
            cosine_reg0 <= 36'sb10100100101111101110100011111111000;
            sine_reg0   <= 36'sb100111100000011011101001000001101100;
        end
        14112: begin
            cosine_reg0 <= 36'sb10100100110100100010010011011100110;
            sine_reg0   <= 36'sb100111100000111011111111110000010010;
        end
        14113: begin
            cosine_reg0 <= 36'sb10100100111001010101111100100011111;
            sine_reg0   <= 36'sb100111100001011100010111011011010011;
        end
        14114: begin
            cosine_reg0 <= 36'sb10100100111110001001011111010100001;
            sine_reg0   <= 36'sb100111100001111100110000000010101110;
        end
        14115: begin
            cosine_reg0 <= 36'sb10100101000010111100111011101101011;
            sine_reg0   <= 36'sb100111100010011101001001100110100000;
        end
        14116: begin
            cosine_reg0 <= 36'sb10100101000111110000010001101111011;
            sine_reg0   <= 36'sb100111100010111101100100000110101010;
        end
        14117: begin
            cosine_reg0 <= 36'sb10100101001100100011100001011001111;
            sine_reg0   <= 36'sb100111100011011101111111100011001000;
        end
        14118: begin
            cosine_reg0 <= 36'sb10100101010001010110101010101100110;
            sine_reg0   <= 36'sb100111100011111110011011111011111100;
        end
        14119: begin
            cosine_reg0 <= 36'sb10100101010110001001101101101000000;
            sine_reg0   <= 36'sb100111100100011110111001010001000010;
        end
        14120: begin
            cosine_reg0 <= 36'sb10100101011010111100101010001011001;
            sine_reg0   <= 36'sb100111100100111111010111100010011010;
        end
        14121: begin
            cosine_reg0 <= 36'sb10100101011111101111100000010110001;
            sine_reg0   <= 36'sb100111100101011111110110110000000011;
        end
        14122: begin
            cosine_reg0 <= 36'sb10100101100100100010010000001000111;
            sine_reg0   <= 36'sb100111100110000000010110111001111011;
        end
        14123: begin
            cosine_reg0 <= 36'sb10100101101001010100111001100011000;
            sine_reg0   <= 36'sb100111100110100000111000000000000001;
        end
        14124: begin
            cosine_reg0 <= 36'sb10100101101110000111011100100100011;
            sine_reg0   <= 36'sb100111100111000001011010000010010100;
        end
        14125: begin
            cosine_reg0 <= 36'sb10100101110010111001111001001101000;
            sine_reg0   <= 36'sb100111100111100001111101000000110010;
        end
        14126: begin
            cosine_reg0 <= 36'sb10100101110111101100001111011100011;
            sine_reg0   <= 36'sb100111101000000010100000111011011011;
        end
        14127: begin
            cosine_reg0 <= 36'sb10100101111100011110011111010010101;
            sine_reg0   <= 36'sb100111101000100011000101110010001101;
        end
        14128: begin
            cosine_reg0 <= 36'sb10100110000001010000101000101111010;
            sine_reg0   <= 36'sb100111101001000011101011100101000110;
        end
        14129: begin
            cosine_reg0 <= 36'sb10100110000110000010101011110010011;
            sine_reg0   <= 36'sb100111101001100100010010010100000111;
        end
        14130: begin
            cosine_reg0 <= 36'sb10100110001010110100101000011011101;
            sine_reg0   <= 36'sb100111101010000100111001111111001100;
        end
        14131: begin
            cosine_reg0 <= 36'sb10100110001111100110011110101010111;
            sine_reg0   <= 36'sb100111101010100101100010100110010101;
        end
        14132: begin
            cosine_reg0 <= 36'sb10100110010100011000001110100000000;
            sine_reg0   <= 36'sb100111101011000110001100001001100010;
        end
        14133: begin
            cosine_reg0 <= 36'sb10100110011001001001110111111010101;
            sine_reg0   <= 36'sb100111101011100110110110101000101111;
        end
        14134: begin
            cosine_reg0 <= 36'sb10100110011101111011011010111010111;
            sine_reg0   <= 36'sb100111101100000111100010000011111101;
        end
        14135: begin
            cosine_reg0 <= 36'sb10100110100010101100110111100000010;
            sine_reg0   <= 36'sb100111101100101000001110011011001010;
        end
        14136: begin
            cosine_reg0 <= 36'sb10100110100111011110001101101010110;
            sine_reg0   <= 36'sb100111101101001000111011101110010101;
        end
        14137: begin
            cosine_reg0 <= 36'sb10100110101100001111011101011010000;
            sine_reg0   <= 36'sb100111101101101001101001111101011100;
        end
        14138: begin
            cosine_reg0 <= 36'sb10100110110001000000100110101110001;
            sine_reg0   <= 36'sb100111101110001010011001001000011110;
        end
        14139: begin
            cosine_reg0 <= 36'sb10100110110101110001101001100110110;
            sine_reg0   <= 36'sb100111101110101011001001001111011011;
        end
        14140: begin
            cosine_reg0 <= 36'sb10100110111010100010100110000011101;
            sine_reg0   <= 36'sb100111101111001011111010010010010000;
        end
        14141: begin
            cosine_reg0 <= 36'sb10100110111111010011011100000100110;
            sine_reg0   <= 36'sb100111101111101100101100010000111100;
        end
        14142: begin
            cosine_reg0 <= 36'sb10100111000100000100001011101001110;
            sine_reg0   <= 36'sb100111110000001101011111001011011110;
        end
        14143: begin
            cosine_reg0 <= 36'sb10100111001000110100110100110010101;
            sine_reg0   <= 36'sb100111110000101110010011000001110110;
        end
        14144: begin
            cosine_reg0 <= 36'sb10100111001101100101010111011111000;
            sine_reg0   <= 36'sb100111110001001111000111110100000001;
        end
        14145: begin
            cosine_reg0 <= 36'sb10100111010010010101110011101110111;
            sine_reg0   <= 36'sb100111110001101111111101100001111110;
        end
        14146: begin
            cosine_reg0 <= 36'sb10100111010111000110001001100010000;
            sine_reg0   <= 36'sb100111110010010000110100001011101101;
        end
        14147: begin
            cosine_reg0 <= 36'sb10100111011011110110011000111000001;
            sine_reg0   <= 36'sb100111110010110001101011110001001011;
        end
        14148: begin
            cosine_reg0 <= 36'sb10100111100000100110100001110001001;
            sine_reg0   <= 36'sb100111110011010010100100010010011000;
        end
        14149: begin
            cosine_reg0 <= 36'sb10100111100101010110100100001100111;
            sine_reg0   <= 36'sb100111110011110011011101101111010010;
        end
        14150: begin
            cosine_reg0 <= 36'sb10100111101010000110100000001011001;
            sine_reg0   <= 36'sb100111110100010100011000000111111000;
        end
        14151: begin
            cosine_reg0 <= 36'sb10100111101110110110010101101011101;
            sine_reg0   <= 36'sb100111110100110101010011011100001001;
        end
        14152: begin
            cosine_reg0 <= 36'sb10100111110011100110000100101110011;
            sine_reg0   <= 36'sb100111110101010110001111101100000011;
        end
        14153: begin
            cosine_reg0 <= 36'sb10100111111000010101101101010011000;
            sine_reg0   <= 36'sb100111110101110111001100110111100110;
        end
        14154: begin
            cosine_reg0 <= 36'sb10100111111101000101001111011001011;
            sine_reg0   <= 36'sb100111110110011000001010111110110000;
        end
        14155: begin
            cosine_reg0 <= 36'sb10101000000001110100101011000001011;
            sine_reg0   <= 36'sb100111110110111001001010000001011111;
        end
        14156: begin
            cosine_reg0 <= 36'sb10101000000110100100000000001010110;
            sine_reg0   <= 36'sb100111110111011010001001111111110010;
        end
        14157: begin
            cosine_reg0 <= 36'sb10101000001011010011001110110101011;
            sine_reg0   <= 36'sb100111110111111011001010111001101001;
        end
        14158: begin
            cosine_reg0 <= 36'sb10101000010000000010010111000001000;
            sine_reg0   <= 36'sb100111111000011100001100101111000010;
        end
        14159: begin
            cosine_reg0 <= 36'sb10101000010100110001011000101101100;
            sine_reg0   <= 36'sb100111111000111101001111011111111011;
        end
        14160: begin
            cosine_reg0 <= 36'sb10101000011001100000010011111010110;
            sine_reg0   <= 36'sb100111111001011110010011001100010011;
        end
        14161: begin
            cosine_reg0 <= 36'sb10101000011110001111001000101000011;
            sine_reg0   <= 36'sb100111111001111111010111110100001010;
        end
        14162: begin
            cosine_reg0 <= 36'sb10101000100010111101110110110110011;
            sine_reg0   <= 36'sb100111111010100000011101010111011101;
        end
        14163: begin
            cosine_reg0 <= 36'sb10101000100111101100011110100100100;
            sine_reg0   <= 36'sb100111111011000001100011110110001100;
        end
        14164: begin
            cosine_reg0 <= 36'sb10101000101100011010111111110010101;
            sine_reg0   <= 36'sb100111111011100010101011010000010101;
        end
        14165: begin
            cosine_reg0 <= 36'sb10101000110001001001011010100000100;
            sine_reg0   <= 36'sb100111111100000011110011100101110111;
        end
        14166: begin
            cosine_reg0 <= 36'sb10101000110101110111101110101101111;
            sine_reg0   <= 36'sb100111111100100100111100110110110000;
        end
        14167: begin
            cosine_reg0 <= 36'sb10101000111010100101111100011010101;
            sine_reg0   <= 36'sb100111111101000110000111000011000000;
        end
        14168: begin
            cosine_reg0 <= 36'sb10101000111111010100000011100110110;
            sine_reg0   <= 36'sb100111111101100111010010001010100101;
        end
        14169: begin
            cosine_reg0 <= 36'sb10101001000100000010000100010001110;
            sine_reg0   <= 36'sb100111111110001000011110001101011110;
        end
        14170: begin
            cosine_reg0 <= 36'sb10101001001000101111111110011011110;
            sine_reg0   <= 36'sb100111111110101001101011001011101001;
        end
        14171: begin
            cosine_reg0 <= 36'sb10101001001101011101110010000100011;
            sine_reg0   <= 36'sb100111111111001010111001000101000110;
        end
        14172: begin
            cosine_reg0 <= 36'sb10101001010010001011011111001011011;
            sine_reg0   <= 36'sb100111111111101100000111111001110011;
        end
        14173: begin
            cosine_reg0 <= 36'sb10101001010110111001000101110000110;
            sine_reg0   <= 36'sb101000000000001101010111101001101110;
        end
        14174: begin
            cosine_reg0 <= 36'sb10101001011011100110100101110100011;
            sine_reg0   <= 36'sb101000000000101110101000010100110110;
        end
        14175: begin
            cosine_reg0 <= 36'sb10101001100000010011111111010101110;
            sine_reg0   <= 36'sb101000000001001111111001111011001011;
        end
        14176: begin
            cosine_reg0 <= 36'sb10101001100101000001010010010101000;
            sine_reg0   <= 36'sb101000000001110001001100011100101011;
        end
        14177: begin
            cosine_reg0 <= 36'sb10101001101001101110011110110001111;
            sine_reg0   <= 36'sb101000000010010010011111111001010100;
        end
        14178: begin
            cosine_reg0 <= 36'sb10101001101110011011100100101100000;
            sine_reg0   <= 36'sb101000000010110011110100010001000110;
        end
        14179: begin
            cosine_reg0 <= 36'sb10101001110011001000100100000011100;
            sine_reg0   <= 36'sb101000000011010101001001100011111110;
        end
        14180: begin
            cosine_reg0 <= 36'sb10101001110111110101011100111000000;
            sine_reg0   <= 36'sb101000000011110110011111110001111100;
        end
        14181: begin
            cosine_reg0 <= 36'sb10101001111100100010001111001001010;
            sine_reg0   <= 36'sb101000000100010111110110111010111111;
        end
        14182: begin
            cosine_reg0 <= 36'sb10101010000001001110111010110111010;
            sine_reg0   <= 36'sb101000000100111001001110111111000101;
        end
        14183: begin
            cosine_reg0 <= 36'sb10101010000101111011100000000001110;
            sine_reg0   <= 36'sb101000000101011010100111111110001100;
        end
        14184: begin
            cosine_reg0 <= 36'sb10101010001010100111111110101000101;
            sine_reg0   <= 36'sb101000000101111100000001111000010101;
        end
        14185: begin
            cosine_reg0 <= 36'sb10101010001111010100010110101011100;
            sine_reg0   <= 36'sb101000000110011101011100101101011100;
        end
        14186: begin
            cosine_reg0 <= 36'sb10101010010100000000101000001010011;
            sine_reg0   <= 36'sb101000000110111110111000011101100010;
        end
        14187: begin
            cosine_reg0 <= 36'sb10101010011000101100110011000101001;
            sine_reg0   <= 36'sb101000000111100000010101001000100100;
        end
        14188: begin
            cosine_reg0 <= 36'sb10101010011101011000110111011011011;
            sine_reg0   <= 36'sb101000001000000001110010101110100001;
        end
        14189: begin
            cosine_reg0 <= 36'sb10101010100010000100110101001101000;
            sine_reg0   <= 36'sb101000001000100011010001001111011001;
        end
        14190: begin
            cosine_reg0 <= 36'sb10101010100110110000101100011001111;
            sine_reg0   <= 36'sb101000001001000100110000101011001010;
        end
        14191: begin
            cosine_reg0 <= 36'sb10101010101011011100011101000001111;
            sine_reg0   <= 36'sb101000001001100110010001000001110010;
        end
        14192: begin
            cosine_reg0 <= 36'sb10101010110000001000000111000100101;
            sine_reg0   <= 36'sb101000001010000111110010010011010000;
        end
        14193: begin
            cosine_reg0 <= 36'sb10101010110100110011101010100010001;
            sine_reg0   <= 36'sb101000001010101001010100011111100011;
        end
        14194: begin
            cosine_reg0 <= 36'sb10101010111001011111000111011010001;
            sine_reg0   <= 36'sb101000001011001010110111100110101010;
        end
        14195: begin
            cosine_reg0 <= 36'sb10101010111110001010011101101100100;
            sine_reg0   <= 36'sb101000001011101100011011101000100011;
        end
        14196: begin
            cosine_reg0 <= 36'sb10101011000010110101101101011000111;
            sine_reg0   <= 36'sb101000001100001110000000100101001110;
        end
        14197: begin
            cosine_reg0 <= 36'sb10101011000111100000110110011111011;
            sine_reg0   <= 36'sb101000001100101111100110011100101000;
        end
        14198: begin
            cosine_reg0 <= 36'sb10101011001100001011111000111111101;
            sine_reg0   <= 36'sb101000001101010001001101001110110001;
        end
        14199: begin
            cosine_reg0 <= 36'sb10101011010000110110110100111001011;
            sine_reg0   <= 36'sb101000001101110010110100111011100110;
        end
        14200: begin
            cosine_reg0 <= 36'sb10101011010101100001101010001100101;
            sine_reg0   <= 36'sb101000001110010100011101100011001000;
        end
        14201: begin
            cosine_reg0 <= 36'sb10101011011010001100011000111001001;
            sine_reg0   <= 36'sb101000001110110110000111000101010100;
        end
        14202: begin
            cosine_reg0 <= 36'sb10101011011110110111000000111110110;
            sine_reg0   <= 36'sb101000001111010111110001100010001010;
        end
        14203: begin
            cosine_reg0 <= 36'sb10101011100011100001100010011101001;
            sine_reg0   <= 36'sb101000001111111001011100111001101000;
        end
        14204: begin
            cosine_reg0 <= 36'sb10101011101000001011111101010100010;
            sine_reg0   <= 36'sb101000010000011011001001001011101100;
        end
        14205: begin
            cosine_reg0 <= 36'sb10101011101100110110010001100100000;
            sine_reg0   <= 36'sb101000010000111100110110011000010110;
        end
        14206: begin
            cosine_reg0 <= 36'sb10101011110001100000011111001100000;
            sine_reg0   <= 36'sb101000010001011110100100011111100011;
        end
        14207: begin
            cosine_reg0 <= 36'sb10101011110110001010100110001100001;
            sine_reg0   <= 36'sb101000010010000000010011100001010100;
        end
        14208: begin
            cosine_reg0 <= 36'sb10101011111010110100100110100100011;
            sine_reg0   <= 36'sb101000010010100010000011011101100110;
        end
        14209: begin
            cosine_reg0 <= 36'sb10101011111111011110100000010100010;
            sine_reg0   <= 36'sb101000010011000011110100010100011000;
        end
        14210: begin
            cosine_reg0 <= 36'sb10101100000100001000010011011011111;
            sine_reg0   <= 36'sb101000010011100101100110000101101010;
        end
        14211: begin
            cosine_reg0 <= 36'sb10101100001000110001111111111011000;
            sine_reg0   <= 36'sb101000010100000111011000110001011000;
        end
        14212: begin
            cosine_reg0 <= 36'sb10101100001101011011100101110001010;
            sine_reg0   <= 36'sb101000010100101001001100010111100100;
        end
        14213: begin
            cosine_reg0 <= 36'sb10101100010010000101000100111110101;
            sine_reg0   <= 36'sb101000010101001011000000111000001010;
        end
        14214: begin
            cosine_reg0 <= 36'sb10101100010110101110011101100011000;
            sine_reg0   <= 36'sb101000010101101100110110010011001001;
        end
        14215: begin
            cosine_reg0 <= 36'sb10101100011011010111101111011110000;
            sine_reg0   <= 36'sb101000010110001110101100101000100010;
        end
        14216: begin
            cosine_reg0 <= 36'sb10101100100000000000111010101111101;
            sine_reg0   <= 36'sb101000010110110000100011111000010001;
        end
        14217: begin
            cosine_reg0 <= 36'sb10101100100100101001111111010111101;
            sine_reg0   <= 36'sb101000010111010010011100000010010110;
        end
        14218: begin
            cosine_reg0 <= 36'sb10101100101001010010111101010101110;
            sine_reg0   <= 36'sb101000010111110100010101000110101111;
        end
        14219: begin
            cosine_reg0 <= 36'sb10101100101101111011110100101010000;
            sine_reg0   <= 36'sb101000011000010110001111000101011100;
        end
        14220: begin
            cosine_reg0 <= 36'sb10101100110010100100100101010100000;
            sine_reg0   <= 36'sb101000011000111000001001111110011011;
        end
        14221: begin
            cosine_reg0 <= 36'sb10101100110111001101001111010011101;
            sine_reg0   <= 36'sb101000011001011010000101110001101010;
        end
        14222: begin
            cosine_reg0 <= 36'sb10101100111011110101110010101000110;
            sine_reg0   <= 36'sb101000011001111100000010011111001000;
        end
        14223: begin
            cosine_reg0 <= 36'sb10101101000000011110001111010011010;
            sine_reg0   <= 36'sb101000011010011110000000000110110100;
        end
        14224: begin
            cosine_reg0 <= 36'sb10101101000101000110100101010010111;
            sine_reg0   <= 36'sb101000011010111111111110101000101101;
        end
        14225: begin
            cosine_reg0 <= 36'sb10101101001001101110110100100111011;
            sine_reg0   <= 36'sb101000011011100001111110000100110001;
        end
        14226: begin
            cosine_reg0 <= 36'sb10101101001110010110111101010000101;
            sine_reg0   <= 36'sb101000011100000011111110011010111111;
        end
        14227: begin
            cosine_reg0 <= 36'sb10101101010010111110111111001110100;
            sine_reg0   <= 36'sb101000011100100101111111101011010110;
        end
        14228: begin
            cosine_reg0 <= 36'sb10101101010111100110111010100000110;
            sine_reg0   <= 36'sb101000011101001000000001110101110100;
        end
        14229: begin
            cosine_reg0 <= 36'sb10101101011100001110101111000111010;
            sine_reg0   <= 36'sb101000011101101010000100111010011000;
        end
        14230: begin
            cosine_reg0 <= 36'sb10101101100000110110011101000001111;
            sine_reg0   <= 36'sb101000011110001100001000111001000010;
        end
        14231: begin
            cosine_reg0 <= 36'sb10101101100101011110000100010000010;
            sine_reg0   <= 36'sb101000011110101110001101110001101110;
        end
        14232: begin
            cosine_reg0 <= 36'sb10101101101010000101100100110010011;
            sine_reg0   <= 36'sb101000011111010000010011100100011101;
        end
        14233: begin
            cosine_reg0 <= 36'sb10101101101110101100111110101000000;
            sine_reg0   <= 36'sb101000011111110010011010010001001100;
        end
        14234: begin
            cosine_reg0 <= 36'sb10101101110011010100010001110001000;
            sine_reg0   <= 36'sb101000100000010100100001110111111011;
        end
        14235: begin
            cosine_reg0 <= 36'sb10101101110111111011011110001101001;
            sine_reg0   <= 36'sb101000100000110110101010011000101000;
        end
        14236: begin
            cosine_reg0 <= 36'sb10101101111100100010100011111100010;
            sine_reg0   <= 36'sb101000100001011000110011110011010010;
        end
        14237: begin
            cosine_reg0 <= 36'sb10101110000001001001100010111110010;
            sine_reg0   <= 36'sb101000100001111010111110000111110111;
        end
        14238: begin
            cosine_reg0 <= 36'sb10101110000101110000011011010010110;
            sine_reg0   <= 36'sb101000100010011101001001010110010111;
        end
        14239: begin
            cosine_reg0 <= 36'sb10101110001010010111001100111001110;
            sine_reg0   <= 36'sb101000100010111111010101011110110000;
        end
        14240: begin
            cosine_reg0 <= 36'sb10101110001110111101110111110011001;
            sine_reg0   <= 36'sb101000100011100001100010100001000000;
        end
        14241: begin
            cosine_reg0 <= 36'sb10101110010011100100011011111110100;
            sine_reg0   <= 36'sb101000100100000011110000011101000110;
        end
        14242: begin
            cosine_reg0 <= 36'sb10101110011000001010111001011011110;
            sine_reg0   <= 36'sb101000100100100101111111010011000010;
        end
        14243: begin
            cosine_reg0 <= 36'sb10101110011100110001010000001010110;
            sine_reg0   <= 36'sb101000100101001000001111000010110001;
        end
        14244: begin
            cosine_reg0 <= 36'sb10101110100001010111100000001011011;
            sine_reg0   <= 36'sb101000100101101010011111101100010010;
        end
        14245: begin
            cosine_reg0 <= 36'sb10101110100101111101101001011101011;
            sine_reg0   <= 36'sb101000100110001100110001001111100101;
        end
        14246: begin
            cosine_reg0 <= 36'sb10101110101010100011101100000000100;
            sine_reg0   <= 36'sb101000100110101111000011101100100111;
        end
        14247: begin
            cosine_reg0 <= 36'sb10101110101111001001100111110100110;
            sine_reg0   <= 36'sb101000100111010001010111000011010111;
        end
        14248: begin
            cosine_reg0 <= 36'sb10101110110011101111011100111001111;
            sine_reg0   <= 36'sb101000100111110011101011010011110101;
        end
        14249: begin
            cosine_reg0 <= 36'sb10101110111000010101001011001111101;
            sine_reg0   <= 36'sb101000101000010110000000011101111110;
        end
        14250: begin
            cosine_reg0 <= 36'sb10101110111100111010110010110101111;
            sine_reg0   <= 36'sb101000101000111000010110100001110001;
        end
        14251: begin
            cosine_reg0 <= 36'sb10101111000001100000010011101100100;
            sine_reg0   <= 36'sb101000101001011010101101011111001110;
        end
        14252: begin
            cosine_reg0 <= 36'sb10101111000110000101101101110011001;
            sine_reg0   <= 36'sb101000101001111101000101010110010010;
        end
        14253: begin
            cosine_reg0 <= 36'sb10101111001010101011000001001001111;
            sine_reg0   <= 36'sb101000101010011111011110000110111101;
        end
        14254: begin
            cosine_reg0 <= 36'sb10101111001111010000001101110000011;
            sine_reg0   <= 36'sb101000101011000001110111110001001101;
        end
        14255: begin
            cosine_reg0 <= 36'sb10101111010011110101010011100110100;
            sine_reg0   <= 36'sb101000101011100100010010010101000000;
        end
        14256: begin
            cosine_reg0 <= 36'sb10101111011000011010010010101100000;
            sine_reg0   <= 36'sb101000101100000110101101110010010111;
        end
        14257: begin
            cosine_reg0 <= 36'sb10101111011100111111001011000000111;
            sine_reg0   <= 36'sb101000101100101001001010001001001110;
        end
        14258: begin
            cosine_reg0 <= 36'sb10101111100001100011111100100100110;
            sine_reg0   <= 36'sb101000101101001011100111011001100101;
        end
        14259: begin
            cosine_reg0 <= 36'sb10101111100110001000100111010111100;
            sine_reg0   <= 36'sb101000101101101110000101100011011010;
        end
        14260: begin
            cosine_reg0 <= 36'sb10101111101010101101001011011001001;
            sine_reg0   <= 36'sb101000101110010000100100100110101100;
        end
        14261: begin
            cosine_reg0 <= 36'sb10101111101111010001101000101001001;
            sine_reg0   <= 36'sb101000101110110011000100100011011011;
        end
        14262: begin
            cosine_reg0 <= 36'sb10101111110011110101111111000111101;
            sine_reg0   <= 36'sb101000101111010101100101011001100011;
        end
        14263: begin
            cosine_reg0 <= 36'sb10101111111000011010001110110100011;
            sine_reg0   <= 36'sb101000101111111000000111001001000101;
        end
        14264: begin
            cosine_reg0 <= 36'sb10101111111100111110010111101111001;
            sine_reg0   <= 36'sb101000110000011010101001110001111111;
        end
        14265: begin
            cosine_reg0 <= 36'sb10110000000001100010011001110111101;
            sine_reg0   <= 36'sb101000110000111101001101010100001111;
        end
        14266: begin
            cosine_reg0 <= 36'sb10110000000110000110010101001101111;
            sine_reg0   <= 36'sb101000110001011111110001101111110100;
        end
        14267: begin
            cosine_reg0 <= 36'sb10110000001010101010001001110001101;
            sine_reg0   <= 36'sb101000110010000010010111000100101101;
        end
        14268: begin
            cosine_reg0 <= 36'sb10110000001111001101110111100010110;
            sine_reg0   <= 36'sb101000110010100100111101010010111001;
        end
        14269: begin
            cosine_reg0 <= 36'sb10110000010011110001011110100001000;
            sine_reg0   <= 36'sb101000110011000111100100011010010101;
        end
        14270: begin
            cosine_reg0 <= 36'sb10110000011000010100111110101100010;
            sine_reg0   <= 36'sb101000110011101010001100011011000010;
        end
        14271: begin
            cosine_reg0 <= 36'sb10110000011100111000011000000100010;
            sine_reg0   <= 36'sb101000110100001100110101010100111101;
        end
        14272: begin
            cosine_reg0 <= 36'sb10110000100001011011101010101000111;
            sine_reg0   <= 36'sb101000110100101111011111001000000101;
        end
        14273: begin
            cosine_reg0 <= 36'sb10110000100101111110110110011001111;
            sine_reg0   <= 36'sb101000110101010010001001110100011001;
        end
        14274: begin
            cosine_reg0 <= 36'sb10110000101010100001111011010111010;
            sine_reg0   <= 36'sb101000110101110100110101011001110111;
        end
        14275: begin
            cosine_reg0 <= 36'sb10110000101111000100111001100000110;
            sine_reg0   <= 36'sb101000110110010111100001111000011110;
        end
        14276: begin
            cosine_reg0 <= 36'sb10110000110011100111110000110110001;
            sine_reg0   <= 36'sb101000110110111010001111010000001101;
        end
        14277: begin
            cosine_reg0 <= 36'sb10110000111000001010100001010111010;
            sine_reg0   <= 36'sb101000110111011100111101100001000011;
        end
        14278: begin
            cosine_reg0 <= 36'sb10110000111100101101001011000011111;
            sine_reg0   <= 36'sb101000110111111111101100101010111110;
        end
        14279: begin
            cosine_reg0 <= 36'sb10110001000001001111101101111100000;
            sine_reg0   <= 36'sb101000111000100010011100101101111100;
        end
        14280: begin
            cosine_reg0 <= 36'sb10110001000101110010001001111111010;
            sine_reg0   <= 36'sb101000111001000101001101101001111101;
        end
        14281: begin
            cosine_reg0 <= 36'sb10110001001010010100011111001101101;
            sine_reg0   <= 36'sb101000111001100111111111011110111111;
        end
        14282: begin
            cosine_reg0 <= 36'sb10110001001110110110101101100110111;
            sine_reg0   <= 36'sb101000111010001010110010001101000001;
        end
        14283: begin
            cosine_reg0 <= 36'sb10110001010011011000110101001010110;
            sine_reg0   <= 36'sb101000111010101101100101110100000001;
        end
        14284: begin
            cosine_reg0 <= 36'sb10110001010111111010110101111001010;
            sine_reg0   <= 36'sb101000111011010000011010010011111110;
        end
        14285: begin
            cosine_reg0 <= 36'sb10110001011100011100101111110010000;
            sine_reg0   <= 36'sb101000111011110011001111101100110111;
        end
        14286: begin
            cosine_reg0 <= 36'sb10110001100000111110100010110101000;
            sine_reg0   <= 36'sb101000111100010110000101111110101011;
        end
        14287: begin
            cosine_reg0 <= 36'sb10110001100101100000001111000010000;
            sine_reg0   <= 36'sb101000111100111000111101001001010111;
        end
        14288: begin
            cosine_reg0 <= 36'sb10110001101010000001110100011000110;
            sine_reg0   <= 36'sb101000111101011011110101001100111011;
        end
        14289: begin
            cosine_reg0 <= 36'sb10110001101110100011010010111001010;
            sine_reg0   <= 36'sb101000111101111110101110001001010101;
        end
        14290: begin
            cosine_reg0 <= 36'sb10110001110011000100101010100011001;
            sine_reg0   <= 36'sb101000111110100001100111111110100101;
        end
        14291: begin
            cosine_reg0 <= 36'sb10110001110111100101111011010110011;
            sine_reg0   <= 36'sb101000111111000100100010101100101000;
        end
        14292: begin
            cosine_reg0 <= 36'sb10110001111100000111000101010010110;
            sine_reg0   <= 36'sb101000111111100111011110010011011101;
        end
        14293: begin
            cosine_reg0 <= 36'sb10110010000000101000001000011000000;
            sine_reg0   <= 36'sb101001000000001010011010110011000011;
        end
        14294: begin
            cosine_reg0 <= 36'sb10110010000101001001000100100110001;
            sine_reg0   <= 36'sb101001000000101101011000001011011001;
        end
        14295: begin
            cosine_reg0 <= 36'sb10110010001001101001111001111100110;
            sine_reg0   <= 36'sb101001000001010000010110011100011101;
        end
        14296: begin
            cosine_reg0 <= 36'sb10110010001110001010101000011011111;
            sine_reg0   <= 36'sb101001000001110011010101100110001110;
        end
        14297: begin
            cosine_reg0 <= 36'sb10110010010010101011010000000011010;
            sine_reg0   <= 36'sb101001000010010110010101101000101011;
        end
        14298: begin
            cosine_reg0 <= 36'sb10110010010111001011110000110010110;
            sine_reg0   <= 36'sb101001000010111001010110100011110010;
        end
        14299: begin
            cosine_reg0 <= 36'sb10110010011011101100001010101010001;
            sine_reg0   <= 36'sb101001000011011100011000010111100010;
        end
        14300: begin
            cosine_reg0 <= 36'sb10110010100000001100011101101001001;
            sine_reg0   <= 36'sb101001000011111111011011000011111001;
        end
        14301: begin
            cosine_reg0 <= 36'sb10110010100100101100101001101111111;
            sine_reg0   <= 36'sb101001000100100010011110101000110110;
        end
        14302: begin
            cosine_reg0 <= 36'sb10110010101001001100101110111101111;
            sine_reg0   <= 36'sb101001000101000101100011000110011001;
        end
        14303: begin
            cosine_reg0 <= 36'sb10110010101101101100101101010011001;
            sine_reg0   <= 36'sb101001000101101000101000011100011110;
        end
        14304: begin
            cosine_reg0 <= 36'sb10110010110010001100100100101111011;
            sine_reg0   <= 36'sb101001000110001011101110101011000110;
        end
        14305: begin
            cosine_reg0 <= 36'sb10110010110110101100010101010010101;
            sine_reg0   <= 36'sb101001000110101110110101110010001111;
        end
        14306: begin
            cosine_reg0 <= 36'sb10110010111011001011111110111100100;
            sine_reg0   <= 36'sb101001000111010001111101110001110111;
        end
        14307: begin
            cosine_reg0 <= 36'sb10110010111111101011100001101100111;
            sine_reg0   <= 36'sb101001000111110101000110101001111101;
        end
        14308: begin
            cosine_reg0 <= 36'sb10110011000100001010111101100011101;
            sine_reg0   <= 36'sb101001001000011000010000011010011111;
        end
        14309: begin
            cosine_reg0 <= 36'sb10110011001000101010010010100000100;
            sine_reg0   <= 36'sb101001001000111011011011000011011101;
        end
        14310: begin
            cosine_reg0 <= 36'sb10110011001101001001100000100011011;
            sine_reg0   <= 36'sb101001001001011110100110100100110101;
        end
        14311: begin
            cosine_reg0 <= 36'sb10110011010001101000100111101100001;
            sine_reg0   <= 36'sb101001001010000001110010111110100110;
        end
        14312: begin
            cosine_reg0 <= 36'sb10110011010110000111100111111010100;
            sine_reg0   <= 36'sb101001001010100101000000010000101110;
        end
        14313: begin
            cosine_reg0 <= 36'sb10110011011010100110100001001110011;
            sine_reg0   <= 36'sb101001001011001000001110011011001100;
        end
        14314: begin
            cosine_reg0 <= 36'sb10110011011111000101010011100111100;
            sine_reg0   <= 36'sb101001001011101011011101011101111110;
        end
        14315: begin
            cosine_reg0 <= 36'sb10110011100011100011111111000101111;
            sine_reg0   <= 36'sb101001001100001110101101011001000100;
        end
        14316: begin
            cosine_reg0 <= 36'sb10110011101000000010100011101001001;
            sine_reg0   <= 36'sb101001001100110001111110001100011011;
        end
        14317: begin
            cosine_reg0 <= 36'sb10110011101100100001000001010001010;
            sine_reg0   <= 36'sb101001001101010101001111111000000011;
        end
        14318: begin
            cosine_reg0 <= 36'sb10110011110000111111010111111101111;
            sine_reg0   <= 36'sb101001001101111000100010011011111010;
        end
        14319: begin
            cosine_reg0 <= 36'sb10110011110101011101100111101111000;
            sine_reg0   <= 36'sb101001001110011011110101110111111111;
        end
        14320: begin
            cosine_reg0 <= 36'sb10110011111001111011110000100100100;
            sine_reg0   <= 36'sb101001001110111111001010001100010000;
        end
        14321: begin
            cosine_reg0 <= 36'sb10110011111110011001110010011110000;
            sine_reg0   <= 36'sb101001001111100010011111011000101101;
        end
        14322: begin
            cosine_reg0 <= 36'sb10110100000010110111101101011011011;
            sine_reg0   <= 36'sb101001010000000101110101011101010010;
        end
        14323: begin
            cosine_reg0 <= 36'sb10110100000111010101100001011100101;
            sine_reg0   <= 36'sb101001010000101001001100011010000001;
        end
        14324: begin
            cosine_reg0 <= 36'sb10110100001011110011001110100001011;
            sine_reg0   <= 36'sb101001010001001100100100001110110110;
        end
        14325: begin
            cosine_reg0 <= 36'sb10110100010000010000110100101001101;
            sine_reg0   <= 36'sb101001010001101111111100111011110001;
        end
        14326: begin
            cosine_reg0 <= 36'sb10110100010100101110010011110101000;
            sine_reg0   <= 36'sb101001010010010011010110100000110000;
        end
        14327: begin
            cosine_reg0 <= 36'sb10110100011001001011101100000011100;
            sine_reg0   <= 36'sb101001010010110110110000111101110001;
        end
        14328: begin
            cosine_reg0 <= 36'sb10110100011101101000111101010101000;
            sine_reg0   <= 36'sb101001010011011010001100010010110101;
        end
        14329: begin
            cosine_reg0 <= 36'sb10110100100010000110000111101001001;
            sine_reg0   <= 36'sb101001010011111101101000011111111000;
        end
        14330: begin
            cosine_reg0 <= 36'sb10110100100110100011001010111111110;
            sine_reg0   <= 36'sb101001010100100001000101100100111010;
        end
        14331: begin
            cosine_reg0 <= 36'sb10110100101011000000000111011000111;
            sine_reg0   <= 36'sb101001010101000100100011100001111010;
        end
        14332: begin
            cosine_reg0 <= 36'sb10110100101111011100111100110100001;
            sine_reg0   <= 36'sb101001010101101000000010010110110110;
        end
        14333: begin
            cosine_reg0 <= 36'sb10110100110011111001101011010001011;
            sine_reg0   <= 36'sb101001010110001011100010000011101100;
        end
        14334: begin
            cosine_reg0 <= 36'sb10110100111000010110010010110000101;
            sine_reg0   <= 36'sb101001010110101111000010101000011011;
        end
        14335: begin
            cosine_reg0 <= 36'sb10110100111100110010110011010001100;
            sine_reg0   <= 36'sb101001010111010010100100000101000011;
        end
        14336: begin
            cosine_reg0 <= 36'sb10110101000001001111001100110011111;
            sine_reg0   <= 36'sb101001010111110110000110011001100001;
        end
        14337: begin
            cosine_reg0 <= 36'sb10110101000101101011011111010111101;
            sine_reg0   <= 36'sb101001011000011001101001100101110100;
        end
        14338: begin
            cosine_reg0 <= 36'sb10110101001010000111101010111100101;
            sine_reg0   <= 36'sb101001011000111101001101101001111011;
        end
        14339: begin
            cosine_reg0 <= 36'sb10110101001110100011101111100010100;
            sine_reg0   <= 36'sb101001011001100000110010100101110101;
        end
        14340: begin
            cosine_reg0 <= 36'sb10110101010010111111101101001001010;
            sine_reg0   <= 36'sb101001011010000100011000011001011111;
        end
        14341: begin
            cosine_reg0 <= 36'sb10110101010111011011100011110000110;
            sine_reg0   <= 36'sb101001011010100111111111000100111001;
        end
        14342: begin
            cosine_reg0 <= 36'sb10110101011011110111010011011000110;
            sine_reg0   <= 36'sb101001011011001011100110101000000010;
        end
        14343: begin
            cosine_reg0 <= 36'sb10110101100000010010111100000001000;
            sine_reg0   <= 36'sb101001011011101111001111000010110111;
        end
        14344: begin
            cosine_reg0 <= 36'sb10110101100100101110011101101001011;
            sine_reg0   <= 36'sb101001011100010010111000010101011000;
        end
        14345: begin
            cosine_reg0 <= 36'sb10110101101001001001111000010001111;
            sine_reg0   <= 36'sb101001011100110110100010011111100100;
        end
        14346: begin
            cosine_reg0 <= 36'sb10110101101101100101001011111010000;
            sine_reg0   <= 36'sb101001011101011010001101100001011000;
        end
        14347: begin
            cosine_reg0 <= 36'sb10110101110010000000011000100001111;
            sine_reg0   <= 36'sb101001011101111101111001011010110011;
        end
        14348: begin
            cosine_reg0 <= 36'sb10110101110110011011011110001001010;
            sine_reg0   <= 36'sb101001011110100001100110001011110101;
        end
        14349: begin
            cosine_reg0 <= 36'sb10110101111010110110011100101111111;
            sine_reg0   <= 36'sb101001011111000101010011110100011011;
        end
        14350: begin
            cosine_reg0 <= 36'sb10110101111111010001010100010101110;
            sine_reg0   <= 36'sb101001011111101001000010010100100101;
        end
        14351: begin
            cosine_reg0 <= 36'sb10110110000011101100000100111010011;
            sine_reg0   <= 36'sb101001100000001100110001101100010000;
        end
        14352: begin
            cosine_reg0 <= 36'sb10110110001000000110101110011110000;
            sine_reg0   <= 36'sb101001100000110000100001111011011100;
        end
        14353: begin
            cosine_reg0 <= 36'sb10110110001100100001010001000000001;
            sine_reg0   <= 36'sb101001100001010100010011000010001000;
        end
        14354: begin
            cosine_reg0 <= 36'sb10110110010000111011101100100000110;
            sine_reg0   <= 36'sb101001100001111000000101000000010001;
        end
        14355: begin
            cosine_reg0 <= 36'sb10110110010101010110000000111111101;
            sine_reg0   <= 36'sb101001100010011011110111110101110110;
        end
        14356: begin
            cosine_reg0 <= 36'sb10110110011001110000001110011100101;
            sine_reg0   <= 36'sb101001100010111111101011100010110111;
        end
        14357: begin
            cosine_reg0 <= 36'sb10110110011110001010010100110111100;
            sine_reg0   <= 36'sb101001100011100011100000000111010001;
        end
        14358: begin
            cosine_reg0 <= 36'sb10110110100010100100010100010000010;
            sine_reg0   <= 36'sb101001100100000111010101100011000100;
        end
        14359: begin
            cosine_reg0 <= 36'sb10110110100110111110001100100110100;
            sine_reg0   <= 36'sb101001100100101011001011110110001101;
        end
        14360: begin
            cosine_reg0 <= 36'sb10110110101011010111111101111010010;
            sine_reg0   <= 36'sb101001100101001111000011000000101100;
        end
        14361: begin
            cosine_reg0 <= 36'sb10110110101111110001101000001011010;
            sine_reg0   <= 36'sb101001100101110010111011000010011111;
        end
        14362: begin
            cosine_reg0 <= 36'sb10110110110100001011001011011001011;
            sine_reg0   <= 36'sb101001100110010110110011111011100101;
        end
        14363: begin
            cosine_reg0 <= 36'sb10110110111000100100100111100100011;
            sine_reg0   <= 36'sb101001100110111010101101101011111100;
        end
        14364: begin
            cosine_reg0 <= 36'sb10110110111100111101111100101100001;
            sine_reg0   <= 36'sb101001100111011110101000010011100011;
        end
        14365: begin
            cosine_reg0 <= 36'sb10110111000001010111001010110000011;
            sine_reg0   <= 36'sb101001101000000010100011110010011001;
        end
        14366: begin
            cosine_reg0 <= 36'sb10110111000101110000010001110001001;
            sine_reg0   <= 36'sb101001101000100110100000001000011100;
        end
        14367: begin
            cosine_reg0 <= 36'sb10110111001010001001010001101110001;
            sine_reg0   <= 36'sb101001101001001010011101010101101011;
        end
        14368: begin
            cosine_reg0 <= 36'sb10110111001110100010001010100111010;
            sine_reg0   <= 36'sb101001101001101110011011011010000101;
        end
        14369: begin
            cosine_reg0 <= 36'sb10110111010010111010111100011100010;
            sine_reg0   <= 36'sb101001101010010010011010010101100111;
        end
        14370: begin
            cosine_reg0 <= 36'sb10110111010111010011100111001100111;
            sine_reg0   <= 36'sb101001101010110110011010001000010001;
        end
        14371: begin
            cosine_reg0 <= 36'sb10110111011011101100001010111001010;
            sine_reg0   <= 36'sb101001101011011010011010110010000001;
        end
        14372: begin
            cosine_reg0 <= 36'sb10110111100000000100100111100000111;
            sine_reg0   <= 36'sb101001101011111110011100010010110111;
        end
        14373: begin
            cosine_reg0 <= 36'sb10110111100100011100111101000011110;
            sine_reg0   <= 36'sb101001101100100010011110101010101111;
        end
        14374: begin
            cosine_reg0 <= 36'sb10110111101000110101001011100001110;
            sine_reg0   <= 36'sb101001101101000110100001111001101010;
        end
        14375: begin
            cosine_reg0 <= 36'sb10110111101101001101010010111010101;
            sine_reg0   <= 36'sb101001101101101010100101111111100110;
        end
        14376: begin
            cosine_reg0 <= 36'sb10110111110001100101010011001110010;
            sine_reg0   <= 36'sb101001101110001110101010111100100001;
        end
        14377: begin
            cosine_reg0 <= 36'sb10110111110101111101001100011100011;
            sine_reg0   <= 36'sb101001101110110010110000110000011010;
        end
        14378: begin
            cosine_reg0 <= 36'sb10110111111010010100111110100100111;
            sine_reg0   <= 36'sb101001101111010110110111011011001111;
        end
        14379: begin
            cosine_reg0 <= 36'sb10110111111110101100101001100111101;
            sine_reg0   <= 36'sb101001101111111010111110111101000000;
        end
        14380: begin
            cosine_reg0 <= 36'sb10111000000011000100001101100100011;
            sine_reg0   <= 36'sb101001110000011111000111010101101010;
        end
        14381: begin
            cosine_reg0 <= 36'sb10111000000111011011101010011011000;
            sine_reg0   <= 36'sb101001110001000011010000100101001101;
        end
        14382: begin
            cosine_reg0 <= 36'sb10111000001011110011000000001011011;
            sine_reg0   <= 36'sb101001110001100111011010101011100111;
        end
        14383: begin
            cosine_reg0 <= 36'sb10111000010000001010001110110101011;
            sine_reg0   <= 36'sb101001110010001011100101101000110110;
        end
        14384: begin
            cosine_reg0 <= 36'sb10111000010100100001010110011000101;
            sine_reg0   <= 36'sb101001110010101111110001011100111010;
        end
        14385: begin
            cosine_reg0 <= 36'sb10111000011000111000010110110101001;
            sine_reg0   <= 36'sb101001110011010011111110000111110000;
        end
        14386: begin
            cosine_reg0 <= 36'sb10111000011101001111010000001010101;
            sine_reg0   <= 36'sb101001110011111000001011101001011000;
        end
        14387: begin
            cosine_reg0 <= 36'sb10111000100001100110000010011001001;
            sine_reg0   <= 36'sb101001110100011100011010000001110000;
        end
        14388: begin
            cosine_reg0 <= 36'sb10111000100101111100101101100000010;
            sine_reg0   <= 36'sb101001110101000000101001010000110110;
        end
        14389: begin
            cosine_reg0 <= 36'sb10111000101010010011010001011111111;
            sine_reg0   <= 36'sb101001110101100100111001010110101010;
        end
        14390: begin
            cosine_reg0 <= 36'sb10111000101110101001101110010111111;
            sine_reg0   <= 36'sb101001110110001001001010010011001001;
        end
        14391: begin
            cosine_reg0 <= 36'sb10111000110011000000000100001000001;
            sine_reg0   <= 36'sb101001110110101101011100000110010011;
        end
        14392: begin
            cosine_reg0 <= 36'sb10111000110111010110010010110000011;
            sine_reg0   <= 36'sb101001110111010001101110110000000110;
        end
        14393: begin
            cosine_reg0 <= 36'sb10111000111011101100011010010000100;
            sine_reg0   <= 36'sb101001110111110110000010010000100000;
        end
        14394: begin
            cosine_reg0 <= 36'sb10111001000000000010011010101000010;
            sine_reg0   <= 36'sb101001111000011010010110100111100001;
        end
        14395: begin
            cosine_reg0 <= 36'sb10111001000100011000010011110111101;
            sine_reg0   <= 36'sb101001111000111110101011110101000110;
        end
        14396: begin
            cosine_reg0 <= 36'sb10111001001000101110000101111110011;
            sine_reg0   <= 36'sb101001111001100011000001111001001111;
        end
        14397: begin
            cosine_reg0 <= 36'sb10111001001101000011110000111100010;
            sine_reg0   <= 36'sb101001111010000111011000110011111010;
        end
        14398: begin
            cosine_reg0 <= 36'sb10111001010001011001010100110001001;
            sine_reg0   <= 36'sb101001111010101011110000100101000110;
        end
        14399: begin
            cosine_reg0 <= 36'sb10111001010101101110110001011100111;
            sine_reg0   <= 36'sb101001111011010000001001001100110001;
        end
        14400: begin
            cosine_reg0 <= 36'sb10111001011010000100000110111111011;
            sine_reg0   <= 36'sb101001111011110100100010101010111001;
        end
        14401: begin
            cosine_reg0 <= 36'sb10111001011110011001010101011000011;
            sine_reg0   <= 36'sb101001111100011000111100111111011110;
        end
        14402: begin
            cosine_reg0 <= 36'sb10111001100010101110011100100111110;
            sine_reg0   <= 36'sb101001111100111101011000001010011110;
        end
        14403: begin
            cosine_reg0 <= 36'sb10111001100111000011011100101101011;
            sine_reg0   <= 36'sb101001111101100001110100001011111000;
        end
        14404: begin
            cosine_reg0 <= 36'sb10111001101011011000010101101000111;
            sine_reg0   <= 36'sb101001111110000110010001000011101010;
        end
        14405: begin
            cosine_reg0 <= 36'sb10111001101111101101000111011010011;
            sine_reg0   <= 36'sb101001111110101010101110110001110011;
        end
        14406: begin
            cosine_reg0 <= 36'sb10111001110100000001110010000001100;
            sine_reg0   <= 36'sb101001111111001111001101010110010001;
        end
        14407: begin
            cosine_reg0 <= 36'sb10111001111000010110010101011110001;
            sine_reg0   <= 36'sb101001111111110011101100110001000011;
        end
        14408: begin
            cosine_reg0 <= 36'sb10111001111100101010110001110000001;
            sine_reg0   <= 36'sb101010000000011000001101000010000111;
        end
        14409: begin
            cosine_reg0 <= 36'sb10111010000000111111000110110111011;
            sine_reg0   <= 36'sb101010000000111100101110001001011101;
        end
        14410: begin
            cosine_reg0 <= 36'sb10111010000101010011010100110011101;
            sine_reg0   <= 36'sb101010000001100001010000000111000011;
        end
        14411: begin
            cosine_reg0 <= 36'sb10111010001001100111011011100100101;
            sine_reg0   <= 36'sb101010000010000101110010111010110111;
        end
        14412: begin
            cosine_reg0 <= 36'sb10111010001101111011011011001010100;
            sine_reg0   <= 36'sb101010000010101010010110100100110111;
        end
        14413: begin
            cosine_reg0 <= 36'sb10111010010010001111010011100100110;
            sine_reg0   <= 36'sb101010000011001110111011000101000100;
        end
        14414: begin
            cosine_reg0 <= 36'sb10111010010110100011000100110011011;
            sine_reg0   <= 36'sb101010000011110011100000011011011010;
        end
        14415: begin
            cosine_reg0 <= 36'sb10111010011010110110101110110110010;
            sine_reg0   <= 36'sb101010000100011000000110100111111001;
        end
        14416: begin
            cosine_reg0 <= 36'sb10111010011111001010010001101101001;
            sine_reg0   <= 36'sb101010000100111100101101101010100000;
        end
        14417: begin
            cosine_reg0 <= 36'sb10111010100011011101101101011000000;
            sine_reg0   <= 36'sb101010000101100001010101100011001100;
        end
        14418: begin
            cosine_reg0 <= 36'sb10111010100111110001000001110110011;
            sine_reg0   <= 36'sb101010000110000101111110010001111101;
        end
        14419: begin
            cosine_reg0 <= 36'sb10111010101100000100001111001000011;
            sine_reg0   <= 36'sb101010000110101010100111110110110001;
        end
        14420: begin
            cosine_reg0 <= 36'sb10111010110000010111010101001101110;
            sine_reg0   <= 36'sb101010000111001111010010010001100111;
        end
        14421: begin
            cosine_reg0 <= 36'sb10111010110100101010010100000110010;
            sine_reg0   <= 36'sb101010000111110011111101100010011100;
        end
        14422: begin
            cosine_reg0 <= 36'sb10111010111000111101001011110001111;
            sine_reg0   <= 36'sb101010001000011000101001101001010001;
        end
        14423: begin
            cosine_reg0 <= 36'sb10111010111101001111111100010000010;
            sine_reg0   <= 36'sb101010001000111101010110100110000011;
        end
        14424: begin
            cosine_reg0 <= 36'sb10111011000001100010100101100001011;
            sine_reg0   <= 36'sb101010001001100010000100011000110001;
        end
        14425: begin
            cosine_reg0 <= 36'sb10111011000101110101000111100101001;
            sine_reg0   <= 36'sb101010001010000110110011000001011010;
        end
        14426: begin
            cosine_reg0 <= 36'sb10111011001010000111100010011011001;
            sine_reg0   <= 36'sb101010001010101011100010011111111100;
        end
        14427: begin
            cosine_reg0 <= 36'sb10111011001110011001110110000011011;
            sine_reg0   <= 36'sb101010001011010000010010110100010101;
        end
        14428: begin
            cosine_reg0 <= 36'sb10111011010010101100000010011101110;
            sine_reg0   <= 36'sb101010001011110101000011111110100101;
        end
        14429: begin
            cosine_reg0 <= 36'sb10111011010110111110000111101001111;
            sine_reg0   <= 36'sb101010001100011001110101111110101010;
        end
        14430: begin
            cosine_reg0 <= 36'sb10111011011011010000000101100111110;
            sine_reg0   <= 36'sb101010001100111110101000110100100010;
        end
        14431: begin
            cosine_reg0 <= 36'sb10111011011111100001111100010111010;
            sine_reg0   <= 36'sb101010001101100011011100100000001100;
        end
        14432: begin
            cosine_reg0 <= 36'sb10111011100011110011101011111000000;
            sine_reg0   <= 36'sb101010001110001000010001000001100111;
        end
        14433: begin
            cosine_reg0 <= 36'sb10111011101000000101010100001010000;
            sine_reg0   <= 36'sb101010001110101101000110011000110010;
        end
        14434: begin
            cosine_reg0 <= 36'sb10111011101100010110110101001101001;
            sine_reg0   <= 36'sb101010001111010001111100100101101010;
        end
        14435: begin
            cosine_reg0 <= 36'sb10111011110000101000001111000001001;
            sine_reg0   <= 36'sb101010001111110110110011101000001110;
        end
        14436: begin
            cosine_reg0 <= 36'sb10111011110100111001100001100101110;
            sine_reg0   <= 36'sb101010010000011011101011100000011110;
        end
        14437: begin
            cosine_reg0 <= 36'sb10111011111001001010101100111011000;
            sine_reg0   <= 36'sb101010010001000000100100001110010111;
        end
        14438: begin
            cosine_reg0 <= 36'sb10111011111101011011110001000000101;
            sine_reg0   <= 36'sb101010010001100101011101110001111000;
        end
        14439: begin
            cosine_reg0 <= 36'sb10111100000001101100101101110110100;
            sine_reg0   <= 36'sb101010010010001010011000001011000000;
        end
        14440: begin
            cosine_reg0 <= 36'sb10111100000101111101100011011100011;
            sine_reg0   <= 36'sb101010010010101111010011011001101101;
        end
        14441: begin
            cosine_reg0 <= 36'sb10111100001010001110010001110010010;
            sine_reg0   <= 36'sb101010010011010100001111011101111110;
        end
        14442: begin
            cosine_reg0 <= 36'sb10111100001110011110111000110111110;
            sine_reg0   <= 36'sb101010010011111001001100010111110001;
        end
        14443: begin
            cosine_reg0 <= 36'sb10111100010010101111011000101101000;
            sine_reg0   <= 36'sb101010010100011110001010000111000110;
        end
        14444: begin
            cosine_reg0 <= 36'sb10111100010110111111110001010001100;
            sine_reg0   <= 36'sb101010010101000011001000101011111010;
        end
        14445: begin
            cosine_reg0 <= 36'sb10111100011011010000000010100101010;
            sine_reg0   <= 36'sb101010010101101000001000000110001100;
        end
        14446: begin
            cosine_reg0 <= 36'sb10111100011111100000001100101000001;
            sine_reg0   <= 36'sb101010010110001101001000010101111011;
        end
        14447: begin
            cosine_reg0 <= 36'sb10111100100011110000001111011001111;
            sine_reg0   <= 36'sb101010010110110010001001011011000101;
        end
        14448: begin
            cosine_reg0 <= 36'sb10111100101000000000001010111010011;
            sine_reg0   <= 36'sb101010010111010111001011010101101001;
        end
        14449: begin
            cosine_reg0 <= 36'sb10111100101100001111111111001001100;
            sine_reg0   <= 36'sb101010010111111100001110000101100110;
        end
        14450: begin
            cosine_reg0 <= 36'sb10111100110000011111101100000111000;
            sine_reg0   <= 36'sb101010011000100001010001101010111010;
        end
        14451: begin
            cosine_reg0 <= 36'sb10111100110100101111010001110010110;
            sine_reg0   <= 36'sb101010011001000110010110000101100011;
        end
        14452: begin
            cosine_reg0 <= 36'sb10111100111000111110110000001100101;
            sine_reg0   <= 36'sb101010011001101011011011010101100000;
        end
        14453: begin
            cosine_reg0 <= 36'sb10111100111101001110000111010100100;
            sine_reg0   <= 36'sb101010011010010000100001011010110000;
        end
        14454: begin
            cosine_reg0 <= 36'sb10111101000001011101010111001010001;
            sine_reg0   <= 36'sb101010011010110101101000010101010010;
        end
        14455: begin
            cosine_reg0 <= 36'sb10111101000101101100011111101101010;
            sine_reg0   <= 36'sb101010011011011010110000000101000011;
        end
        14456: begin
            cosine_reg0 <= 36'sb10111101001001111011100000111101111;
            sine_reg0   <= 36'sb101010011011111111111000101010000011;
        end
        14457: begin
            cosine_reg0 <= 36'sb10111101001110001010011010111011110;
            sine_reg0   <= 36'sb101010011100100101000010000100010000;
        end
        14458: begin
            cosine_reg0 <= 36'sb10111101010010011001001101100110111;
            sine_reg0   <= 36'sb101010011101001010001100010011101000;
        end
        14459: begin
            cosine_reg0 <= 36'sb10111101010110100111111000111110110;
            sine_reg0   <= 36'sb101010011101101111010111011000001011;
        end
        14460: begin
            cosine_reg0 <= 36'sb10111101011010110110011101000011100;
            sine_reg0   <= 36'sb101010011110010100100011010001110110;
        end
        14461: begin
            cosine_reg0 <= 36'sb10111101011111000100111001110101000;
            sine_reg0   <= 36'sb101010011110111001110000000000101000;
        end
        14462: begin
            cosine_reg0 <= 36'sb10111101100011010011001111010010110;
            sine_reg0   <= 36'sb101010011111011110111101100100100001;
        end
        14463: begin
            cosine_reg0 <= 36'sb10111101100111100001011101011101000;
            sine_reg0   <= 36'sb101010100000000100001011111101011110;
        end
        14464: begin
            cosine_reg0 <= 36'sb10111101101011101111100100010011010;
            sine_reg0   <= 36'sb101010100000101001011011001011011101;
        end
        14465: begin
            cosine_reg0 <= 36'sb10111101101111111101100011110101100;
            sine_reg0   <= 36'sb101010100001001110101011001110011111;
        end
        14466: begin
            cosine_reg0 <= 36'sb10111101110100001011011100000011101;
            sine_reg0   <= 36'sb101010100001110011111100000110100000;
        end
        14467: begin
            cosine_reg0 <= 36'sb10111101111000011001001100111101010;
            sine_reg0   <= 36'sb101010100010011001001101110011100000;
        end
        14468: begin
            cosine_reg0 <= 36'sb10111101111100100110110110100010100;
            sine_reg0   <= 36'sb101010100010111110100000010101011110;
        end
        14469: begin
            cosine_reg0 <= 36'sb10111110000000110100011000110011000;
            sine_reg0   <= 36'sb101010100011100011110011101100010111;
        end
        14470: begin
            cosine_reg0 <= 36'sb10111110000101000001110011101110110;
            sine_reg0   <= 36'sb101010100100001001000111111000001010;
        end
        14471: begin
            cosine_reg0 <= 36'sb10111110001001001111000111010101100;
            sine_reg0   <= 36'sb101010100100101110011100111000110111;
        end
        14472: begin
            cosine_reg0 <= 36'sb10111110001101011100010011100111000;
            sine_reg0   <= 36'sb101010100101010011110010101110011011;
        end
        14473: begin
            cosine_reg0 <= 36'sb10111110010001101001011000100011010;
            sine_reg0   <= 36'sb101010100101111001001001011000110101;
        end
        14474: begin
            cosine_reg0 <= 36'sb10111110010101110110010110001001111;
            sine_reg0   <= 36'sb101010100110011110100000111000000011;
        end
        14475: begin
            cosine_reg0 <= 36'sb10111110011010000011001100011011000;
            sine_reg0   <= 36'sb101010100111000011111001001100000101;
        end
        14476: begin
            cosine_reg0 <= 36'sb10111110011110001111111011010110010;
            sine_reg0   <= 36'sb101010100111101001010010010100111001;
        end
        14477: begin
            cosine_reg0 <= 36'sb10111110100010011100100010111011101;
            sine_reg0   <= 36'sb101010101000001110101100010010011100;
        end
        14478: begin
            cosine_reg0 <= 36'sb10111110100110101001000011001010110;
            sine_reg0   <= 36'sb101010101000110100000111000100101111;
        end
        14479: begin
            cosine_reg0 <= 36'sb10111110101010110101011100000011101;
            sine_reg0   <= 36'sb101010101001011001100010101011101111;
        end
        14480: begin
            cosine_reg0 <= 36'sb10111110101111000001101101100110000;
            sine_reg0   <= 36'sb101010101001111110111111000111011011;
        end
        14481: begin
            cosine_reg0 <= 36'sb10111110110011001101110111110001110;
            sine_reg0   <= 36'sb101010101010100100011100010111110001;
        end
        14482: begin
            cosine_reg0 <= 36'sb10111110110111011001111010100110110;
            sine_reg0   <= 36'sb101010101011001001111010011100110001;
        end
        14483: begin
            cosine_reg0 <= 36'sb10111110111011100101110110000100111;
            sine_reg0   <= 36'sb101010101011101111011001010110011000;
        end
        14484: begin
            cosine_reg0 <= 36'sb10111110111111110001101010001011111;
            sine_reg0   <= 36'sb101010101100010100111001000100100101;
        end
        14485: begin
            cosine_reg0 <= 36'sb10111111000011111101010110111011100;
            sine_reg0   <= 36'sb101010101100111010011001100111010111;
        end
        14486: begin
            cosine_reg0 <= 36'sb10111111001000001000111100010011110;
            sine_reg0   <= 36'sb101010101101011111111010111110101101;
        end
        14487: begin
            cosine_reg0 <= 36'sb10111111001100010100011010010100100;
            sine_reg0   <= 36'sb101010101110000101011101001010100100;
        end
        14488: begin
            cosine_reg0 <= 36'sb10111111010000011111110000111101011;
            sine_reg0   <= 36'sb101010101110101011000000001010111011;
        end
        14489: begin
            cosine_reg0 <= 36'sb10111111010100101011000000001110100;
            sine_reg0   <= 36'sb101010101111010000100011111111110010;
        end
        14490: begin
            cosine_reg0 <= 36'sb10111111011000110110001000000111011;
            sine_reg0   <= 36'sb101010101111110110001000101001000110;
        end
        14491: begin
            cosine_reg0 <= 36'sb10111111011101000001001000101000001;
            sine_reg0   <= 36'sb101010110000011011101110000110110110;
        end
        14492: begin
            cosine_reg0 <= 36'sb10111111100001001100000001110000100;
            sine_reg0   <= 36'sb101010110001000001010100011001000000;
        end
        14493: begin
            cosine_reg0 <= 36'sb10111111100101010110110011100000010;
            sine_reg0   <= 36'sb101010110001100110111011011111100100;
        end
        14494: begin
            cosine_reg0 <= 36'sb10111111101001100001011101110111010;
            sine_reg0   <= 36'sb101010110010001100100011011010100000;
        end
        14495: begin
            cosine_reg0 <= 36'sb10111111101101101100000000110101100;
            sine_reg0   <= 36'sb101010110010110010001100001001110001;
        end
        14496: begin
            cosine_reg0 <= 36'sb10111111110001110110011100011010101;
            sine_reg0   <= 36'sb101010110011010111110101101101011000;
        end
        14497: begin
            cosine_reg0 <= 36'sb10111111110110000000110000100110101;
            sine_reg0   <= 36'sb101010110011111101100000000101010010;
        end
        14498: begin
            cosine_reg0 <= 36'sb10111111111010001010111101011001010;
            sine_reg0   <= 36'sb101010110100100011001011010001011101;
        end
        14499: begin
            cosine_reg0 <= 36'sb10111111111110010101000010110010010;
            sine_reg0   <= 36'sb101010110101001000110111010001111010;
        end
        14500: begin
            cosine_reg0 <= 36'sb11000000000010011111000000110001101;
            sine_reg0   <= 36'sb101010110101101110100100000110100101;
        end
        14501: begin
            cosine_reg0 <= 36'sb11000000000110101000110111010111010;
            sine_reg0   <= 36'sb101010110110010100010001101111011101;
        end
        14502: begin
            cosine_reg0 <= 36'sb11000000001010110010100110100010111;
            sine_reg0   <= 36'sb101010110110111010000000001100100010;
        end
        14503: begin
            cosine_reg0 <= 36'sb11000000001110111100001110010100010;
            sine_reg0   <= 36'sb101010110111011111101111011101110010;
        end
        14504: begin
            cosine_reg0 <= 36'sb11000000010011000101101110101011011;
            sine_reg0   <= 36'sb101010111000000101011111100011001010;
        end
        14505: begin
            cosine_reg0 <= 36'sb11000000010111001111000111101000000;
            sine_reg0   <= 36'sb101010111000101011010000011100101011;
        end
        14506: begin
            cosine_reg0 <= 36'sb11000000011011011000011001001010000;
            sine_reg0   <= 36'sb101010111001010001000010001010010001;
        end
        14507: begin
            cosine_reg0 <= 36'sb11000000011111100001100011010001001;
            sine_reg0   <= 36'sb101010111001110110110100101011111100;
        end
        14508: begin
            cosine_reg0 <= 36'sb11000000100011101010100101111101011;
            sine_reg0   <= 36'sb101010111010011100101000000001101011;
        end
        14509: begin
            cosine_reg0 <= 36'sb11000000100111110011100001001110100;
            sine_reg0   <= 36'sb101010111011000010011100001011011100;
        end
        14510: begin
            cosine_reg0 <= 36'sb11000000101011111100010101000100011;
            sine_reg0   <= 36'sb101010111011101000010001001001001101;
        end
        14511: begin
            cosine_reg0 <= 36'sb11000000110000000101000001011110110;
            sine_reg0   <= 36'sb101010111100001110000110111010111101;
        end
        14512: begin
            cosine_reg0 <= 36'sb11000000110100001101100110011101101;
            sine_reg0   <= 36'sb101010111100110011111101100000101010;
        end
        14513: begin
            cosine_reg0 <= 36'sb11000000111000010110000100000000101;
            sine_reg0   <= 36'sb101010111101011001110100111010010100;
        end
        14514: begin
            cosine_reg0 <= 36'sb11000000111100011110011010000111110;
            sine_reg0   <= 36'sb101010111101111111101101000111111000;
        end
        14515: begin
            cosine_reg0 <= 36'sb11000001000000100110101000110010111;
            sine_reg0   <= 36'sb101010111110100101100110001001010101;
        end
        14516: begin
            cosine_reg0 <= 36'sb11000001000100101110110000000001110;
            sine_reg0   <= 36'sb101010111111001011011111111110101010;
        end
        14517: begin
            cosine_reg0 <= 36'sb11000001001000110110101111110100001;
            sine_reg0   <= 36'sb101010111111110001011010100111110101;
        end
        14518: begin
            cosine_reg0 <= 36'sb11000001001100111110101000001010000;
            sine_reg0   <= 36'sb101011000000010111010110000100110101;
        end
        14519: begin
            cosine_reg0 <= 36'sb11000001010001000110011001000011010;
            sine_reg0   <= 36'sb101011000000111101010010010101101000;
        end
        14520: begin
            cosine_reg0 <= 36'sb11000001010101001110000010011111101;
            sine_reg0   <= 36'sb101011000001100011001111011010001101;
        end
        14521: begin
            cosine_reg0 <= 36'sb11000001011001010101100100011110111;
            sine_reg0   <= 36'sb101011000010001001001101010010100011;
        end
        14522: begin
            cosine_reg0 <= 36'sb11000001011101011100111111000001000;
            sine_reg0   <= 36'sb101011000010101111001011111110100111;
        end
        14523: begin
            cosine_reg0 <= 36'sb11000001100001100100010010000101110;
            sine_reg0   <= 36'sb101011000011010101001011011110011001;
        end
        14524: begin
            cosine_reg0 <= 36'sb11000001100101101011011101101101000;
            sine_reg0   <= 36'sb101011000011111011001011110001110111;
        end
        14525: begin
            cosine_reg0 <= 36'sb11000001101001110010100001110110101;
            sine_reg0   <= 36'sb101011000100100001001100111000111111;
        end
        14526: begin
            cosine_reg0 <= 36'sb11000001101101111001011110100010011;
            sine_reg0   <= 36'sb101011000101000111001110110011110000;
        end
        14527: begin
            cosine_reg0 <= 36'sb11000001110010000000010011110000010;
            sine_reg0   <= 36'sb101011000101101101010001100010001001;
        end
        14528: begin
            cosine_reg0 <= 36'sb11000001110110000111000001011111111;
            sine_reg0   <= 36'sb101011000110010011010101000100001000;
        end
        14529: begin
            cosine_reg0 <= 36'sb11000001111010001101100111110001010;
            sine_reg0   <= 36'sb101011000110111001011001011001101011;
        end
        14530: begin
            cosine_reg0 <= 36'sb11000001111110010100000110100100010;
            sine_reg0   <= 36'sb101011000111011111011110100010110010;
        end
        14531: begin
            cosine_reg0 <= 36'sb11000010000010011010011101111000100;
            sine_reg0   <= 36'sb101011001000000101100100011111011010;
        end
        14532: begin
            cosine_reg0 <= 36'sb11000010000110100000101101101110000;
            sine_reg0   <= 36'sb101011001000101011101011001111100011;
        end
        14533: begin
            cosine_reg0 <= 36'sb11000010001010100110110110000100101;
            sine_reg0   <= 36'sb101011001001010001110010110011001010;
        end
        14534: begin
            cosine_reg0 <= 36'sb11000010001110101100110110111100010;
            sine_reg0   <= 36'sb101011001001110111111011001010001111;
        end
        14535: begin
            cosine_reg0 <= 36'sb11000010010010110010110000010100100;
            sine_reg0   <= 36'sb101011001010011110000100010100110000;
        end
        14536: begin
            cosine_reg0 <= 36'sb11000010010110111000100010001101011;
            sine_reg0   <= 36'sb101011001011000100001110010010101010;
        end
        14537: begin
            cosine_reg0 <= 36'sb11000010011010111110001100100110110;
            sine_reg0   <= 36'sb101011001011101010011001000011111110;
        end
        14538: begin
            cosine_reg0 <= 36'sb11000010011111000011101111100000011;
            sine_reg0   <= 36'sb101011001100010000100100101000101001;
        end
        14539: begin
            cosine_reg0 <= 36'sb11000010100011001001001010111010001;
            sine_reg0   <= 36'sb101011001100110110110001000000101011;
        end
        14540: begin
            cosine_reg0 <= 36'sb11000010100111001110011110110011110;
            sine_reg0   <= 36'sb101011001101011100111110001100000000;
        end
        14541: begin
            cosine_reg0 <= 36'sb11000010101011010011101011001101011;
            sine_reg0   <= 36'sb101011001110000011001100001010101001;
        end
        14542: begin
            cosine_reg0 <= 36'sb11000010101111011000110000000110100;
            sine_reg0   <= 36'sb101011001110101001011010111100100011;
        end
        14543: begin
            cosine_reg0 <= 36'sb11000010110011011101101101011111001;
            sine_reg0   <= 36'sb101011001111001111101010100001101101;
        end
        14544: begin
            cosine_reg0 <= 36'sb11000010110111100010100011010111010;
            sine_reg0   <= 36'sb101011001111110101111010111010000110;
        end
        14545: begin
            cosine_reg0 <= 36'sb11000010111011100111010001101110011;
            sine_reg0   <= 36'sb101011010000011100001100000101101011;
        end
        14546: begin
            cosine_reg0 <= 36'sb11000010111111101011111000100100101;
            sine_reg0   <= 36'sb101011010001000010011110000100011101;
        end
        14547: begin
            cosine_reg0 <= 36'sb11000011000011110000010111111001110;
            sine_reg0   <= 36'sb101011010001101000110000110110011000;
        end
        14548: begin
            cosine_reg0 <= 36'sb11000011000111110100101111101101100;
            sine_reg0   <= 36'sb101011010010001111000100011011011101;
        end
        14549: begin
            cosine_reg0 <= 36'sb11000011001011111000111111111111111;
            sine_reg0   <= 36'sb101011010010110101011000110011101000;
        end
        14550: begin
            cosine_reg0 <= 36'sb11000011001111111101001000110000101;
            sine_reg0   <= 36'sb101011010011011011101101111110111001;
        end
        14551: begin
            cosine_reg0 <= 36'sb11000011010100000001001001111111101;
            sine_reg0   <= 36'sb101011010100000010000011111101001111;
        end
        14552: begin
            cosine_reg0 <= 36'sb11000011011000000101000011101100110;
            sine_reg0   <= 36'sb101011010100101000011010101110100111;
        end
        14553: begin
            cosine_reg0 <= 36'sb11000011011100001000110101110111110;
            sine_reg0   <= 36'sb101011010101001110110010010011000000;
        end
        14554: begin
            cosine_reg0 <= 36'sb11000011100000001100100000100000100;
            sine_reg0   <= 36'sb101011010101110101001010101010011010;
        end
        14555: begin
            cosine_reg0 <= 36'sb11000011100100010000000011100111000;
            sine_reg0   <= 36'sb101011010110011011100011110100110001;
        end
        14556: begin
            cosine_reg0 <= 36'sb11000011101000010011011111001010110;
            sine_reg0   <= 36'sb101011010111000001111101110010000101;
        end
        14557: begin
            cosine_reg0 <= 36'sb11000011101100010110110011001100000;
            sine_reg0   <= 36'sb101011010111101000011000100010010101;
        end
        14558: begin
            cosine_reg0 <= 36'sb11000011110000011001111111101010010;
            sine_reg0   <= 36'sb101011011000001110110100000101011111;
        end
        14559: begin
            cosine_reg0 <= 36'sb11000011110100011101000100100101101;
            sine_reg0   <= 36'sb101011011000110101010000011011100001;
        end
        14560: begin
            cosine_reg0 <= 36'sb11000011111000100000000001111101110;
            sine_reg0   <= 36'sb101011011001011011101101100100011010;
        end
        14561: begin
            cosine_reg0 <= 36'sb11000011111100100010110111110010100;
            sine_reg0   <= 36'sb101011011010000010001011100000001000;
        end
        14562: begin
            cosine_reg0 <= 36'sb11000100000000100101100110000011111;
            sine_reg0   <= 36'sb101011011010101000101010001110101011;
        end
        14563: begin
            cosine_reg0 <= 36'sb11000100000100101000001100110001101;
            sine_reg0   <= 36'sb101011011011001111001001101111111111;
        end
        14564: begin
            cosine_reg0 <= 36'sb11000100001000101010101011111011100;
            sine_reg0   <= 36'sb101011011011110101101010000100000101;
        end
        14565: begin
            cosine_reg0 <= 36'sb11000100001100101101000011100001100;
            sine_reg0   <= 36'sb101011011100011100001011001010111010;
        end
        14566: begin
            cosine_reg0 <= 36'sb11000100010000101111010011100011011;
            sine_reg0   <= 36'sb101011011101000010101101000100011110;
        end
        14567: begin
            cosine_reg0 <= 36'sb11000100010100110001011100000001000;
            sine_reg0   <= 36'sb101011011101101001001111110000101110;
        end
        14568: begin
            cosine_reg0 <= 36'sb11000100011000110011011100111010001;
            sine_reg0   <= 36'sb101011011110001111110011001111101000;
        end
        14569: begin
            cosine_reg0 <= 36'sb11000100011100110101010110001110110;
            sine_reg0   <= 36'sb101011011110110110010111100001001101;
        end
        14570: begin
            cosine_reg0 <= 36'sb11000100100000110111000111111110110;
            sine_reg0   <= 36'sb101011011111011100111100100101011001;
        end
        14571: begin
            cosine_reg0 <= 36'sb11000100100100111000110010001001110;
            sine_reg0   <= 36'sb101011100000000011100010011100001101;
        end
        14572: begin
            cosine_reg0 <= 36'sb11000100101000111010010100101111110;
            sine_reg0   <= 36'sb101011100000101010001001000101100101;
        end
        14573: begin
            cosine_reg0 <= 36'sb11000100101100111011101111110000101;
            sine_reg0   <= 36'sb101011100001010000110000100001100000;
        end
        14574: begin
            cosine_reg0 <= 36'sb11000100110000111101000011001100000;
            sine_reg0   <= 36'sb101011100001110111011000101111111110;
        end
        14575: begin
            cosine_reg0 <= 36'sb11000100110100111110001111000010000;
            sine_reg0   <= 36'sb101011100010011110000001110000111101;
        end
        14576: begin
            cosine_reg0 <= 36'sb11000100111000111111010011010010011;
            sine_reg0   <= 36'sb101011100011000100101011100100011011;
        end
        14577: begin
            cosine_reg0 <= 36'sb11000100111101000000001111111100111;
            sine_reg0   <= 36'sb101011100011101011010110001010010110;
        end
        14578: begin
            cosine_reg0 <= 36'sb11000101000001000001000101000001011;
            sine_reg0   <= 36'sb101011100100010010000001100010101101;
        end
        14579: begin
            cosine_reg0 <= 36'sb11000101000101000001110010011111111;
            sine_reg0   <= 36'sb101011100100111000101101101101011111;
        end
        14580: begin
            cosine_reg0 <= 36'sb11000101001001000010011000011000000;
            sine_reg0   <= 36'sb101011100101011111011010101010101011;
        end
        14581: begin
            cosine_reg0 <= 36'sb11000101001101000010110110101001110;
            sine_reg0   <= 36'sb101011100110000110001000011010001110;
        end
        14582: begin
            cosine_reg0 <= 36'sb11000101010001000011001101010100111;
            sine_reg0   <= 36'sb101011100110101100110110111100000111;
        end
        14583: begin
            cosine_reg0 <= 36'sb11000101010101000011011100011001011;
            sine_reg0   <= 36'sb101011100111010011100110010000010101;
        end
        14584: begin
            cosine_reg0 <= 36'sb11000101011001000011100011110110111;
            sine_reg0   <= 36'sb101011100111111010010110010110110110;
        end
        14585: begin
            cosine_reg0 <= 36'sb11000101011101000011100011101101011;
            sine_reg0   <= 36'sb101011101000100001000111001111101001;
        end
        14586: begin
            cosine_reg0 <= 36'sb11000101100001000011011011111100101;
            sine_reg0   <= 36'sb101011101001000111111000111010101100;
        end
        14587: begin
            cosine_reg0 <= 36'sb11000101100101000011001100100100100;
            sine_reg0   <= 36'sb101011101001101110101011010111111101;
        end
        14588: begin
            cosine_reg0 <= 36'sb11000101101001000010110101100101000;
            sine_reg0   <= 36'sb101011101010010101011110100111011100;
        end
        14589: begin
            cosine_reg0 <= 36'sb11000101101101000010010110111101110;
            sine_reg0   <= 36'sb101011101010111100010010101001000111;
        end
        14590: begin
            cosine_reg0 <= 36'sb11000101110001000001110000101110110;
            sine_reg0   <= 36'sb101011101011100011000111011100111100;
        end
        14591: begin
            cosine_reg0 <= 36'sb11000101110101000001000010110111110;
            sine_reg0   <= 36'sb101011101100001001111101000010111001;
        end
        14592: begin
            cosine_reg0 <= 36'sb11000101111001000000001101011000100;
            sine_reg0   <= 36'sb101011101100110000110011011010111110;
        end
        14593: begin
            cosine_reg0 <= 36'sb11000101111100111111010000010001001;
            sine_reg0   <= 36'sb101011101101010111101010100101001001;
        end
        14594: begin
            cosine_reg0 <= 36'sb11000110000000111110001011100001010;
            sine_reg0   <= 36'sb101011101101111110100010100001011000;
        end
        14595: begin
            cosine_reg0 <= 36'sb11000110000100111100111111001000111;
            sine_reg0   <= 36'sb101011101110100101011011001111101001;
        end
        14596: begin
            cosine_reg0 <= 36'sb11000110001000111011101011000111110;
            sine_reg0   <= 36'sb101011101111001100010100101111111100;
        end
        14597: begin
            cosine_reg0 <= 36'sb11000110001100111010001111011101101;
            sine_reg0   <= 36'sb101011101111110011001111000010001111;
        end
        14598: begin
            cosine_reg0 <= 36'sb11000110010000111000101100001010101;
            sine_reg0   <= 36'sb101011110000011010001010000110100000;
        end
        14599: begin
            cosine_reg0 <= 36'sb11000110010100110111000001001110010;
            sine_reg0   <= 36'sb101011110001000001000101111100101101;
        end
        14600: begin
            cosine_reg0 <= 36'sb11000110011000110101001110101000101;
            sine_reg0   <= 36'sb101011110001101000000010100100110110;
        end
        14601: begin
            cosine_reg0 <= 36'sb11000110011100110011010100011001100;
            sine_reg0   <= 36'sb101011110010001110111111111110111001;
        end
        14602: begin
            cosine_reg0 <= 36'sb11000110100000110001010010100000110;
            sine_reg0   <= 36'sb101011110010110101111110001010110011;
        end
        14603: begin
            cosine_reg0 <= 36'sb11000110100100101111001000111110001;
            sine_reg0   <= 36'sb101011110011011100111101001000100101;
        end
        14604: begin
            cosine_reg0 <= 36'sb11000110101000101100110111110001100;
            sine_reg0   <= 36'sb101011110100000011111100111000001100;
        end
        14605: begin
            cosine_reg0 <= 36'sb11000110101100101010011110111010111;
            sine_reg0   <= 36'sb101011110100101010111101011001100110;
        end
        14606: begin
            cosine_reg0 <= 36'sb11000110110000100111111110011001111;
            sine_reg0   <= 36'sb101011110101010001111110101100110011;
        end
        14607: begin
            cosine_reg0 <= 36'sb11000110110100100101010110001110100;
            sine_reg0   <= 36'sb101011110101111001000000110001110000;
        end
        14608: begin
            cosine_reg0 <= 36'sb11000110111000100010100110011000101;
            sine_reg0   <= 36'sb101011110110100000000011101000011101;
        end
        14609: begin
            cosine_reg0 <= 36'sb11000110111100011111101110111000000;
            sine_reg0   <= 36'sb101011110111000111000111010000110111;
        end
        14610: begin
            cosine_reg0 <= 36'sb11000111000000011100101111101100011;
            sine_reg0   <= 36'sb101011110111101110001011101010111110;
        end
        14611: begin
            cosine_reg0 <= 36'sb11000111000100011001101000110101111;
            sine_reg0   <= 36'sb101011111000010101010000110110101111;
        end
        14612: begin
            cosine_reg0 <= 36'sb11000111001000010110011010010100001;
            sine_reg0   <= 36'sb101011111000111100010110110100001010;
        end
        14613: begin
            cosine_reg0 <= 36'sb11000111001100010011000100000111000;
            sine_reg0   <= 36'sb101011111001100011011101100011001100;
        end
        14614: begin
            cosine_reg0 <= 36'sb11000111010000001111100110001110011;
            sine_reg0   <= 36'sb101011111010001010100101000011110100;
        end
        14615: begin
            cosine_reg0 <= 36'sb11000111010100001100000000101010001;
            sine_reg0   <= 36'sb101011111010110001101101010110000001;
        end
        14616: begin
            cosine_reg0 <= 36'sb11000111011000001000010011011010001;
            sine_reg0   <= 36'sb101011111011011000110110011001110001;
        end
        14617: begin
            cosine_reg0 <= 36'sb11000111011100000100011110011110010;
            sine_reg0   <= 36'sb101011111100000000000000001111000011;
        end
        14618: begin
            cosine_reg0 <= 36'sb11000111100000000000100001110110001;
            sine_reg0   <= 36'sb101011111100100111001010110101110101;
        end
        14619: begin
            cosine_reg0 <= 36'sb11000111100011111100011101100001111;
            sine_reg0   <= 36'sb101011111101001110010110001110000110;
        end
        14620: begin
            cosine_reg0 <= 36'sb11000111100111111000010001100001001;
            sine_reg0   <= 36'sb101011111101110101100010010111110011;
        end
        14621: begin
            cosine_reg0 <= 36'sb11000111101011110011111101110011111;
            sine_reg0   <= 36'sb101011111110011100101111010010111101;
        end
        14622: begin
            cosine_reg0 <= 36'sb11000111101111101111100010011010000;
            sine_reg0   <= 36'sb101011111111000011111100111111100000;
        end
        14623: begin
            cosine_reg0 <= 36'sb11000111110011101010111111010011010;
            sine_reg0   <= 36'sb101011111111101011001011011101011100;
        end
        14624: begin
            cosine_reg0 <= 36'sb11000111110111100110010100011111011;
            sine_reg0   <= 36'sb101100000000010010011010101100101111;
        end
        14625: begin
            cosine_reg0 <= 36'sb11000111111011100001100001111110011;
            sine_reg0   <= 36'sb101100000000111001101010101101011000;
        end
        14626: begin
            cosine_reg0 <= 36'sb11000111111111011100100111110000001;
            sine_reg0   <= 36'sb101100000001100000111011011111010101;
        end
        14627: begin
            cosine_reg0 <= 36'sb11001000000011010111100101110100011;
            sine_reg0   <= 36'sb101100000010001000001101000010100100;
        end
        14628: begin
            cosine_reg0 <= 36'sb11001000000111010010011100001011001;
            sine_reg0   <= 36'sb101100000010101111011111010111000100;
        end
        14629: begin
            cosine_reg0 <= 36'sb11001000001011001101001010110100000;
            sine_reg0   <= 36'sb101100000011010110110010011100110100;
        end
        14630: begin
            cosine_reg0 <= 36'sb11001000001111000111110001101111000;
            sine_reg0   <= 36'sb101100000011111110000110010011110010;
        end
        14631: begin
            cosine_reg0 <= 36'sb11001000010011000010010000111011111;
            sine_reg0   <= 36'sb101100000100100101011010111011111100;
        end
        14632: begin
            cosine_reg0 <= 36'sb11001000010110111100101000011010101;
            sine_reg0   <= 36'sb101100000101001100110000010101010001;
        end
        14633: begin
            cosine_reg0 <= 36'sb11001000011010110110111000001011000;
            sine_reg0   <= 36'sb101100000101110100000110011111110000;
        end
        14634: begin
            cosine_reg0 <= 36'sb11001000011110110001000000001100111;
            sine_reg0   <= 36'sb101100000110011011011101011011010110;
        end
        14635: begin
            cosine_reg0 <= 36'sb11001000100010101011000000100000000;
            sine_reg0   <= 36'sb101100000111000010110101001000000011;
        end
        14636: begin
            cosine_reg0 <= 36'sb11001000100110100100111001000100011;
            sine_reg0   <= 36'sb101100000111101010001101100101110101;
        end
        14637: begin
            cosine_reg0 <= 36'sb11001000101010011110101001111001110;
            sine_reg0   <= 36'sb101100001000010001100110110100101010;
        end
        14638: begin
            cosine_reg0 <= 36'sb11001000101110011000010011000000000;
            sine_reg0   <= 36'sb101100001000111001000000110100100010;
        end
        14639: begin
            cosine_reg0 <= 36'sb11001000110010010001110100010111000;
            sine_reg0   <= 36'sb101100001001100000011011100101011001;
        end
        14640: begin
            cosine_reg0 <= 36'sb11001000110110001011001101111110100;
            sine_reg0   <= 36'sb101100001010000111110111000111001111;
        end
        14641: begin
            cosine_reg0 <= 36'sb11001000111010000100011111110110100;
            sine_reg0   <= 36'sb101100001010101111010011011010000011;
        end
        14642: begin
            cosine_reg0 <= 36'sb11001000111101111101101001111110111;
            sine_reg0   <= 36'sb101100001011010110110000011101110010;
        end
        14643: begin
            cosine_reg0 <= 36'sb11001001000001110110101100010111010;
            sine_reg0   <= 36'sb101100001011111110001110010010011100;
        end
        14644: begin
            cosine_reg0 <= 36'sb11001001000101101111100110111111101;
            sine_reg0   <= 36'sb101100001100100101101100110111111110;
        end
        14645: begin
            cosine_reg0 <= 36'sb11001001001001101000011001110111111;
            sine_reg0   <= 36'sb101100001101001101001100001110011000;
        end
        14646: begin
            cosine_reg0 <= 36'sb11001001001101100001000100111111110;
            sine_reg0   <= 36'sb101100001101110100101100010101100111;
        end
        14647: begin
            cosine_reg0 <= 36'sb11001001010001011001101000010111010;
            sine_reg0   <= 36'sb101100001110011100001101001101101010;
        end
        14648: begin
            cosine_reg0 <= 36'sb11001001010101010010000011111110001;
            sine_reg0   <= 36'sb101100001111000011101110110110100000;
        end
        14649: begin
            cosine_reg0 <= 36'sb11001001011001001010010111110100001;
            sine_reg0   <= 36'sb101100001111101011010001010000000111;
        end
        14650: begin
            cosine_reg0 <= 36'sb11001001011101000010100011111001010;
            sine_reg0   <= 36'sb101100010000010010110100011010011110;
        end
        14651: begin
            cosine_reg0 <= 36'sb11001001100000111010101000001101011;
            sine_reg0   <= 36'sb101100010000111010011000010101100011;
        end
        14652: begin
            cosine_reg0 <= 36'sb11001001100100110010100100110000010;
            sine_reg0   <= 36'sb101100010001100001111101000001010100;
        end
        14653: begin
            cosine_reg0 <= 36'sb11001001101000101010011001100001110;
            sine_reg0   <= 36'sb101100010010001001100010011101110001;
        end
        14654: begin
            cosine_reg0 <= 36'sb11001001101100100010000110100001101;
            sine_reg0   <= 36'sb101100010010110001001000101010110110;
        end
        14655: begin
            cosine_reg0 <= 36'sb11001001110000011001101011110000000;
            sine_reg0   <= 36'sb101100010011011000101111101000100100;
        end
        14656: begin
            cosine_reg0 <= 36'sb11001001110100010001001001001100100;
            sine_reg0   <= 36'sb101100010100000000010111010110111001;
        end
        14657: begin
            cosine_reg0 <= 36'sb11001001111000001000011110110111000;
            sine_reg0   <= 36'sb101100010100100111111111110101110010;
        end
        14658: begin
            cosine_reg0 <= 36'sb11001001111011111111101100101111011;
            sine_reg0   <= 36'sb101100010101001111101001000101001110;
        end
        14659: begin
            cosine_reg0 <= 36'sb11001001111111110110110010110101101;
            sine_reg0   <= 36'sb101100010101110111010011000101001101;
        end
        14660: begin
            cosine_reg0 <= 36'sb11001010000011101101110001001001011;
            sine_reg0   <= 36'sb101100010110011110111101110101101011;
        end
        14661: begin
            cosine_reg0 <= 36'sb11001010000111100100100111101010100;
            sine_reg0   <= 36'sb101100010111000110101001010110101001;
        end
        14662: begin
            cosine_reg0 <= 36'sb11001010001011011011010110011001000;
            sine_reg0   <= 36'sb101100010111101110010101101000000100;
        end
        14663: begin
            cosine_reg0 <= 36'sb11001010001111010001111101010100101;
            sine_reg0   <= 36'sb101100011000010110000010101001111010;
        end
        14664: begin
            cosine_reg0 <= 36'sb11001010010011001000011100011101010;
            sine_reg0   <= 36'sb101100011000111101110000011100001011;
        end
        14665: begin
            cosine_reg0 <= 36'sb11001010010110111110110011110010110;
            sine_reg0   <= 36'sb101100011001100101011110111110110100;
        end
        14666: begin
            cosine_reg0 <= 36'sb11001010011010110101000011010100111;
            sine_reg0   <= 36'sb101100011010001101001110010001110101;
        end
        14667: begin
            cosine_reg0 <= 36'sb11001010011110101011001011000011101;
            sine_reg0   <= 36'sb101100011010110100111110010101001011;
        end
        14668: begin
            cosine_reg0 <= 36'sb11001010100010100001001010111110110;
            sine_reg0   <= 36'sb101100011011011100101111001000110101;
        end
        14669: begin
            cosine_reg0 <= 36'sb11001010100110010111000011000110001;
            sine_reg0   <= 36'sb101100011100000100100000101100110010;
        end
        14670: begin
            cosine_reg0 <= 36'sb11001010101010001100110011011001101;
            sine_reg0   <= 36'sb101100011100101100010011000001000000;
        end
        14671: begin
            cosine_reg0 <= 36'sb11001010101110000010011011111001001;
            sine_reg0   <= 36'sb101100011101010100000110000101011101;
        end
        14672: begin
            cosine_reg0 <= 36'sb11001010110001110111111100100100011;
            sine_reg0   <= 36'sb101100011101111011111001111010001001;
        end
        14673: begin
            cosine_reg0 <= 36'sb11001010110101101101010101011011010;
            sine_reg0   <= 36'sb101100011110100011101110011111000000;
        end
        14674: begin
            cosine_reg0 <= 36'sb11001010111001100010100110011101110;
            sine_reg0   <= 36'sb101100011111001011100011110100000011;
        end
        14675: begin
            cosine_reg0 <= 36'sb11001010111101010111101111101011100;
            sine_reg0   <= 36'sb101100011111110011011001111001001111;
        end
        14676: begin
            cosine_reg0 <= 36'sb11001011000001001100110001000100100;
            sine_reg0   <= 36'sb101100100000011011010000101110100010;
        end
        14677: begin
            cosine_reg0 <= 36'sb11001011000101000001101010101000101;
            sine_reg0   <= 36'sb101100100001000011001000010011111100;
        end
        14678: begin
            cosine_reg0 <= 36'sb11001011001000110110011100010111101;
            sine_reg0   <= 36'sb101100100001101011000000101001011011;
        end
        14679: begin
            cosine_reg0 <= 36'sb11001011001100101011000110010001011;
            sine_reg0   <= 36'sb101100100010010010111001101110111101;
        end
        14680: begin
            cosine_reg0 <= 36'sb11001011010000011111101000010101111;
            sine_reg0   <= 36'sb101100100010111010110011100100100000;
        end
        14681: begin
            cosine_reg0 <= 36'sb11001011010100010100000010100100110;
            sine_reg0   <= 36'sb101100100011100010101110001010000100;
        end
        14682: begin
            cosine_reg0 <= 36'sb11001011011000001000010100111110000;
            sine_reg0   <= 36'sb101100100100001010101001011111100110;
        end
        14683: begin
            cosine_reg0 <= 36'sb11001011011011111100011111100001011;
            sine_reg0   <= 36'sb101100100100110010100101100101000101;
        end
        14684: begin
            cosine_reg0 <= 36'sb11001011011111110000100010001110111;
            sine_reg0   <= 36'sb101100100101011010100010011010100000;
        end
        14685: begin
            cosine_reg0 <= 36'sb11001011100011100100011101000110010;
            sine_reg0   <= 36'sb101100100110000010011111111111110101;
        end
        14686: begin
            cosine_reg0 <= 36'sb11001011100111011000010000000111010;
            sine_reg0   <= 36'sb101100100110101010011110010101000010;
        end
        14687: begin
            cosine_reg0 <= 36'sb11001011101011001011111011010010000;
            sine_reg0   <= 36'sb101100100111010010011101011010000110;
        end
        14688: begin
            cosine_reg0 <= 36'sb11001011101110111111011110100110001;
            sine_reg0   <= 36'sb101100100111111010011101001110111111;
        end
        14689: begin
            cosine_reg0 <= 36'sb11001011110010110010111010000011101;
            sine_reg0   <= 36'sb101100101000100010011101110011101100;
        end
        14690: begin
            cosine_reg0 <= 36'sb11001011110110100110001101101010010;
            sine_reg0   <= 36'sb101100101001001010011111001000001011;
        end
        14691: begin
            cosine_reg0 <= 36'sb11001011111010011001011001011001111;
            sine_reg0   <= 36'sb101100101001110010100001001100011011;
        end
        14692: begin
            cosine_reg0 <= 36'sb11001011111110001100011101010010011;
            sine_reg0   <= 36'sb101100101010011010100100000000011011;
        end
        14693: begin
            cosine_reg0 <= 36'sb11001100000001111111011001010011101;
            sine_reg0   <= 36'sb101100101011000010100111100100001000;
        end
        14694: begin
            cosine_reg0 <= 36'sb11001100000101110010001101011101011;
            sine_reg0   <= 36'sb101100101011101010101011110111100000;
        end
        14695: begin
            cosine_reg0 <= 36'sb11001100001001100100111001101111101;
            sine_reg0   <= 36'sb101100101100010010110000111010100100;
        end
        14696: begin
            cosine_reg0 <= 36'sb11001100001101010111011110001010001;
            sine_reg0   <= 36'sb101100101100111010110110101101010000;
        end
        14697: begin
            cosine_reg0 <= 36'sb11001100010001001001111010101100110;
            sine_reg0   <= 36'sb101100101101100010111101001111100100;
        end
        14698: begin
            cosine_reg0 <= 36'sb11001100010100111100001111010111011;
            sine_reg0   <= 36'sb101100101110001011000100100001011110;
        end
        14699: begin
            cosine_reg0 <= 36'sb11001100011000101110011100001001110;
            sine_reg0   <= 36'sb101100101110110011001100100010111100;
        end
        14700: begin
            cosine_reg0 <= 36'sb11001100011100100000100001000100000;
            sine_reg0   <= 36'sb101100101111011011010101010011111101;
        end
        14701: begin
            cosine_reg0 <= 36'sb11001100100000010010011110000101101;
            sine_reg0   <= 36'sb101100110000000011011110110100011111;
        end
        14702: begin
            cosine_reg0 <= 36'sb11001100100100000100010011001110110;
            sine_reg0   <= 36'sb101100110000101011101001000100100001;
        end
        14703: begin
            cosine_reg0 <= 36'sb11001100100111110110000000011111001;
            sine_reg0   <= 36'sb101100110001010011110100000100000001;
        end
        14704: begin
            cosine_reg0 <= 36'sb11001100101011100111100101110110101;
            sine_reg0   <= 36'sb101100110001111011111111110010111101;
        end
        14705: begin
            cosine_reg0 <= 36'sb11001100101111011001000011010101001;
            sine_reg0   <= 36'sb101100110010100100001100010001010101;
        end
        14706: begin
            cosine_reg0 <= 36'sb11001100110011001010011000111010011;
            sine_reg0   <= 36'sb101100110011001100011001011111000110;
        end
        14707: begin
            cosine_reg0 <= 36'sb11001100110110111011100110100110011;
            sine_reg0   <= 36'sb101100110011110100100111011100001111;
        end
        14708: begin
            cosine_reg0 <= 36'sb11001100111010101100101100011000111;
            sine_reg0   <= 36'sb101100110100011100110110001000101111;
        end
        14709: begin
            cosine_reg0 <= 36'sb11001100111110011101101010010001110;
            sine_reg0   <= 36'sb101100110101000101000101100100100011;
        end
        14710: begin
            cosine_reg0 <= 36'sb11001101000010001110100000010000111;
            sine_reg0   <= 36'sb101100110101101101010101101111101011;
        end
        14711: begin
            cosine_reg0 <= 36'sb11001101000101111111001110010110001;
            sine_reg0   <= 36'sb101100110110010101100110101010000101;
        end
        14712: begin
            cosine_reg0 <= 36'sb11001101001001101111110100100001010;
            sine_reg0   <= 36'sb101100110110111101111000010011101110;
        end
        14713: begin
            cosine_reg0 <= 36'sb11001101001101100000010010110010010;
            sine_reg0   <= 36'sb101100110111100110001010101100100110;
        end
        14714: begin
            cosine_reg0 <= 36'sb11001101010001010000101001001000111;
            sine_reg0   <= 36'sb101100111000001110011101110100101100;
        end
        14715: begin
            cosine_reg0 <= 36'sb11001101010101000000110111100101000;
            sine_reg0   <= 36'sb101100111000110110110001101011111101;
        end
        14716: begin
            cosine_reg0 <= 36'sb11001101011000110000111110000110100;
            sine_reg0   <= 36'sb101100111001011111000110010010011000;
        end
        14717: begin
            cosine_reg0 <= 36'sb11001101011100100000111100101101010;
            sine_reg0   <= 36'sb101100111010000111011011100111111011;
        end
        14718: begin
            cosine_reg0 <= 36'sb11001101100000010000110011011001001;
            sine_reg0   <= 36'sb101100111010101111110001101100100101;
        end
        14719: begin
            cosine_reg0 <= 36'sb11001101100100000000100010001001111;
            sine_reg0   <= 36'sb101100111011011000001000100000010101;
        end
        14720: begin
            cosine_reg0 <= 36'sb11001101100111110000001000111111100;
            sine_reg0   <= 36'sb101100111100000000100000000011001000;
        end
        14721: begin
            cosine_reg0 <= 36'sb11001101101011011111100111111001110;
            sine_reg0   <= 36'sb101100111100101000111000010100111110;
        end
        14722: begin
            cosine_reg0 <= 36'sb11001101101111001110111110111000100;
            sine_reg0   <= 36'sb101100111101010001010001010101110100;
        end
        14723: begin
            cosine_reg0 <= 36'sb11001101110010111110001101111011100;
            sine_reg0   <= 36'sb101100111101111001101011000101101001;
        end
        14724: begin
            cosine_reg0 <= 36'sb11001101110110101101010101000010111;
            sine_reg0   <= 36'sb101100111110100010000101100100011100;
        end
        14725: begin
            cosine_reg0 <= 36'sb11001101111010011100010100001110010;
            sine_reg0   <= 36'sb101100111111001010100000110010001011;
        end
        14726: begin
            cosine_reg0 <= 36'sb11001101111110001011001011011101101;
            sine_reg0   <= 36'sb101100111111110010111100101110110100;
        end
        14727: begin
            cosine_reg0 <= 36'sb11001110000001111001111010110000101;
            sine_reg0   <= 36'sb101101000000011011011001011010010110;
        end
        14728: begin
            cosine_reg0 <= 36'sb11001110000101101000100010000111011;
            sine_reg0   <= 36'sb101101000001000011110110110100110000;
        end
        14729: begin
            cosine_reg0 <= 36'sb11001110001001010111000001100001101;
            sine_reg0   <= 36'sb101101000001101100010100111101111111;
        end
        14730: begin
            cosine_reg0 <= 36'sb11001110001101000101011000111111010;
            sine_reg0   <= 36'sb101101000010010100110011110110000010;
        end
        14731: begin
            cosine_reg0 <= 36'sb11001110010000110011101000100000000;
            sine_reg0   <= 36'sb101101000010111101010011011100111000;
        end
        14732: begin
            cosine_reg0 <= 36'sb11001110010100100001110000000011111;
            sine_reg0   <= 36'sb101101000011100101110011110010011111;
        end
        14733: begin
            cosine_reg0 <= 36'sb11001110011000001111101111101010110;
            sine_reg0   <= 36'sb101101000100001110010100110110110101;
        end
        14734: begin
            cosine_reg0 <= 36'sb11001110011011111101100111010100010;
            sine_reg0   <= 36'sb101101000100110110110110101001111010;
        end
        14735: begin
            cosine_reg0 <= 36'sb11001110011111101011010111000000100;
            sine_reg0   <= 36'sb101101000101011111011001001011101011;
        end
        14736: begin
            cosine_reg0 <= 36'sb11001110100011011000111110101111010;
            sine_reg0   <= 36'sb101101000110000111111100011100000110;
        end
        14737: begin
            cosine_reg0 <= 36'sb11001110100111000110011110100000010;
            sine_reg0   <= 36'sb101101000110110000100000011011001011;
        end
        14738: begin
            cosine_reg0 <= 36'sb11001110101010110011110110010011100;
            sine_reg0   <= 36'sb101101000111011001000101001000111000;
        end
        14739: begin
            cosine_reg0 <= 36'sb11001110101110100001000110001000111;
            sine_reg0   <= 36'sb101101001000000001101010100101001010;
        end
        14740: begin
            cosine_reg0 <= 36'sb11001110110010001110001110000000001;
            sine_reg0   <= 36'sb101101001000101010010000110000000010;
        end
        14741: begin
            cosine_reg0 <= 36'sb11001110110101111011001101111001001;
            sine_reg0   <= 36'sb101101001001010010110111101001011100;
        end
        14742: begin
            cosine_reg0 <= 36'sb11001110111001101000000101110011111;
            sine_reg0   <= 36'sb101101001001111011011111010001011000;
        end
        14743: begin
            cosine_reg0 <= 36'sb11001110111101010100110101110000000;
            sine_reg0   <= 36'sb101101001010100100000111100111110011;
        end
        14744: begin
            cosine_reg0 <= 36'sb11001111000001000001011101101101100;
            sine_reg0   <= 36'sb101101001011001100110000101100101101;
        end
        14745: begin
            cosine_reg0 <= 36'sb11001111000100101101111101101100010;
            sine_reg0   <= 36'sb101101001011110101011010100000000011;
        end
        14746: begin
            cosine_reg0 <= 36'sb11001111001000011010010101101100000;
            sine_reg0   <= 36'sb101101001100011110000101000001110101;
        end
        14747: begin
            cosine_reg0 <= 36'sb11001111001100000110100101101100110;
            sine_reg0   <= 36'sb101101001101000110110000010010000000;
        end
        14748: begin
            cosine_reg0 <= 36'sb11001111001111110010101101101110010;
            sine_reg0   <= 36'sb101101001101101111011100010000100100;
        end
        14749: begin
            cosine_reg0 <= 36'sb11001111010011011110101101110000011;
            sine_reg0   <= 36'sb101101001110011000001000111101011110;
        end
        14750: begin
            cosine_reg0 <= 36'sb11001111010111001010100101110011000;
            sine_reg0   <= 36'sb101101001111000000110110011000101100;
        end
        14751: begin
            cosine_reg0 <= 36'sb11001111011010110110010101110110000;
            sine_reg0   <= 36'sb101101001111101001100100100010001110;
        end
        14752: begin
            cosine_reg0 <= 36'sb11001111011110100001111101111001010;
            sine_reg0   <= 36'sb101101010000010010010011011010000010;
        end
        14753: begin
            cosine_reg0 <= 36'sb11001111100010001101011101111100100;
            sine_reg0   <= 36'sb101101010000111011000011000000000110;
        end
        14754: begin
            cosine_reg0 <= 36'sb11001111100101111000110101111111101;
            sine_reg0   <= 36'sb101101010001100011110011010100011000;
        end
        14755: begin
            cosine_reg0 <= 36'sb11001111101001100100000110000010101;
            sine_reg0   <= 36'sb101101010010001100100100010110111000;
        end
        14756: begin
            cosine_reg0 <= 36'sb11001111101101001111001110000101010;
            sine_reg0   <= 36'sb101101010010110101010110000111100011;
        end
        14757: begin
            cosine_reg0 <= 36'sb11001111110000111010001110000111011;
            sine_reg0   <= 36'sb101101010011011110001000100110011000;
        end
        14758: begin
            cosine_reg0 <= 36'sb11001111110100100101000110001000111;
            sine_reg0   <= 36'sb101101010100000110111011110011010101;
        end
        14759: begin
            cosine_reg0 <= 36'sb11001111111000001111110110001001101;
            sine_reg0   <= 36'sb101101010100101111101111101110011001;
        end
        14760: begin
            cosine_reg0 <= 36'sb11001111111011111010011110001001100;
            sine_reg0   <= 36'sb101101010101011000100100010111100010;
        end
        14761: begin
            cosine_reg0 <= 36'sb11001111111111100100111110001000001;
            sine_reg0   <= 36'sb101101010110000001011001101110101111;
        end
        14762: begin
            cosine_reg0 <= 36'sb11010000000011001111010110000101110;
            sine_reg0   <= 36'sb101101010110101010001111110011111101;
        end
        14763: begin
            cosine_reg0 <= 36'sb11010000000110111001100110000001111;
            sine_reg0   <= 36'sb101101010111010011000110100111001100;
        end
        14764: begin
            cosine_reg0 <= 36'sb11010000001010100011101101111100101;
            sine_reg0   <= 36'sb101101010111111011111110001000011011;
        end
        14765: begin
            cosine_reg0 <= 36'sb11010000001110001101101101110101101;
            sine_reg0   <= 36'sb101101011000100100110110010111100110;
        end
        14766: begin
            cosine_reg0 <= 36'sb11010000010001110111100101101101000;
            sine_reg0   <= 36'sb101101011001001101101111010100101101;
        end
        14767: begin
            cosine_reg0 <= 36'sb11010000010101100001010101100010011;
            sine_reg0   <= 36'sb101101011001110110101000111111101110;
        end
        14768: begin
            cosine_reg0 <= 36'sb11010000011001001010111101010101110;
            sine_reg0   <= 36'sb101101011010011111100011011000101000;
        end
        14769: begin
            cosine_reg0 <= 36'sb11010000011100110100011101000110111;
            sine_reg0   <= 36'sb101101011011001000011110011111011001;
        end
        14770: begin
            cosine_reg0 <= 36'sb11010000100000011101110100110101110;
            sine_reg0   <= 36'sb101101011011110001011010010011111111;
        end
        14771: begin
            cosine_reg0 <= 36'sb11010000100100000111000100100010001;
            sine_reg0   <= 36'sb101101011100011010010110110110011001;
        end
        14772: begin
            cosine_reg0 <= 36'sb11010000100111110000001100001011111;
            sine_reg0   <= 36'sb101101011101000011010100000110100101;
        end
        14773: begin
            cosine_reg0 <= 36'sb11010000101011011001001011110010111;
            sine_reg0   <= 36'sb101101011101101100010010000100100010;
        end
        14774: begin
            cosine_reg0 <= 36'sb11010000101111000010000011010111000;
            sine_reg0   <= 36'sb101101011110010101010000110000001110;
        end
        14775: begin
            cosine_reg0 <= 36'sb11010000110010101010110010111000000;
            sine_reg0   <= 36'sb101101011110111110010000001001101000;
        end
        14776: begin
            cosine_reg0 <= 36'sb11010000110110010011011010010101111;
            sine_reg0   <= 36'sb101101011111100111010000010000101101;
        end
        14777: begin
            cosine_reg0 <= 36'sb11010000111001111011111001110000100;
            sine_reg0   <= 36'sb101101100000010000010001000101011101;
        end
        14778: begin
            cosine_reg0 <= 36'sb11010000111101100100010001000111101;
            sine_reg0   <= 36'sb101101100000111001010010100111110110;
        end
        14779: begin
            cosine_reg0 <= 36'sb11010001000001001100100000011011001;
            sine_reg0   <= 36'sb101101100001100010010100110111110110;
        end
        14780: begin
            cosine_reg0 <= 36'sb11010001000100110100100111101011000;
            sine_reg0   <= 36'sb101101100010001011010111110101011011;
        end
        14781: begin
            cosine_reg0 <= 36'sb11010001001000011100100110110110111;
            sine_reg0   <= 36'sb101101100010110100011011100000100101;
        end
        14782: begin
            cosine_reg0 <= 36'sb11010001001100000100011101111110111;
            sine_reg0   <= 36'sb101101100011011101011111111001010000;
        end
        14783: begin
            cosine_reg0 <= 36'sb11010001001111101100001101000010101;
            sine_reg0   <= 36'sb101101100100000110100100111111011101;
        end
        14784: begin
            cosine_reg0 <= 36'sb11010001010011010011110100000010001;
            sine_reg0   <= 36'sb101101100100101111101010110011001001;
        end
        14785: begin
            cosine_reg0 <= 36'sb11010001010110111011010010111101001;
            sine_reg0   <= 36'sb101101100101011000110001010100010011;
        end
        14786: begin
            cosine_reg0 <= 36'sb11010001011010100010101001110011101;
            sine_reg0   <= 36'sb101101100110000001111000100010111001;
        end
        14787: begin
            cosine_reg0 <= 36'sb11010001011110001001111000100101011;
            sine_reg0   <= 36'sb101101100110101011000000011110111001;
        end
        14788: begin
            cosine_reg0 <= 36'sb11010001100001110000111111010010010;
            sine_reg0   <= 36'sb101101100111010100001001001000010011;
        end
        14789: begin
            cosine_reg0 <= 36'sb11010001100101010111111101111010010;
            sine_reg0   <= 36'sb101101100111111101010010011111000011;
        end
        14790: begin
            cosine_reg0 <= 36'sb11010001101000111110110100011101000;
            sine_reg0   <= 36'sb101101101000100110011100100011001010;
        end
        14791: begin
            cosine_reg0 <= 36'sb11010001101100100101100010111010100;
            sine_reg0   <= 36'sb101101101001001111100111010100100100;
        end
        14792: begin
            cosine_reg0 <= 36'sb11010001110000001100001001010010101;
            sine_reg0   <= 36'sb101101101001111000110010110011010010;
        end
        14793: begin
            cosine_reg0 <= 36'sb11010001110011110010100111100101010;
            sine_reg0   <= 36'sb101101101010100001111110111111010000;
        end
        14794: begin
            cosine_reg0 <= 36'sb11010001110111011000111101110010001;
            sine_reg0   <= 36'sb101101101011001011001011111000011110;
        end
        14795: begin
            cosine_reg0 <= 36'sb11010001111010111111001011111001010;
            sine_reg0   <= 36'sb101101101011110100011001011110111001;
        end
        14796: begin
            cosine_reg0 <= 36'sb11010001111110100101010001111010011;
            sine_reg0   <= 36'sb101101101100011101100111110010100001;
        end
        14797: begin
            cosine_reg0 <= 36'sb11010010000010001011001111110101011;
            sine_reg0   <= 36'sb101101101101000110110110110011010011;
        end
        14798: begin
            cosine_reg0 <= 36'sb11010010000101110001000101101010001;
            sine_reg0   <= 36'sb101101101101110000000110100001001111;
        end
        14799: begin
            cosine_reg0 <= 36'sb11010010001001010110110011011000100;
            sine_reg0   <= 36'sb101101101110011001010110111100010010;
        end
        14800: begin
            cosine_reg0 <= 36'sb11010010001100111100011001000000100;
            sine_reg0   <= 36'sb101101101111000010101000000100011010;
        end
        14801: begin
            cosine_reg0 <= 36'sb11010010010000100001110110100001101;
            sine_reg0   <= 36'sb101101101111101011111001111001100111;
        end
        14802: begin
            cosine_reg0 <= 36'sb11010010010100000111001011111100001;
            sine_reg0   <= 36'sb101101110000010101001100011011110111;
        end
        14803: begin
            cosine_reg0 <= 36'sb11010010010111101100011001001111101;
            sine_reg0   <= 36'sb101101110000111110011111101011001000;
        end
        14804: begin
            cosine_reg0 <= 36'sb11010010011011010001011110011100001;
            sine_reg0   <= 36'sb101101110001100111110011100111011001;
        end
        14805: begin
            cosine_reg0 <= 36'sb11010010011110110110011011100001011;
            sine_reg0   <= 36'sb101101110010010001001000010000100111;
        end
        14806: begin
            cosine_reg0 <= 36'sb11010010100010011011010000011111010;
            sine_reg0   <= 36'sb101101110010111010011101100110110010;
        end
        14807: begin
            cosine_reg0 <= 36'sb11010010100101111111111101010101101;
            sine_reg0   <= 36'sb101101110011100011110011101001110111;
        end
        14808: begin
            cosine_reg0 <= 36'sb11010010101001100100100010000100011;
            sine_reg0   <= 36'sb101101110100001101001010011001110110;
        end
        14809: begin
            cosine_reg0 <= 36'sb11010010101101001000111110101011100;
            sine_reg0   <= 36'sb101101110100110110100001110110101100;
        end
        14810: begin
            cosine_reg0 <= 36'sb11010010110000101101010011001010101;
            sine_reg0   <= 36'sb101101110101011111111010000000011000;
        end
        14811: begin
            cosine_reg0 <= 36'sb11010010110100010001011111100001110;
            sine_reg0   <= 36'sb101101110110001001010010110110111000;
        end
        14812: begin
            cosine_reg0 <= 36'sb11010010110111110101100011110000101;
            sine_reg0   <= 36'sb101101110110110010101100011010001011;
        end
        14813: begin
            cosine_reg0 <= 36'sb11010010111011011001011111110111010;
            sine_reg0   <= 36'sb101101110111011100000110101010010000;
        end
        14814: begin
            cosine_reg0 <= 36'sb11010010111110111101010011110101100;
            sine_reg0   <= 36'sb101101111000000101100001100111000011;
        end
        14815: begin
            cosine_reg0 <= 36'sb11010011000010100000111111101011001;
            sine_reg0   <= 36'sb101101111000101110111101010000100101;
        end
        14816: begin
            cosine_reg0 <= 36'sb11010011000110000100100011011000000;
            sine_reg0   <= 36'sb101101111001011000011001100110110100;
        end
        14817: begin
            cosine_reg0 <= 36'sb11010011001001100111111110111100000;
            sine_reg0   <= 36'sb101101111010000001110110101001101101;
        end
        14818: begin
            cosine_reg0 <= 36'sb11010011001101001011010010010111001;
            sine_reg0   <= 36'sb101101111010101011010100011001001111;
        end
        14819: begin
            cosine_reg0 <= 36'sb11010011010000101110011101101001000;
            sine_reg0   <= 36'sb101101111011010100110010110101011001;
        end
        14820: begin
            cosine_reg0 <= 36'sb11010011010100010001100000110001101;
            sine_reg0   <= 36'sb101101111011111110010001111110001000;
        end
        14821: begin
            cosine_reg0 <= 36'sb11010011010111110100011011110000111;
            sine_reg0   <= 36'sb101101111100100111110001110011011100;
        end
        14822: begin
            cosine_reg0 <= 36'sb11010011011011010111001110100110101;
            sine_reg0   <= 36'sb101101111101010001010010010101010011;
        end
        14823: begin
            cosine_reg0 <= 36'sb11010011011110111001111001010010101;
            sine_reg0   <= 36'sb101101111101111010110011100011101100;
        end
        14824: begin
            cosine_reg0 <= 36'sb11010011100010011100011011110100111;
            sine_reg0   <= 36'sb101101111110100100010101011110100011;
        end
        14825: begin
            cosine_reg0 <= 36'sb11010011100101111110110110001101001;
            sine_reg0   <= 36'sb101101111111001101111000000101111001;
        end
        14826: begin
            cosine_reg0 <= 36'sb11010011101001100001001000011011010;
            sine_reg0   <= 36'sb101101111111110111011011011001101011;
        end
        14827: begin
            cosine_reg0 <= 36'sb11010011101101000011010010011111010;
            sine_reg0   <= 36'sb101110000000100000111111011001111000;
        end
        14828: begin
            cosine_reg0 <= 36'sb11010011110000100101010100011000110;
            sine_reg0   <= 36'sb101110000001001010100100000110011110;
        end
        14829: begin
            cosine_reg0 <= 36'sb11010011110100000111001110000111111;
            sine_reg0   <= 36'sb101110000001110100001001011111011011;
        end
        14830: begin
            cosine_reg0 <= 36'sb11010011110111101000111111101100011;
            sine_reg0   <= 36'sb101110000010011101101111100100101111;
        end
        14831: begin
            cosine_reg0 <= 36'sb11010011111011001010101001000110001;
            sine_reg0   <= 36'sb101110000011000111010110010110010111;
        end
        14832: begin
            cosine_reg0 <= 36'sb11010011111110101100001010010100111;
            sine_reg0   <= 36'sb101110000011110000111101110100010001;
        end
        14833: begin
            cosine_reg0 <= 36'sb11010100000010001101100011011000101;
            sine_reg0   <= 36'sb101110000100011010100101111110011101;
        end
        14834: begin
            cosine_reg0 <= 36'sb11010100000101101110110100010001010;
            sine_reg0   <= 36'sb101110000101000100001110110100111001;
        end
        14835: begin
            cosine_reg0 <= 36'sb11010100001001001111111100111110100;
            sine_reg0   <= 36'sb101110000101101101111000010111100010;
        end
        14836: begin
            cosine_reg0 <= 36'sb11010100001100110000111101100000011;
            sine_reg0   <= 36'sb101110000110010111100010100110011000;
        end
        14837: begin
            cosine_reg0 <= 36'sb11010100010000010001110101110110101;
            sine_reg0   <= 36'sb101110000111000001001101100001011000;
        end
        14838: begin
            cosine_reg0 <= 36'sb11010100010011110010100110000001001;
            sine_reg0   <= 36'sb101110000111101010111001001000100001;
        end
        14839: begin
            cosine_reg0 <= 36'sb11010100010111010011001101111111111;
            sine_reg0   <= 36'sb101110001000010100100101011011110011;
        end
        14840: begin
            cosine_reg0 <= 36'sb11010100011010110011101101110010100;
            sine_reg0   <= 36'sb101110001000111110010010011011001001;
        end
        14841: begin
            cosine_reg0 <= 36'sb11010100011110010100000101011001001;
            sine_reg0   <= 36'sb101110001001101000000000000110100101;
        end
        14842: begin
            cosine_reg0 <= 36'sb11010100100001110100010100110011011;
            sine_reg0   <= 36'sb101110001010010001101110011110000011;
        end
        14843: begin
            cosine_reg0 <= 36'sb11010100100101010100011100000001011;
            sine_reg0   <= 36'sb101110001010111011011101100001100010;
        end
        14844: begin
            cosine_reg0 <= 36'sb11010100101000110100011011000010110;
            sine_reg0   <= 36'sb101110001011100101001101010001000000;
        end
        14845: begin
            cosine_reg0 <= 36'sb11010100101100010100010001110111100;
            sine_reg0   <= 36'sb101110001100001110111101101100011101;
        end
        14846: begin
            cosine_reg0 <= 36'sb11010100101111110100000000011111011;
            sine_reg0   <= 36'sb101110001100111000101110110011110101;
        end
        14847: begin
            cosine_reg0 <= 36'sb11010100110011010011100110111010011;
            sine_reg0   <= 36'sb101110001101100010100000100111001001;
        end
        14848: begin
            cosine_reg0 <= 36'sb11010100110110110011000101001000011;
            sine_reg0   <= 36'sb101110001110001100010011000110010101;
        end
        14849: begin
            cosine_reg0 <= 36'sb11010100111010010010011011001001001;
            sine_reg0   <= 36'sb101110001110110110000110010001011001;
        end
        14850: begin
            cosine_reg0 <= 36'sb11010100111101110001101000111100100;
            sine_reg0   <= 36'sb101110001111011111111010001000010010;
        end
        14851: begin
            cosine_reg0 <= 36'sb11010101000001010000101110100010011;
            sine_reg0   <= 36'sb101110010000001001101110101011000000;
        end
        14852: begin
            cosine_reg0 <= 36'sb11010101000100101111101011111010110;
            sine_reg0   <= 36'sb101110010000110011100011111001100000;
        end
        14853: begin
            cosine_reg0 <= 36'sb11010101001000001110100001000101011;
            sine_reg0   <= 36'sb101110010001011101011001110011110010;
        end
        14854: begin
            cosine_reg0 <= 36'sb11010101001011101101001110000010000;
            sine_reg0   <= 36'sb101110010010000111010000011001110011;
        end
        14855: begin
            cosine_reg0 <= 36'sb11010101001111001011110010110000110;
            sine_reg0   <= 36'sb101110010010110001000111101011100001;
        end
        14856: begin
            cosine_reg0 <= 36'sb11010101010010101010001111010001010;
            sine_reg0   <= 36'sb101110010011011010111111101000111100;
        end
        14857: begin
            cosine_reg0 <= 36'sb11010101010110001000100011100011101;
            sine_reg0   <= 36'sb101110010100000100111000010010000001;
        end
        14858: begin
            cosine_reg0 <= 36'sb11010101011001100110101111100111100;
            sine_reg0   <= 36'sb101110010100101110110001100110101111;
        end
        14859: begin
            cosine_reg0 <= 36'sb11010101011101000100110011011100110;
            sine_reg0   <= 36'sb101110010101011000101011100111000100;
        end
        14860: begin
            cosine_reg0 <= 36'sb11010101100000100010101111000011100;
            sine_reg0   <= 36'sb101110010110000010100110010010111111;
        end
        14861: begin
            cosine_reg0 <= 36'sb11010101100100000000100010011011010;
            sine_reg0   <= 36'sb101110010110101100100001101010011110;
        end
        14862: begin
            cosine_reg0 <= 36'sb11010101100111011110001101100100001;
            sine_reg0   <= 36'sb101110010111010110011101101101100000;
        end
        14863: begin
            cosine_reg0 <= 36'sb11010101101010111011110000011110000;
            sine_reg0   <= 36'sb101110011000000000011010011100000010;
        end
        14864: begin
            cosine_reg0 <= 36'sb11010101101110011001001011001000101;
            sine_reg0   <= 36'sb101110011000101010010111110110000100;
        end
        14865: begin
            cosine_reg0 <= 36'sb11010101110001110110011101100011111;
            sine_reg0   <= 36'sb101110011001010100010101111011100011;
        end
        14866: begin
            cosine_reg0 <= 36'sb11010101110101010011100111101111101;
            sine_reg0   <= 36'sb101110011001111110010100101100011110;
        end
        14867: begin
            cosine_reg0 <= 36'sb11010101111000110000101001101011111;
            sine_reg0   <= 36'sb101110011010101000010100001000110100;
        end
        14868: begin
            cosine_reg0 <= 36'sb11010101111100001101100011011000010;
            sine_reg0   <= 36'sb101110011011010010010100010000100010;
        end
        14869: begin
            cosine_reg0 <= 36'sb11010101111111101010010100110100110;
            sine_reg0   <= 36'sb101110011011111100010101000011100111;
        end
        14870: begin
            cosine_reg0 <= 36'sb11010110000011000110111110000001011;
            sine_reg0   <= 36'sb101110011100100110010110100010000010;
        end
        14871: begin
            cosine_reg0 <= 36'sb11010110000110100011011110111101110;
            sine_reg0   <= 36'sb101110011101010000011000101011110001;
        end
        14872: begin
            cosine_reg0 <= 36'sb11010110001001111111110111101001111;
            sine_reg0   <= 36'sb101110011101111010011011100000110010;
        end
        14873: begin
            cosine_reg0 <= 36'sb11010110001101011100001000000101101;
            sine_reg0   <= 36'sb101110011110100100011111000001000100;
        end
        14874: begin
            cosine_reg0 <= 36'sb11010110010000111000010000010000110;
            sine_reg0   <= 36'sb101110011111001110100011001100100100;
        end
        14875: begin
            cosine_reg0 <= 36'sb11010110010100010100010000001011010;
            sine_reg0   <= 36'sb101110011111111000101000000011010010;
        end
        14876: begin
            cosine_reg0 <= 36'sb11010110010111110000000111110100111;
            sine_reg0   <= 36'sb101110100000100010101101100101001100;
        end
        14877: begin
            cosine_reg0 <= 36'sb11010110011011001011110111001101101;
            sine_reg0   <= 36'sb101110100001001100110011110010010000;
        end
        14878: begin
            cosine_reg0 <= 36'sb11010110011110100111011110010101011;
            sine_reg0   <= 36'sb101110100001110110111010101010011101;
        end
        14879: begin
            cosine_reg0 <= 36'sb11010110100010000010111101001011111;
            sine_reg0   <= 36'sb101110100010100001000010001101110000;
        end
        14880: begin
            cosine_reg0 <= 36'sb11010110100101011110010011110001000;
            sine_reg0   <= 36'sb101110100011001011001010011100001001;
        end
        14881: begin
            cosine_reg0 <= 36'sb11010110101000111001100010000100101;
            sine_reg0   <= 36'sb101110100011110101010011010101100101;
        end
        14882: begin
            cosine_reg0 <= 36'sb11010110101100010100101000000110101;
            sine_reg0   <= 36'sb101110100100011111011100111010000100;
        end
        14883: begin
            cosine_reg0 <= 36'sb11010110101111101111100101110111000;
            sine_reg0   <= 36'sb101110100101001001100111001001100010;
        end
        14884: begin
            cosine_reg0 <= 36'sb11010110110011001010011011010101100;
            sine_reg0   <= 36'sb101110100101110011110010000100000000;
        end
        14885: begin
            cosine_reg0 <= 36'sb11010110110110100101001000100010000;
            sine_reg0   <= 36'sb101110100110011101111101101001011011;
        end
        14886: begin
            cosine_reg0 <= 36'sb11010110111001111111101101011100010;
            sine_reg0   <= 36'sb101110100111001000001001111001110001;
        end
        14887: begin
            cosine_reg0 <= 36'sb11010110111101011010001010000100011;
            sine_reg0   <= 36'sb101110100111110010010110110101000001;
        end
        14888: begin
            cosine_reg0 <= 36'sb11010111000000110100011110011010001;
            sine_reg0   <= 36'sb101110101000011100100100011011001010;
        end
        14889: begin
            cosine_reg0 <= 36'sb11010111000100001110101010011101010;
            sine_reg0   <= 36'sb101110101001000110110010101100001001;
        end
        14890: begin
            cosine_reg0 <= 36'sb11010111000111101000101110001101110;
            sine_reg0   <= 36'sb101110101001110001000001100111111101;
        end
        14891: begin
            cosine_reg0 <= 36'sb11010111001011000010101001101011100;
            sine_reg0   <= 36'sb101110101010011011010001001110100100;
        end
        14892: begin
            cosine_reg0 <= 36'sb11010111001110011100011100110110010;
            sine_reg0   <= 36'sb101110101011000101100001011111111110;
        end
        14893: begin
            cosine_reg0 <= 36'sb11010111010001110110000111101110001;
            sine_reg0   <= 36'sb101110101011101111110010011100000111;
        end
        14894: begin
            cosine_reg0 <= 36'sb11010111010101001111101010010010101;
            sine_reg0   <= 36'sb101110101100011010000100000010111111;
        end
        14895: begin
            cosine_reg0 <= 36'sb11010111011000101001000100100100000;
            sine_reg0   <= 36'sb101110101101000100010110010100100100;
        end
        14896: begin
            cosine_reg0 <= 36'sb11010111011100000010010110100001110;
            sine_reg0   <= 36'sb101110101101101110101001010000110100;
        end
        14897: begin
            cosine_reg0 <= 36'sb11010111011111011011100000001100000;
            sine_reg0   <= 36'sb101110101110011000111100110111101101;
        end
        14898: begin
            cosine_reg0 <= 36'sb11010111100010110100100001100010101;
            sine_reg0   <= 36'sb101110101111000011010001001001001111;
        end
        14899: begin
            cosine_reg0 <= 36'sb11010111100110001101011010100101011;
            sine_reg0   <= 36'sb101110101111101101100110000101010111;
        end
        14900: begin
            cosine_reg0 <= 36'sb11010111101001100110001011010100001;
            sine_reg0   <= 36'sb101110110000010111111011101100000100;
        end
        14901: begin
            cosine_reg0 <= 36'sb11010111101100111110110011101110110;
            sine_reg0   <= 36'sb101110110001000010010001111101010011;
        end
        14902: begin
            cosine_reg0 <= 36'sb11010111110000010111010011110101010;
            sine_reg0   <= 36'sb101110110001101100101000111001000101;
        end
        14903: begin
            cosine_reg0 <= 36'sb11010111110011101111101011100111010;
            sine_reg0   <= 36'sb101110110010010111000000011111010110;
        end
        14904: begin
            cosine_reg0 <= 36'sb11010111110111000111111011000100111;
            sine_reg0   <= 36'sb101110110011000001011000110000000101;
        end
        14905: begin
            cosine_reg0 <= 36'sb11010111111010100000000010001101111;
            sine_reg0   <= 36'sb101110110011101011110001101011010001;
        end
        14906: begin
            cosine_reg0 <= 36'sb11010111111101111000000001000010001;
            sine_reg0   <= 36'sb101110110100010110001011010000111000;
        end
        14907: begin
            cosine_reg0 <= 36'sb11011000000001001111110111100001100;
            sine_reg0   <= 36'sb101110110101000000100101100000111000;
        end
        14908: begin
            cosine_reg0 <= 36'sb11011000000100100111100101101011110;
            sine_reg0   <= 36'sb101110110101101011000000011011001111;
        end
        14909: begin
            cosine_reg0 <= 36'sb11011000000111111111001011100001000;
            sine_reg0   <= 36'sb101110110110010101011011111111111101;
        end
        14910: begin
            cosine_reg0 <= 36'sb11011000001011010110101001000001000;
            sine_reg0   <= 36'sb101110110110111111111000001110111111;
        end
        14911: begin
            cosine_reg0 <= 36'sb11011000001110101101111110001011100;
            sine_reg0   <= 36'sb101110110111101010010101001000010100;
        end
        14912: begin
            cosine_reg0 <= 36'sb11011000010010000101001011000000100;
            sine_reg0   <= 36'sb101110111000010100110010101011111010;
        end
        14913: begin
            cosine_reg0 <= 36'sb11011000010101011100001111011111111;
            sine_reg0   <= 36'sb101110111000111111010000111001101111;
        end
        14914: begin
            cosine_reg0 <= 36'sb11011000011000110011001011101001100;
            sine_reg0   <= 36'sb101110111001101001101111110001110010;
        end
        14915: begin
            cosine_reg0 <= 36'sb11011000011100001001111111011101001;
            sine_reg0   <= 36'sb101110111010010100001111010100000010;
        end
        14916: begin
            cosine_reg0 <= 36'sb11011000011111100000101010111010110;
            sine_reg0   <= 36'sb101110111010111110101111100000011100;
        end
        14917: begin
            cosine_reg0 <= 36'sb11011000100010110111001110000010010;
            sine_reg0   <= 36'sb101110111011101001010000010110111111;
        end
        14918: begin
            cosine_reg0 <= 36'sb11011000100110001101101000110011011;
            sine_reg0   <= 36'sb101110111100010011110001110111101001;
        end
        14919: begin
            cosine_reg0 <= 36'sb11011000101001100011111011001110001;
            sine_reg0   <= 36'sb101110111100111110010100000010011001;
        end
        14920: begin
            cosine_reg0 <= 36'sb11011000101100111010000101010010010;
            sine_reg0   <= 36'sb101110111101101000110110110111001100;
        end
        14921: begin
            cosine_reg0 <= 36'sb11011000110000010000000110111111110;
            sine_reg0   <= 36'sb101110111110010011011010010110000011;
        end
        14922: begin
            cosine_reg0 <= 36'sb11011000110011100110000000010110011;
            sine_reg0   <= 36'sb101110111110111101111110011110111001;
        end
        14923: begin
            cosine_reg0 <= 36'sb11011000110110111011110001010110001;
            sine_reg0   <= 36'sb101110111111101000100011010001101111;
        end
        14924: begin
            cosine_reg0 <= 36'sb11011000111010010001011001111110110;
            sine_reg0   <= 36'sb101111000000010011001000101110100011;
        end
        14925: begin
            cosine_reg0 <= 36'sb11011000111101100110111010010000001;
            sine_reg0   <= 36'sb101111000000111101101110110101010010;
        end
        14926: begin
            cosine_reg0 <= 36'sb11011001000000111100010010001010010;
            sine_reg0   <= 36'sb101111000001101000010101100101111011;
        end
        14927: begin
            cosine_reg0 <= 36'sb11011001000100010001100001101100111;
            sine_reg0   <= 36'sb101111000010010010111101000000011101;
        end
        14928: begin
            cosine_reg0 <= 36'sb11011001000111100110101000110111111;
            sine_reg0   <= 36'sb101111000010111101100101000100110110;
        end
        14929: begin
            cosine_reg0 <= 36'sb11011001001010111011100111101011010;
            sine_reg0   <= 36'sb101111000011101000001101110011000100;
        end
        14930: begin
            cosine_reg0 <= 36'sb11011001001110010000011110000110101;
            sine_reg0   <= 36'sb101111000100010010110111001011000101;
        end
        14931: begin
            cosine_reg0 <= 36'sb11011001010001100101001100001010001;
            sine_reg0   <= 36'sb101111000100111101100001001100111001;
        end
        14932: begin
            cosine_reg0 <= 36'sb11011001010100111001110001110101100;
            sine_reg0   <= 36'sb101111000101101000001011111000011101;
        end
        14933: begin
            cosine_reg0 <= 36'sb11011001011000001110001111001000110;
            sine_reg0   <= 36'sb101111000110010010110111001101101111;
        end
        14934: begin
            cosine_reg0 <= 36'sb11011001011011100010100100000011100;
            sine_reg0   <= 36'sb101111000110111101100011001100101110;
        end
        14935: begin
            cosine_reg0 <= 36'sb11011001011110110110110000100101110;
            sine_reg0   <= 36'sb101111000111101000001111110101011001;
        end
        14936: begin
            cosine_reg0 <= 36'sb11011001100010001010110100101111100;
            sine_reg0   <= 36'sb101111001000010010111101000111101110;
        end
        14937: begin
            cosine_reg0 <= 36'sb11011001100101011110110000100000100;
            sine_reg0   <= 36'sb101111001000111101101011000011101010;
        end
        14938: begin
            cosine_reg0 <= 36'sb11011001101000110010100011111000100;
            sine_reg0   <= 36'sb101111001001101000011001101001001101;
        end
        14939: begin
            cosine_reg0 <= 36'sb11011001101100000110001110110111101;
            sine_reg0   <= 36'sb101111001010010011001000111000010101;
        end
        14940: begin
            cosine_reg0 <= 36'sb11011001101111011001110001011101100;
            sine_reg0   <= 36'sb101111001010111101111000110001000000;
        end
        14941: begin
            cosine_reg0 <= 36'sb11011001110010101101001011101010010;
            sine_reg0   <= 36'sb101111001011101000101001010011001100;
        end
        14942: begin
            cosine_reg0 <= 36'sb11011001110110000000011101011101101;
            sine_reg0   <= 36'sb101111001100010011011010011110111000;
        end
        14943: begin
            cosine_reg0 <= 36'sb11011001111001010011100110110111011;
            sine_reg0   <= 36'sb101111001100111110001100010100000010;
        end
        14944: begin
            cosine_reg0 <= 36'sb11011001111100100110100111110111100;
            sine_reg0   <= 36'sb101111001101101000111110110010101001;
        end
        14945: begin
            cosine_reg0 <= 36'sb11011001111111111001100000011110000;
            sine_reg0   <= 36'sb101111001110010011110001111010101011;
        end
        14946: begin
            cosine_reg0 <= 36'sb11011010000011001100010000101010100;
            sine_reg0   <= 36'sb101111001110111110100101101100000110;
        end
        14947: begin
            cosine_reg0 <= 36'sb11011010000110011110111000011101000;
            sine_reg0   <= 36'sb101111001111101001011010000110111000;
        end
        14948: begin
            cosine_reg0 <= 36'sb11011010001001110001010111110101011;
            sine_reg0   <= 36'sb101111010000010100001111001011000001;
        end
        14949: begin
            cosine_reg0 <= 36'sb11011010001101000011101110110011100;
            sine_reg0   <= 36'sb101111010000111111000100111000011101;
        end
        14950: begin
            cosine_reg0 <= 36'sb11011010010000010101111101010111001;
            sine_reg0   <= 36'sb101111010001101001111011001111001101;
        end
        14951: begin
            cosine_reg0 <= 36'sb11011010010011101000000011100000011;
            sine_reg0   <= 36'sb101111010010010100110010001111001101;
        end
        14952: begin
            cosine_reg0 <= 36'sb11011010010110111010000001001110111;
            sine_reg0   <= 36'sb101111010010111111101001111000011101;
        end
        14953: begin
            cosine_reg0 <= 36'sb11011010011010001011110110100010101;
            sine_reg0   <= 36'sb101111010011101010100010001010111010;
        end
        14954: begin
            cosine_reg0 <= 36'sb11011010011101011101100011011011011;
            sine_reg0   <= 36'sb101111010100010101011011000110100011;
        end
        14955: begin
            cosine_reg0 <= 36'sb11011010100000101111000111111001010;
            sine_reg0   <= 36'sb101111010101000000010100101011010111;
        end
        14956: begin
            cosine_reg0 <= 36'sb11011010100100000000100011111011111;
            sine_reg0   <= 36'sb101111010101101011001110111001010011;
        end
        14957: begin
            cosine_reg0 <= 36'sb11011010100111010001110111100011010;
            sine_reg0   <= 36'sb101111010110010110001001110000010111;
        end
        14958: begin
            cosine_reg0 <= 36'sb11011010101010100011000010101111010;
            sine_reg0   <= 36'sb101111010111000001000101010000011111;
        end
        14959: begin
            cosine_reg0 <= 36'sb11011010101101110100000101011111101;
            sine_reg0   <= 36'sb101111010111101100000001011001101100;
        end
        14960: begin
            cosine_reg0 <= 36'sb11011010110001000100111111110100100;
            sine_reg0   <= 36'sb101111011000010110111110001011111011;
        end
        14961: begin
            cosine_reg0 <= 36'sb11011010110100010101110001101101100;
            sine_reg0   <= 36'sb101111011001000001111011100111001010;
        end
        14962: begin
            cosine_reg0 <= 36'sb11011010110111100110011011001010100;
            sine_reg0   <= 36'sb101111011001101100111001101011010111;
        end
        14963: begin
            cosine_reg0 <= 36'sb11011010111010110110111100001011101;
            sine_reg0   <= 36'sb101111011010010111111000011000100010;
        end
        14964: begin
            cosine_reg0 <= 36'sb11011010111110000111010100110000100;
            sine_reg0   <= 36'sb101111011011000010110111101110101001;
        end
        14965: begin
            cosine_reg0 <= 36'sb11011011000001010111100100111001000;
            sine_reg0   <= 36'sb101111011011101101110111101101101001;
        end
        14966: begin
            cosine_reg0 <= 36'sb11011011000100100111101100100101010;
            sine_reg0   <= 36'sb101111011100011000111000010101100001;
        end
        14967: begin
            cosine_reg0 <= 36'sb11011011000111110111101011110100111;
            sine_reg0   <= 36'sb101111011101000011111001100110010000;
        end
        14968: begin
            cosine_reg0 <= 36'sb11011011001011000111100010100111111;
            sine_reg0   <= 36'sb101111011101101110111011011111110100;
        end
        14969: begin
            cosine_reg0 <= 36'sb11011011001110010111010000111110000;
            sine_reg0   <= 36'sb101111011110011001111110000010001011;
        end
        14970: begin
            cosine_reg0 <= 36'sb11011011010001100110110110110111010;
            sine_reg0   <= 36'sb101111011111000101000001001101010011;
        end
        14971: begin
            cosine_reg0 <= 36'sb11011011010100110110010100010011100;
            sine_reg0   <= 36'sb101111011111110000000101000001001011;
        end
        14972: begin
            cosine_reg0 <= 36'sb11011011011000000101101001010010101;
            sine_reg0   <= 36'sb101111100000011011001001011101110010;
        end
        14973: begin
            cosine_reg0 <= 36'sb11011011011011010100110101110100011;
            sine_reg0   <= 36'sb101111100001000110001110100011000100;
        end
        14974: begin
            cosine_reg0 <= 36'sb11011011011110100011111001111000110;
            sine_reg0   <= 36'sb101111100001110001010100010001000010;
        end
        14975: begin
            cosine_reg0 <= 36'sb11011011100001110010110101011111100;
            sine_reg0   <= 36'sb101111100010011100011010100111101001;
        end
        14976: begin
            cosine_reg0 <= 36'sb11011011100101000001101000101000101;
            sine_reg0   <= 36'sb101111100011000111100001100110111000;
        end
        14977: begin
            cosine_reg0 <= 36'sb11011011101000010000010011010100000;
            sine_reg0   <= 36'sb101111100011110010101001001110101100;
        end
        14978: begin
            cosine_reg0 <= 36'sb11011011101011011110110101100001100;
            sine_reg0   <= 36'sb101111100100011101110001011111000101;
        end
        14979: begin
            cosine_reg0 <= 36'sb11011011101110101101001111010000111;
            sine_reg0   <= 36'sb101111100101001000111010011000000000;
        end
        14980: begin
            cosine_reg0 <= 36'sb11011011110001111011100000100010010;
            sine_reg0   <= 36'sb101111100101110100000011111001011100;
        end
        14981: begin
            cosine_reg0 <= 36'sb11011011110101001001101001010101001;
            sine_reg0   <= 36'sb101111100110011111001110000011010111;
        end
        14982: begin
            cosine_reg0 <= 36'sb11011011111000010111101001101001110;
            sine_reg0   <= 36'sb101111100111001010011000110101110000;
        end
        14983: begin
            cosine_reg0 <= 36'sb11011011111011100101100001011111110;
            sine_reg0   <= 36'sb101111100111110101100100010000100101;
        end
        14984: begin
            cosine_reg0 <= 36'sb11011011111110110011010000110111001;
            sine_reg0   <= 36'sb101111101000100000110000010011110100;
        end
        14985: begin
            cosine_reg0 <= 36'sb11011100000010000000110111101111110;
            sine_reg0   <= 36'sb101111101001001011111100111111011100;
        end
        14986: begin
            cosine_reg0 <= 36'sb11011100000101001110010110001001011;
            sine_reg0   <= 36'sb101111101001110111001010010011011010;
        end
        14987: begin
            cosine_reg0 <= 36'sb11011100001000011011101100000100000;
            sine_reg0   <= 36'sb101111101010100010011000001111101110;
        end
        14988: begin
            cosine_reg0 <= 36'sb11011100001011101000111001011111100;
            sine_reg0   <= 36'sb101111101011001101100110110100010101;
        end
        14989: begin
            cosine_reg0 <= 36'sb11011100001110110101111110011011110;
            sine_reg0   <= 36'sb101111101011111000110110000001001110;
        end
        14990: begin
            cosine_reg0 <= 36'sb11011100010010000010111010111000101;
            sine_reg0   <= 36'sb101111101100100100000101110110011000;
        end
        14991: begin
            cosine_reg0 <= 36'sb11011100010101001111101110110101111;
            sine_reg0   <= 36'sb101111101101001111010110010011110000;
        end
        14992: begin
            cosine_reg0 <= 36'sb11011100011000011100011010010011100;
            sine_reg0   <= 36'sb101111101101111010100111011001010101;
        end
        14993: begin
            cosine_reg0 <= 36'sb11011100011011101000111101010001011;
            sine_reg0   <= 36'sb101111101110100101111001000111000101;
        end
        14994: begin
            cosine_reg0 <= 36'sb11011100011110110101010111101111011;
            sine_reg0   <= 36'sb101111101111010001001011011100111111;
        end
        14995: begin
            cosine_reg0 <= 36'sb11011100100010000001101001101101011;
            sine_reg0   <= 36'sb101111101111111100011110011011000001;
        end
        14996: begin
            cosine_reg0 <= 36'sb11011100100101001101110011001011010;
            sine_reg0   <= 36'sb101111110000100111110010000001001001;
        end
        14997: begin
            cosine_reg0 <= 36'sb11011100101000011001110100001000110;
            sine_reg0   <= 36'sb101111110001010011000110001111010101;
        end
        14998: begin
            cosine_reg0 <= 36'sb11011100101011100101101100100110000;
            sine_reg0   <= 36'sb101111110001111110011011000101100100;
        end
        14999: begin
            cosine_reg0 <= 36'sb11011100101110110001011100100010101;
            sine_reg0   <= 36'sb101111110010101001110000100011110101;
        end
        15000: begin
            cosine_reg0 <= 36'sb11011100110001111101000011111110101;
            sine_reg0   <= 36'sb101111110011010101000110101010000101;
        end
        15001: begin
            cosine_reg0 <= 36'sb11011100110101001000100010111010000;
            sine_reg0   <= 36'sb101111110100000000011101011000010011;
        end
        15002: begin
            cosine_reg0 <= 36'sb11011100111000010011111001010100011;
            sine_reg0   <= 36'sb101111110100101011110100101110011101;
        end
        15003: begin
            cosine_reg0 <= 36'sb11011100111011011111000111001101110;
            sine_reg0   <= 36'sb101111110101010111001100101100100010;
        end
        15004: begin
            cosine_reg0 <= 36'sb11011100111110101010001100100110001;
            sine_reg0   <= 36'sb101111110110000010100101010010100000;
        end
        15005: begin
            cosine_reg0 <= 36'sb11011101000001110101001001011101001;
            sine_reg0   <= 36'sb101111110110101101111110100000010101;
        end
        15006: begin
            cosine_reg0 <= 36'sb11011101000100111111111101110010110;
            sine_reg0   <= 36'sb101111110111011001011000010101111111;
        end
        15007: begin
            cosine_reg0 <= 36'sb11011101001000001010101001100111000;
            sine_reg0   <= 36'sb101111111000000100110010110011011101;
        end
        15008: begin
            cosine_reg0 <= 36'sb11011101001011010101001100111001101;
            sine_reg0   <= 36'sb101111111000110000001101111000101101;
        end
        15009: begin
            cosine_reg0 <= 36'sb11011101001110011111100111101010011;
            sine_reg0   <= 36'sb101111111001011011101001100101101110;
        end
        15010: begin
            cosine_reg0 <= 36'sb11011101010001101001111001111001011;
            sine_reg0   <= 36'sb101111111010000111000101111010011110;
        end
        15011: begin
            cosine_reg0 <= 36'sb11011101010100110100000011100110011;
            sine_reg0   <= 36'sb101111111010110010100010110110111011;
        end
        15012: begin
            cosine_reg0 <= 36'sb11011101010111111110000100110001011;
            sine_reg0   <= 36'sb101111111011011110000000011011000011;
        end
        15013: begin
            cosine_reg0 <= 36'sb11011101011011000111111101011010000;
            sine_reg0   <= 36'sb101111111100001001011110100110110101;
        end
        15014: begin
            cosine_reg0 <= 36'sb11011101011110010001101101100000011;
            sine_reg0   <= 36'sb101111111100110100111101011010001111;
        end
        15015: begin
            cosine_reg0 <= 36'sb11011101100001011011010101000100010;
            sine_reg0   <= 36'sb101111111101100000011100110101010000;
        end
        15016: begin
            cosine_reg0 <= 36'sb11011101100100100100110100000101101;
            sine_reg0   <= 36'sb101111111110001011111100110111110110;
        end
        15017: begin
            cosine_reg0 <= 36'sb11011101100111101110001010100100010;
            sine_reg0   <= 36'sb101111111110110111011101100001111110;
        end
        15018: begin
            cosine_reg0 <= 36'sb11011101101010110111011000100000000;
            sine_reg0   <= 36'sb101111111111100010111110110011101000;
        end
        15019: begin
            cosine_reg0 <= 36'sb11011101101110000000011101111000111;
            sine_reg0   <= 36'sb110000000000001110100000101100110010;
        end
        15020: begin
            cosine_reg0 <= 36'sb11011101110001001001011010101110101;
            sine_reg0   <= 36'sb110000000000111010000011001101011010;
        end
        15021: begin
            cosine_reg0 <= 36'sb11011101110100010010001111000001001;
            sine_reg0   <= 36'sb110000000001100101100110010101011110;
        end
        15022: begin
            cosine_reg0 <= 36'sb11011101110111011010111010110000011;
            sine_reg0   <= 36'sb110000000010010001001010000100111101;
        end
        15023: begin
            cosine_reg0 <= 36'sb11011101111010100011011101111100010;
            sine_reg0   <= 36'sb110000000010111100101110011011110100;
        end
        15024: begin
            cosine_reg0 <= 36'sb11011101111101101011111000100100100;
            sine_reg0   <= 36'sb110000000011101000010011011010000100;
        end
        15025: begin
            cosine_reg0 <= 36'sb11011110000000110100001010101001001;
            sine_reg0   <= 36'sb110000000100010011111000111111101000;
        end
        15026: begin
            cosine_reg0 <= 36'sb11011110000011111100010100001001111;
            sine_reg0   <= 36'sb110000000100111111011111001100100001;
        end
        15027: begin
            cosine_reg0 <= 36'sb11011110000111000100010101000110110;
            sine_reg0   <= 36'sb110000000101101011000110000000101100;
        end
        15028: begin
            cosine_reg0 <= 36'sb11011110001010001100001101011111101;
            sine_reg0   <= 36'sb110000000110010110101101011100001000;
        end
        15029: begin
            cosine_reg0 <= 36'sb11011110001101010011111101010100011;
            sine_reg0   <= 36'sb110000000111000010010101011110110011;
        end
        15030: begin
            cosine_reg0 <= 36'sb11011110010000011011100100100100110;
            sine_reg0   <= 36'sb110000000111101101111110001000101011;
        end
        15031: begin
            cosine_reg0 <= 36'sb11011110010011100011000011010000110;
            sine_reg0   <= 36'sb110000001000011001100111011001101110;
        end
        15032: begin
            cosine_reg0 <= 36'sb11011110010110101010011001011000010;
            sine_reg0   <= 36'sb110000001001000101010001010001111100;
        end
        15033: begin
            cosine_reg0 <= 36'sb11011110011001110001100110111011001;
            sine_reg0   <= 36'sb110000001001110000111011110001010010;
        end
        15034: begin
            cosine_reg0 <= 36'sb11011110011100111000101011111001010;
            sine_reg0   <= 36'sb110000001010011100100110110111101110;
        end
        15035: begin
            cosine_reg0 <= 36'sb11011110011111111111101000010010100;
            sine_reg0   <= 36'sb110000001011001000010010100101001111;
        end
        15036: begin
            cosine_reg0 <= 36'sb11011110100011000110011100000110110;
            sine_reg0   <= 36'sb110000001011110011111110111001110011;
        end
        15037: begin
            cosine_reg0 <= 36'sb11011110100110001101000111010101111;
            sine_reg0   <= 36'sb110000001100011111101011110101011001;
        end
        15038: begin
            cosine_reg0 <= 36'sb11011110101001010011101001111111110;
            sine_reg0   <= 36'sb110000001101001011011001010111111110;
        end
        15039: begin
            cosine_reg0 <= 36'sb11011110101100011010000100000100011;
            sine_reg0   <= 36'sb110000001101110111000111100001100001;
        end
        15040: begin
            cosine_reg0 <= 36'sb11011110101111100000010101100011011;
            sine_reg0   <= 36'sb110000001110100010110110010010000001;
        end
        15041: begin
            cosine_reg0 <= 36'sb11011110110010100110011110011100111;
            sine_reg0   <= 36'sb110000001111001110100101101001011100;
        end
        15042: begin
            cosine_reg0 <= 36'sb11011110110101101100011110110000101;
            sine_reg0   <= 36'sb110000001111111010010101100111110000;
        end
        15043: begin
            cosine_reg0 <= 36'sb11011110111000110010010110011110100;
            sine_reg0   <= 36'sb110000010000100110000110001100111011;
        end
        15044: begin
            cosine_reg0 <= 36'sb11011110111011111000000101100110100;
            sine_reg0   <= 36'sb110000010001010001110111011000111100;
        end
        15045: begin
            cosine_reg0 <= 36'sb11011110111110111101101100001000011;
            sine_reg0   <= 36'sb110000010001111101101001001011110000;
        end
        15046: begin
            cosine_reg0 <= 36'sb11011111000010000011001010000100001;
            sine_reg0   <= 36'sb110000010010101001011011100101010111;
        end
        15047: begin
            cosine_reg0 <= 36'sb11011111000101001000011111011001100;
            sine_reg0   <= 36'sb110000010011010101001110100101101111;
        end
        15048: begin
            cosine_reg0 <= 36'sb11011111001000001101101100001000011;
            sine_reg0   <= 36'sb110000010100000001000010001100110110;
        end
        15049: begin
            cosine_reg0 <= 36'sb11011111001011010010110000010000111;
            sine_reg0   <= 36'sb110000010100101100110110011010101001;
        end
        15050: begin
            cosine_reg0 <= 36'sb11011111001110010111101011110010101;
            sine_reg0   <= 36'sb110000010101011000101011001111001001;
        end
        15051: begin
            cosine_reg0 <= 36'sb11011111010001011100011110101101101;
            sine_reg0   <= 36'sb110000010110000100100000101010010010;
        end
        15052: begin
            cosine_reg0 <= 36'sb11011111010100100001001001000001101;
            sine_reg0   <= 36'sb110000010110110000010110101100000011;
        end
        15053: begin
            cosine_reg0 <= 36'sb11011111010111100101101010101110101;
            sine_reg0   <= 36'sb110000010111011100001101010100011011;
        end
        15054: begin
            cosine_reg0 <= 36'sb11011111011010101010000011110100101;
            sine_reg0   <= 36'sb110000011000001000000100100011011000;
        end
        15055: begin
            cosine_reg0 <= 36'sb11011111011101101110010100010011010;
            sine_reg0   <= 36'sb110000011000110011111100011000110111;
        end
        15056: begin
            cosine_reg0 <= 36'sb11011111100000110010011100001010100;
            sine_reg0   <= 36'sb110000011001011111110100110100111001;
        end
        15057: begin
            cosine_reg0 <= 36'sb11011111100011110110011011011010010;
            sine_reg0   <= 36'sb110000011010001011101101110111011001;
        end
        15058: begin
            cosine_reg0 <= 36'sb11011111100110111010010010000010011;
            sine_reg0   <= 36'sb110000011010110111100111100000011000;
        end
        15059: begin
            cosine_reg0 <= 36'sb11011111101001111110000000000010111;
            sine_reg0   <= 36'sb110000011011100011100001101111110011;
        end
        15060: begin
            cosine_reg0 <= 36'sb11011111101101000001100101011011100;
            sine_reg0   <= 36'sb110000011100001111011100100101101001;
        end
        15061: begin
            cosine_reg0 <= 36'sb11011111110000000101000010001100001;
            sine_reg0   <= 36'sb110000011100111011011000000001111000;
        end
        15062: begin
            cosine_reg0 <= 36'sb11011111110011001000010110010100101;
            sine_reg0   <= 36'sb110000011101100111010100000100011110;
        end
        15063: begin
            cosine_reg0 <= 36'sb11011111110110001011100001110100111;
            sine_reg0   <= 36'sb110000011110010011010000101101011001;
        end
        15064: begin
            cosine_reg0 <= 36'sb11011111111001001110100100101101000;
            sine_reg0   <= 36'sb110000011110111111001101111100101000;
        end
        15065: begin
            cosine_reg0 <= 36'sb11011111111100010001011110111100100;
            sine_reg0   <= 36'sb110000011111101011001011110010001010;
        end
        15066: begin
            cosine_reg0 <= 36'sb11011111111111010100010000100011100;
            sine_reg0   <= 36'sb110000100000010111001010001101111100;
        end
        15067: begin
            cosine_reg0 <= 36'sb11100000000010010110111001100001111;
            sine_reg0   <= 36'sb110000100001000011001001001111111101;
        end
        15068: begin
            cosine_reg0 <= 36'sb11100000000101011001011001110111100;
            sine_reg0   <= 36'sb110000100001101111001000111000001011;
        end
        15069: begin
            cosine_reg0 <= 36'sb11100000001000011011110001100100001;
            sine_reg0   <= 36'sb110000100010011011001001000110100100;
        end
        15070: begin
            cosine_reg0 <= 36'sb11100000001011011110000000100111110;
            sine_reg0   <= 36'sb110000100011000111001001111011000111;
        end
        15071: begin
            cosine_reg0 <= 36'sb11100000001110100000000111000010010;
            sine_reg0   <= 36'sb110000100011110011001011010101110001;
        end
        15072: begin
            cosine_reg0 <= 36'sb11100000010001100010000100110011100;
            sine_reg0   <= 36'sb110000100100011111001101010110100011;
        end
        15073: begin
            cosine_reg0 <= 36'sb11100000010100100011111001111011011;
            sine_reg0   <= 36'sb110000100101001011001111111101011000;
        end
        15074: begin
            cosine_reg0 <= 36'sb11100000010111100101100110011001110;
            sine_reg0   <= 36'sb110000100101110111010011001010010001;
        end
        15075: begin
            cosine_reg0 <= 36'sb11100000011010100111001010001110100;
            sine_reg0   <= 36'sb110000100110100011010110111101001011;
        end
        15076: begin
            cosine_reg0 <= 36'sb11100000011101101000100101011001100;
            sine_reg0   <= 36'sb110000100111001111011011010110000100;
        end
        15077: begin
            cosine_reg0 <= 36'sb11100000100000101001110111111010110;
            sine_reg0   <= 36'sb110000100111111011100000010100111011;
        end
        15078: begin
            cosine_reg0 <= 36'sb11100000100011101011000001110010000;
            sine_reg0   <= 36'sb110000101000100111100101111001101110;
        end
        15079: begin
            cosine_reg0 <= 36'sb11100000100110101100000010111111001;
            sine_reg0   <= 36'sb110000101001010011101100000100011100;
        end
        15080: begin
            cosine_reg0 <= 36'sb11100000101001101100111011100010001;
            sine_reg0   <= 36'sb110000101001111111110010110101000010;
        end
        15081: begin
            cosine_reg0 <= 36'sb11100000101100101101101011011010110;
            sine_reg0   <= 36'sb110000101010101011111010001011011111;
        end
        15082: begin
            cosine_reg0 <= 36'sb11100000101111101110010010101001000;
            sine_reg0   <= 36'sb110000101011011000000010000111110010;
        end
        15083: begin
            cosine_reg0 <= 36'sb11100000110010101110110001001100110;
            sine_reg0   <= 36'sb110000101100000100001010101001111000;
        end
        15084: begin
            cosine_reg0 <= 36'sb11100000110101101111000111000101110;
            sine_reg0   <= 36'sb110000101100110000010011110001110000;
        end
        15085: begin
            cosine_reg0 <= 36'sb11100000111000101111010100010100001;
            sine_reg0   <= 36'sb110000101101011100011101011111011001;
        end
        15086: begin
            cosine_reg0 <= 36'sb11100000111011101111011000110111100;
            sine_reg0   <= 36'sb110000101110001000100111110010101111;
        end
        15087: begin
            cosine_reg0 <= 36'sb11100000111110101111010100101111111;
            sine_reg0   <= 36'sb110000101110110100110010101011110011;
        end
        15088: begin
            cosine_reg0 <= 36'sb11100001000001101111000111111101001;
            sine_reg0   <= 36'sb110000101111100000111110001010100001;
        end
        15089: begin
            cosine_reg0 <= 36'sb11100001000100101110110010011111010;
            sine_reg0   <= 36'sb110000110000001101001010001110111001;
        end
        15090: begin
            cosine_reg0 <= 36'sb11100001000111101110010100010110000;
            sine_reg0   <= 36'sb110000110000111001010110111000111001;
        end
        15091: begin
            cosine_reg0 <= 36'sb11100001001010101101101101100001010;
            sine_reg0   <= 36'sb110000110001100101100100001000011111;
        end
        15092: begin
            cosine_reg0 <= 36'sb11100001001101101100111110000000111;
            sine_reg0   <= 36'sb110000110010010001110001111101101001;
        end
        15093: begin
            cosine_reg0 <= 36'sb11100001010000101100000101110100111;
            sine_reg0   <= 36'sb110000110010111110000000011000010101;
        end
        15094: begin
            cosine_reg0 <= 36'sb11100001010011101011000100111101000;
            sine_reg0   <= 36'sb110000110011101010001111011000100010;
        end
        15095: begin
            cosine_reg0 <= 36'sb11100001010110101001111011011001010;
            sine_reg0   <= 36'sb110000110100010110011110111110001111;
        end
        15096: begin
            cosine_reg0 <= 36'sb11100001011001101000101001001001100;
            sine_reg0   <= 36'sb110000110101000010101111001001011001;
        end
        15097: begin
            cosine_reg0 <= 36'sb11100001011100100111001110001101100;
            sine_reg0   <= 36'sb110000110101101110111111111001111111;
        end
        15098: begin
            cosine_reg0 <= 36'sb11100001011111100101101010100101010;
            sine_reg0   <= 36'sb110000110110011011010001001111111110;
        end
        15099: begin
            cosine_reg0 <= 36'sb11100001100010100011111110010000101;
            sine_reg0   <= 36'sb110000110111000111100011001011010110;
        end
        15100: begin
            cosine_reg0 <= 36'sb11100001100101100010001001001111101;
            sine_reg0   <= 36'sb110000110111110011110101101100000101;
        end
        15101: begin
            cosine_reg0 <= 36'sb11100001101000100000001011100001111;
            sine_reg0   <= 36'sb110000111000100000001000110010001001;
        end
        15102: begin
            cosine_reg0 <= 36'sb11100001101011011110000101000111011;
            sine_reg0   <= 36'sb110000111001001100011100011101011111;
        end
        15103: begin
            cosine_reg0 <= 36'sb11100001101110011011110110000000001;
            sine_reg0   <= 36'sb110000111001111000110000101110001000;
        end
        15104: begin
            cosine_reg0 <= 36'sb11100001110001011001011110001011111;
            sine_reg0   <= 36'sb110000111010100101000101100100000000;
        end
        15105: begin
            cosine_reg0 <= 36'sb11100001110100010110111101101010101;
            sine_reg0   <= 36'sb110000111011010001011010111111000110;
        end
        15106: begin
            cosine_reg0 <= 36'sb11100001110111010100010100011100001;
            sine_reg0   <= 36'sb110000111011111101110000111111011000;
        end
        15107: begin
            cosine_reg0 <= 36'sb11100001111010010001100010100000011;
            sine_reg0   <= 36'sb110000111100101010000111100100110101;
        end
        15108: begin
            cosine_reg0 <= 36'sb11100001111101001110100111110111001;
            sine_reg0   <= 36'sb110000111101010110011110101111011100;
        end
        15109: begin
            cosine_reg0 <= 36'sb11100010000000001011100100100000011;
            sine_reg0   <= 36'sb110000111110000010110110011111001001;
        end
        15110: begin
            cosine_reg0 <= 36'sb11100010000011001000011000011100000;
            sine_reg0   <= 36'sb110000111110101111001110110011111100;
        end
        15111: begin
            cosine_reg0 <= 36'sb11100010000110000101000011101001111;
            sine_reg0   <= 36'sb110000111111011011100111101101110010;
        end
        15112: begin
            cosine_reg0 <= 36'sb11100010001001000001100110001010000;
            sine_reg0   <= 36'sb110001000000001000000001001100101011;
        end
        15113: begin
            cosine_reg0 <= 36'sb11100010001011111101111111111100000;
            sine_reg0   <= 36'sb110001000000110100011011010000100101;
        end
        15114: begin
            cosine_reg0 <= 36'sb11100010001110111010010000111111111;
            sine_reg0   <= 36'sb110001000001100000110101111001011100;
        end
        15115: begin
            cosine_reg0 <= 36'sb11100010010001110110011001010101101;
            sine_reg0   <= 36'sb110001000010001101010001000111010001;
        end
        15116: begin
            cosine_reg0 <= 36'sb11100010010100110010011000111101001;
            sine_reg0   <= 36'sb110001000010111001101100111010000001;
        end
        15117: begin
            cosine_reg0 <= 36'sb11100010010111101110001111110110000;
            sine_reg0   <= 36'sb110001000011100110001001010001101011;
        end
        15118: begin
            cosine_reg0 <= 36'sb11100010011010101001111110000000100;
            sine_reg0   <= 36'sb110001000100010010100110001110001101;
        end
        15119: begin
            cosine_reg0 <= 36'sb11100010011101100101100011011100010;
            sine_reg0   <= 36'sb110001000100111111000011101111100100;
        end
        15120: begin
            cosine_reg0 <= 36'sb11100010100000100001000000001001010;
            sine_reg0   <= 36'sb110001000101101011100001110101110000;
        end
        15121: begin
            cosine_reg0 <= 36'sb11100010100011011100010100000111011;
            sine_reg0   <= 36'sb110001000110011000000000100000101111;
        end
        15122: begin
            cosine_reg0 <= 36'sb11100010100110010111011111010110100;
            sine_reg0   <= 36'sb110001000111000100011111110000011111;
        end
        15123: begin
            cosine_reg0 <= 36'sb11100010101001010010100001110110100;
            sine_reg0   <= 36'sb110001000111110000111111100100111110;
        end
        15124: begin
            cosine_reg0 <= 36'sb11100010101100001101011011100111010;
            sine_reg0   <= 36'sb110001001000011101011111111110001010;
        end
        15125: begin
            cosine_reg0 <= 36'sb11100010101111001000001100101000101;
            sine_reg0   <= 36'sb110001001001001010000000111100000010;
        end
        15126: begin
            cosine_reg0 <= 36'sb11100010110010000010110100111010101;
            sine_reg0   <= 36'sb110001001001110110100010011110100101;
        end
        15127: begin
            cosine_reg0 <= 36'sb11100010110100111101010100011101001;
            sine_reg0   <= 36'sb110001001010100011000100100101110000;
        end
        15128: begin
            cosine_reg0 <= 36'sb11100010110111110111101011001111111;
            sine_reg0   <= 36'sb110001001011001111100111010001100001;
        end
        15129: begin
            cosine_reg0 <= 36'sb11100010111010110001111001010010111;
            sine_reg0   <= 36'sb110001001011111100001010100001111000;
        end
        15130: begin
            cosine_reg0 <= 36'sb11100010111101101011111110100101111;
            sine_reg0   <= 36'sb110001001100101000101110010110110001;
        end
        15131: begin
            cosine_reg0 <= 36'sb11100011000000100101111011001001000;
            sine_reg0   <= 36'sb110001001101010101010010110000001101;
        end
        15132: begin
            cosine_reg0 <= 36'sb11100011000011011111101110111011111;
            sine_reg0   <= 36'sb110001001110000001110111101110001000;
        end
        15133: begin
            cosine_reg0 <= 36'sb11100011000110011001011001111110101;
            sine_reg0   <= 36'sb110001001110101110011101010000100001;
        end
        15134: begin
            cosine_reg0 <= 36'sb11100011001001010010111100010000111;
            sine_reg0   <= 36'sb110001001111011011000011010111010110;
        end
        15135: begin
            cosine_reg0 <= 36'sb11100011001100001100010101110010111;
            sine_reg0   <= 36'sb110001010000000111101010000010100111;
        end
        15136: begin
            cosine_reg0 <= 36'sb11100011001111000101100110100100001;
            sine_reg0   <= 36'sb110001010000110100010001010010010000;
        end
        15137: begin
            cosine_reg0 <= 36'sb11100011010001111110101110100100110;
            sine_reg0   <= 36'sb110001010001100000111001000110010000;
        end
        15138: begin
            cosine_reg0 <= 36'sb11100011010100110111101101110100101;
            sine_reg0   <= 36'sb110001010010001101100001011110100110;
        end
        15139: begin
            cosine_reg0 <= 36'sb11100011010111110000100100010011101;
            sine_reg0   <= 36'sb110001010010111010001010011011001111;
        end
        15140: begin
            cosine_reg0 <= 36'sb11100011011010101001010010000001100;
            sine_reg0   <= 36'sb110001010011100110110011111100001011;
        end
        15141: begin
            cosine_reg0 <= 36'sb11100011011101100001110110111110011;
            sine_reg0   <= 36'sb110001010100010011011110000001010111;
        end
        15142: begin
            cosine_reg0 <= 36'sb11100011100000011010010011001001111;
            sine_reg0   <= 36'sb110001010101000000001000101010110001;
        end
        15143: begin
            cosine_reg0 <= 36'sb11100011100011010010100110100100001;
            sine_reg0   <= 36'sb110001010101101100110011111000011001;
        end
        15144: begin
            cosine_reg0 <= 36'sb11100011100110001010110001001100111;
            sine_reg0   <= 36'sb110001010110011001011111101010001011;
        end
        15145: begin
            cosine_reg0 <= 36'sb11100011101001000010110011000100000;
            sine_reg0   <= 36'sb110001010111000110001100000000000111;
        end
        15146: begin
            cosine_reg0 <= 36'sb11100011101011111010101100001001100;
            sine_reg0   <= 36'sb110001010111110010111000111010001011;
        end
        15147: begin
            cosine_reg0 <= 36'sb11100011101110110010011100011101010;
            sine_reg0   <= 36'sb110001011000011111100110011000010101;
        end
        15148: begin
            cosine_reg0 <= 36'sb11100011110001101010000011111111000;
            sine_reg0   <= 36'sb110001011001001100010100011010100011;
        end
        15149: begin
            cosine_reg0 <= 36'sb11100011110100100001100010101110111;
            sine_reg0   <= 36'sb110001011001111001000011000000110100;
        end
        15150: begin
            cosine_reg0 <= 36'sb11100011110111011000111000101100100;
            sine_reg0   <= 36'sb110001011010100101110010001011000101;
        end
        15151: begin
            cosine_reg0 <= 36'sb11100011111010010000000101110111111;
            sine_reg0   <= 36'sb110001011011010010100001111001010101;
        end
        15152: begin
            cosine_reg0 <= 36'sb11100011111101000111001010010001000;
            sine_reg0   <= 36'sb110001011011111111010010001011100011;
        end
        15153: begin
            cosine_reg0 <= 36'sb11100011111111111110000101110111101;
            sine_reg0   <= 36'sb110001011100101100000011000001101101;
        end
        15154: begin
            cosine_reg0 <= 36'sb11100100000010110100111000101011101;
            sine_reg0   <= 36'sb110001011101011000110100011011110000;
        end
        15155: begin
            cosine_reg0 <= 36'sb11100100000101101011100010101101000;
            sine_reg0   <= 36'sb110001011110000101100110011001101100;
        end
        15156: begin
            cosine_reg0 <= 36'sb11100100001000100010000011111011101;
            sine_reg0   <= 36'sb110001011110110010011000111011011110;
        end
        15157: begin
            cosine_reg0 <= 36'sb11100100001011011000011100010111011;
            sine_reg0   <= 36'sb110001011111011111001100000001000101;
        end
        15158: begin
            cosine_reg0 <= 36'sb11100100001110001110101100000000000;
            sine_reg0   <= 36'sb110001100000001011111111101010011110;
        end
        15159: begin
            cosine_reg0 <= 36'sb11100100010001000100110010110101101;
            sine_reg0   <= 36'sb110001100000111000110011110111101010;
        end
        15160: begin
            cosine_reg0 <= 36'sb11100100010011111010110000111000000;
            sine_reg0   <= 36'sb110001100001100101101000101000100100;
        end
        15161: begin
            cosine_reg0 <= 36'sb11100100010110110000100110000111000;
            sine_reg0   <= 36'sb110001100010010010011101111101001101;
        end
        15162: begin
            cosine_reg0 <= 36'sb11100100011001100110010010100010100;
            sine_reg0   <= 36'sb110001100010111111010011110101100001;
        end
        15163: begin
            cosine_reg0 <= 36'sb11100100011100011011110110001010101;
            sine_reg0   <= 36'sb110001100011101100001010010001100000;
        end
        15164: begin
            cosine_reg0 <= 36'sb11100100011111010001010000111110111;
            sine_reg0   <= 36'sb110001100100011001000001010001001000;
        end
        15165: begin
            cosine_reg0 <= 36'sb11100100100010000110100010111111100;
            sine_reg0   <= 36'sb110001100101000101111000110100010110;
        end
        15166: begin
            cosine_reg0 <= 36'sb11100100100100111011101100001100010;
            sine_reg0   <= 36'sb110001100101110010110000111011001010;
        end
        15167: begin
            cosine_reg0 <= 36'sb11100100100111110000101100100100111;
            sine_reg0   <= 36'sb110001100110011111101001100101100001;
        end
        15168: begin
            cosine_reg0 <= 36'sb11100100101010100101100100001001100;
            sine_reg0   <= 36'sb110001100111001100100010110011011010;
        end
        15169: begin
            cosine_reg0 <= 36'sb11100100101101011010010010111001111;
            sine_reg0   <= 36'sb110001100111111001011100100100110011;
        end
        15170: begin
            cosine_reg0 <= 36'sb11100100110000001110111000110110000;
            sine_reg0   <= 36'sb110001101000100110010110111001101010;
        end
        15171: begin
            cosine_reg0 <= 36'sb11100100110011000011010101111101101;
            sine_reg0   <= 36'sb110001101001010011010001110001111110;
        end
        15172: begin
            cosine_reg0 <= 36'sb11100100110101110111101010010000110;
            sine_reg0   <= 36'sb110001101010000000001101001101101100;
        end
        15173: begin
            cosine_reg0 <= 36'sb11100100111000101011110101101111010;
            sine_reg0   <= 36'sb110001101010101101001001001100110100;
        end
        15174: begin
            cosine_reg0 <= 36'sb11100100111011011111111000011001000;
            sine_reg0   <= 36'sb110001101011011010000101101111010011;
        end
        15175: begin
            cosine_reg0 <= 36'sb11100100111110010011110010001101110;
            sine_reg0   <= 36'sb110001101100000111000010110101000111;
        end
        15176: begin
            cosine_reg0 <= 36'sb11100101000001000111100011001101110;
            sine_reg0   <= 36'sb110001101100110100000000011110010000;
        end
        15177: begin
            cosine_reg0 <= 36'sb11100101000011111011001011011000100;
            sine_reg0   <= 36'sb110001101101100000111110101010101010;
        end
        15178: begin
            cosine_reg0 <= 36'sb11100101000110101110101010101110001;
            sine_reg0   <= 36'sb110001101110001101111101011010010101;
        end
        15179: begin
            cosine_reg0 <= 36'sb11100101001001100010000001001110100;
            sine_reg0   <= 36'sb110001101110111010111100101101001111;
        end
        15180: begin
            cosine_reg0 <= 36'sb11100101001100010101001110111001011;
            sine_reg0   <= 36'sb110001101111100111111100100011010101;
        end
        15181: begin
            cosine_reg0 <= 36'sb11100101001111001000010011101110110;
            sine_reg0   <= 36'sb110001110000010100111100111100100111;
        end
        15182: begin
            cosine_reg0 <= 36'sb11100101010001111011001111101110101;
            sine_reg0   <= 36'sb110001110001000001111101111001000010;
        end
        15183: begin
            cosine_reg0 <= 36'sb11100101010100101110000010111000101;
            sine_reg0   <= 36'sb110001110001101110111111011000100101;
        end
        15184: begin
            cosine_reg0 <= 36'sb11100101010111100000101101001100111;
            sine_reg0   <= 36'sb110001110010011100000001011011001110;
        end
        15185: begin
            cosine_reg0 <= 36'sb11100101011010010011001110101011010;
            sine_reg0   <= 36'sb110001110011001001000100000000111011;
        end
        15186: begin
            cosine_reg0 <= 36'sb11100101011101000101100111010011100;
            sine_reg0   <= 36'sb110001110011110110000111001001101010;
        end
        15187: begin
            cosine_reg0 <= 36'sb11100101011111110111110111000101100;
            sine_reg0   <= 36'sb110001110100100011001010110101011011;
        end
        15188: begin
            cosine_reg0 <= 36'sb11100101100010101001111110000001011;
            sine_reg0   <= 36'sb110001110101010000001111000100001010;
        end
        15189: begin
            cosine_reg0 <= 36'sb11100101100101011011111100000110111;
            sine_reg0   <= 36'sb110001110101111101010011110101110111;
        end
        15190: begin
            cosine_reg0 <= 36'sb11100101101000001101110001010101111;
            sine_reg0   <= 36'sb110001110110101010011001001010011111;
        end
        15191: begin
            cosine_reg0 <= 36'sb11100101101010111111011101101110010;
            sine_reg0   <= 36'sb110001110111010111011111000010000001;
        end
        15192: begin
            cosine_reg0 <= 36'sb11100101101101110001000001001111111;
            sine_reg0   <= 36'sb110001111000000100100101011100011100;
        end
        15193: begin
            cosine_reg0 <= 36'sb11100101110000100010011011111010111;
            sine_reg0   <= 36'sb110001111000110001101100011001101100;
        end
        15194: begin
            cosine_reg0 <= 36'sb11100101110011010011101101101110111;
            sine_reg0   <= 36'sb110001111001011110110011111001110001;
        end
        15195: begin
            cosine_reg0 <= 36'sb11100101110110000100110110101011110;
            sine_reg0   <= 36'sb110001111010001011111011111100101010;
        end
        15196: begin
            cosine_reg0 <= 36'sb11100101111000110101110110110001101;
            sine_reg0   <= 36'sb110001111010111001000100100010010011;
        end
        15197: begin
            cosine_reg0 <= 36'sb11100101111011100110101110000000010;
            sine_reg0   <= 36'sb110001111011100110001101101010101011;
        end
        15198: begin
            cosine_reg0 <= 36'sb11100101111110010111011100010111101;
            sine_reg0   <= 36'sb110001111100010011010111010101110010;
        end
        15199: begin
            cosine_reg0 <= 36'sb11100110000001001000000001110111100;
            sine_reg0   <= 36'sb110001111101000000100001100011100100;
        end
        15200: begin
            cosine_reg0 <= 36'sb11100110000011111000011110011111110;
            sine_reg0   <= 36'sb110001111101101101101100010100000000;
        end
        15201: begin
            cosine_reg0 <= 36'sb11100110000110101000110010010000100;
            sine_reg0   <= 36'sb110001111110011010110111100111000101;
        end
        15202: begin
            cosine_reg0 <= 36'sb11100110001001011000111101001001011;
            sine_reg0   <= 36'sb110001111111001000000011011100110001;
        end
        15203: begin
            cosine_reg0 <= 36'sb11100110001100001000111111001010011;
            sine_reg0   <= 36'sb110001111111110101001111110101000001;
        end
        15204: begin
            cosine_reg0 <= 36'sb11100110001110111000111000010011100;
            sine_reg0   <= 36'sb110010000000100010011100101111110101;
        end
        15205: begin
            cosine_reg0 <= 36'sb11100110010001101000101000100100100;
            sine_reg0   <= 36'sb110010000001001111101010001101001010;
        end
        15206: begin
            cosine_reg0 <= 36'sb11100110010100011000001111111101010;
            sine_reg0   <= 36'sb110010000001111100111000001100111111;
        end
        15207: begin
            cosine_reg0 <= 36'sb11100110010111000111101110011101111;
            sine_reg0   <= 36'sb110010000010101010000110101111010001;
        end
        15208: begin
            cosine_reg0 <= 36'sb11100110011001110111000100000110000;
            sine_reg0   <= 36'sb110010000011010111010101110100000000;
        end
        15209: begin
            cosine_reg0 <= 36'sb11100110011100100110010000110101101;
            sine_reg0   <= 36'sb110010000100000100100101011011001010;
        end
        15210: begin
            cosine_reg0 <= 36'sb11100110011111010101010100101100101;
            sine_reg0   <= 36'sb110010000100110001110101100100101100;
        end
        15211: begin
            cosine_reg0 <= 36'sb11100110100010000100001111101011000;
            sine_reg0   <= 36'sb110010000101011111000110010000100110;
        end
        15212: begin
            cosine_reg0 <= 36'sb11100110100100110011000001110000100;
            sine_reg0   <= 36'sb110010000110001100010111011110110100;
        end
        15213: begin
            cosine_reg0 <= 36'sb11100110100111100001101010111101000;
            sine_reg0   <= 36'sb110010000110111001101001001111010110;
        end
        15214: begin
            cosine_reg0 <= 36'sb11100110101010010000001011010000101;
            sine_reg0   <= 36'sb110010000111100110111011100010001010;
        end
        15215: begin
            cosine_reg0 <= 36'sb11100110101100111110100010101011000;
            sine_reg0   <= 36'sb110010001000010100001110010111001110;
        end
        15216: begin
            cosine_reg0 <= 36'sb11100110101111101100110001001100010;
            sine_reg0   <= 36'sb110010001001000001100001101110100000;
        end
        15217: begin
            cosine_reg0 <= 36'sb11100110110010011010110110110100001;
            sine_reg0   <= 36'sb110010001001101110110101100111111110;
        end
        15218: begin
            cosine_reg0 <= 36'sb11100110110101001000110011100010100;
            sine_reg0   <= 36'sb110010001010011100001010000011101000;
        end
        15219: begin
            cosine_reg0 <= 36'sb11100110110111110110100111010111011;
            sine_reg0   <= 36'sb110010001011001001011111000001011010;
        end
        15220: begin
            cosine_reg0 <= 36'sb11100110111010100100010010010010100;
            sine_reg0   <= 36'sb110010001011110110110100100001010100;
        end
        15221: begin
            cosine_reg0 <= 36'sb11100110111101010001110100010100000;
            sine_reg0   <= 36'sb110010001100100100001010100011010011;
        end
        15222: begin
            cosine_reg0 <= 36'sb11100110111111111111001101011011100;
            sine_reg0   <= 36'sb110010001101010001100001000111010110;
        end
        15223: begin
            cosine_reg0 <= 36'sb11100111000010101100011101101001001;
            sine_reg0   <= 36'sb110010001101111110111000001101011011;
        end
        15224: begin
            cosine_reg0 <= 36'sb11100111000101011001100100111100110;
            sine_reg0   <= 36'sb110010001110101100001111110101100001;
        end
        15225: begin
            cosine_reg0 <= 36'sb11100111001000000110100011010110000;
            sine_reg0   <= 36'sb110010001111011001100111111111100101;
        end
        15226: begin
            cosine_reg0 <= 36'sb11100111001010110011011000110101001;
            sine_reg0   <= 36'sb110010010000000111000000101011100101;
        end
        15227: begin
            cosine_reg0 <= 36'sb11100111001101100000000101011001110;
            sine_reg0   <= 36'sb110010010000110100011001111001100001;
        end
        15228: begin
            cosine_reg0 <= 36'sb11100111010000001100101001000100000;
            sine_reg0   <= 36'sb110010010001100001110011101001010110;
        end
        15229: begin
            cosine_reg0 <= 36'sb11100111010010111001000011110011101;
            sine_reg0   <= 36'sb110010010010001111001101111011000011;
        end
        15230: begin
            cosine_reg0 <= 36'sb11100111010101100101010101101000100;
            sine_reg0   <= 36'sb110010010010111100101000101110100101;
        end
        15231: begin
            cosine_reg0 <= 36'sb11100111011000010001011110100010101;
            sine_reg0   <= 36'sb110010010011101010000100000011111100;
        end
        15232: begin
            cosine_reg0 <= 36'sb11100111011010111101011110100001110;
            sine_reg0   <= 36'sb110010010100010111011111111011000100;
        end
        15233: begin
            cosine_reg0 <= 36'sb11100111011101101001010101100110000;
            sine_reg0   <= 36'sb110010010101000100111100010011111101;
        end
        15234: begin
            cosine_reg0 <= 36'sb11100111100000010101000011101111000;
            sine_reg0   <= 36'sb110010010101110010011001001110100110;
        end
        15235: begin
            cosine_reg0 <= 36'sb11100111100011000000101000111100111;
            sine_reg0   <= 36'sb110010010110011111110110101010111011;
        end
        15236: begin
            cosine_reg0 <= 36'sb11100111100101101100000101001111100;
            sine_reg0   <= 36'sb110010010111001101010100101000111011;
        end
        15237: begin
            cosine_reg0 <= 36'sb11100111101000010111011000100110100;
            sine_reg0   <= 36'sb110010010111111010110011001000100101;
        end
        15238: begin
            cosine_reg0 <= 36'sb11100111101011000010100011000010001;
            sine_reg0   <= 36'sb110010011000101000010010001001110110;
        end
        15239: begin
            cosine_reg0 <= 36'sb11100111101101101101100100100010001;
            sine_reg0   <= 36'sb110010011001010101110001101100101110;
        end
        15240: begin
            cosine_reg0 <= 36'sb11100111110000011000011101000110011;
            sine_reg0   <= 36'sb110010011010000011010001110001001010;
        end
        15241: begin
            cosine_reg0 <= 36'sb11100111110011000011001100101110110;
            sine_reg0   <= 36'sb110010011010110000110010010111001000;
        end
        15242: begin
            cosine_reg0 <= 36'sb11100111110101101101110011011011001;
            sine_reg0   <= 36'sb110010011011011110010011011110101000;
        end
        15243: begin
            cosine_reg0 <= 36'sb11100111111000011000010001001011101;
            sine_reg0   <= 36'sb110010011100001011110101000111100110;
        end
        15244: begin
            cosine_reg0 <= 36'sb11100111111011000010100101111111111;
            sine_reg0   <= 36'sb110010011100111001010111010010000001;
        end
        15245: begin
            cosine_reg0 <= 36'sb11100111111101101100110001110111111;
            sine_reg0   <= 36'sb110010011101100110111001111101111000;
        end
        15246: begin
            cosine_reg0 <= 36'sb11101000000000010110110100110011101;
            sine_reg0   <= 36'sb110010011110010100011101001011001001;
        end
        15247: begin
            cosine_reg0 <= 36'sb11101000000011000000101110110010110;
            sine_reg0   <= 36'sb110010011111000010000000111001110010;
        end
        15248: begin
            cosine_reg0 <= 36'sb11101000000101101010011111110101100;
            sine_reg0   <= 36'sb110010011111101111100101001001110001;
        end
        15249: begin
            cosine_reg0 <= 36'sb11101000001000010100000111111011100;
            sine_reg0   <= 36'sb110010100000011101001001111011000100;
        end
        15250: begin
            cosine_reg0 <= 36'sb11101000001010111101100111000100110;
            sine_reg0   <= 36'sb110010100001001010101111001101101010;
        end
        15251: begin
            cosine_reg0 <= 36'sb11101000001101100110111101010001001;
            sine_reg0   <= 36'sb110010100001111000010101000001100001;
        end
        15252: begin
            cosine_reg0 <= 36'sb11101000010000010000001010100000101;
            sine_reg0   <= 36'sb110010100010100101111011010110100111;
        end
        15253: begin
            cosine_reg0 <= 36'sb11101000010010111001001110110011000;
            sine_reg0   <= 36'sb110010100011010011100010001100111011;
        end
        15254: begin
            cosine_reg0 <= 36'sb11101000010101100010001010001000001;
            sine_reg0   <= 36'sb110010100100000001001001100100011010;
        end
        15255: begin
            cosine_reg0 <= 36'sb11101000011000001010111100100000001;
            sine_reg0   <= 36'sb110010100100101110110001011101000011;
        end
        15256: begin
            cosine_reg0 <= 36'sb11101000011010110011100101111010110;
            sine_reg0   <= 36'sb110010100101011100011001110110110101;
        end
        15257: begin
            cosine_reg0 <= 36'sb11101000011101011100000110010111110;
            sine_reg0   <= 36'sb110010100110001010000010110001101101;
        end
        15258: begin
            cosine_reg0 <= 36'sb11101000100000000100011101110111011;
            sine_reg0   <= 36'sb110010100110110111101100001101101001;
        end
        15259: begin
            cosine_reg0 <= 36'sb11101000100010101100101100011001001;
            sine_reg0   <= 36'sb110010100111100101010110001010101000;
        end
        15260: begin
            cosine_reg0 <= 36'sb11101000100101010100110001111101010;
            sine_reg0   <= 36'sb110010101000010011000000101000101001;
        end
        15261: begin
            cosine_reg0 <= 36'sb11101000100111111100101110100011100;
            sine_reg0   <= 36'sb110010101001000000101011100111101001;
        end
        15262: begin
            cosine_reg0 <= 36'sb11101000101010100100100010001011110;
            sine_reg0   <= 36'sb110010101001101110010111000111100110;
        end
        15263: begin
            cosine_reg0 <= 36'sb11101000101101001100001100110101111;
            sine_reg0   <= 36'sb110010101010011100000011001000011111;
        end
        15264: begin
            cosine_reg0 <= 36'sb11101000101111110011101110100001111;
            sine_reg0   <= 36'sb110010101011001001101111101010010011;
        end
        15265: begin
            cosine_reg0 <= 36'sb11101000110010011011000111001111100;
            sine_reg0   <= 36'sb110010101011110111011100101100111110;
        end
        15266: begin
            cosine_reg0 <= 36'sb11101000110101000010010110111110111;
            sine_reg0   <= 36'sb110010101100100101001010010000100001;
        end
        15267: begin
            cosine_reg0 <= 36'sb11101000110111101001011101101111101;
            sine_reg0   <= 36'sb110010101101010010111000010100111000;
        end
        15268: begin
            cosine_reg0 <= 36'sb11101000111010010000011011100001111;
            sine_reg0   <= 36'sb110010101110000000100110111010000010;
        end
        15269: begin
            cosine_reg0 <= 36'sb11101000111100110111010000010101100;
            sine_reg0   <= 36'sb110010101110101110010101111111111101;
        end
        15270: begin
            cosine_reg0 <= 36'sb11101000111111011101111100001010010;
            sine_reg0   <= 36'sb110010101111011100000101100110101000;
        end
        15271: begin
            cosine_reg0 <= 36'sb11101001000010000100011111000000001;
            sine_reg0   <= 36'sb110010110000001001110101101110000000;
        end
        15272: begin
            cosine_reg0 <= 36'sb11101001000100101010111000110111001;
            sine_reg0   <= 36'sb110010110000110111100110010110000101;
        end
        15273: begin
            cosine_reg0 <= 36'sb11101001000111010001001001101110111;
            sine_reg0   <= 36'sb110010110001100101010111011110110100;
        end
        15274: begin
            cosine_reg0 <= 36'sb11101001001001110111010001100111100;
            sine_reg0   <= 36'sb110010110010010011001001001000001011;
        end
        15275: begin
            cosine_reg0 <= 36'sb11101001001100011101010000100000111;
            sine_reg0   <= 36'sb110010110011000000111011010010001001;
        end
        15276: begin
            cosine_reg0 <= 36'sb11101001001111000011000110011010111;
            sine_reg0   <= 36'sb110010110011101110101101111100101100;
        end
        15277: begin
            cosine_reg0 <= 36'sb11101001010001101000110011010101011;
            sine_reg0   <= 36'sb110010110100011100100001000111110001;
        end
        15278: begin
            cosine_reg0 <= 36'sb11101001010100001110010111010000010;
            sine_reg0   <= 36'sb110010110101001010010100110011011001;
        end
        15279: begin
            cosine_reg0 <= 36'sb11101001010110110011110010001011100;
            sine_reg0   <= 36'sb110010110101111000001000111111100000;
        end
        15280: begin
            cosine_reg0 <= 36'sb11101001011001011001000100000110111;
            sine_reg0   <= 36'sb110010110110100101111101101100000101;
        end
        15281: begin
            cosine_reg0 <= 36'sb11101001011011111110001101000010100;
            sine_reg0   <= 36'sb110010110111010011110010111001000101;
        end
        15282: begin
            cosine_reg0 <= 36'sb11101001011110100011001100111110000;
            sine_reg0   <= 36'sb110010111000000001101000100110100001;
        end
        15283: begin
            cosine_reg0 <= 36'sb11101001100001001000000011111001100;
            sine_reg0   <= 36'sb110010111000101111011110110100010100;
        end
        15284: begin
            cosine_reg0 <= 36'sb11101001100011101100110001110100111;
            sine_reg0   <= 36'sb110010111001011101010101100010011111;
        end
        15285: begin
            cosine_reg0 <= 36'sb11101001100110010001010110101111111;
            sine_reg0   <= 36'sb110010111010001011001100110000111111;
        end
        15286: begin
            cosine_reg0 <= 36'sb11101001101000110101110010101010100;
            sine_reg0   <= 36'sb110010111010111001000100011111110001;
        end
        15287: begin
            cosine_reg0 <= 36'sb11101001101011011010000101100100101;
            sine_reg0   <= 36'sb110010111011100110111100101110110110;
        end
        15288: begin
            cosine_reg0 <= 36'sb11101001101101111110001111011110010;
            sine_reg0   <= 36'sb110010111100010100110101011110001010;
        end
        15289: begin
            cosine_reg0 <= 36'sb11101001110000100010010000010111001;
            sine_reg0   <= 36'sb110010111101000010101110101101101100;
        end
        15290: begin
            cosine_reg0 <= 36'sb11101001110011000110001000001111010;
            sine_reg0   <= 36'sb110010111101110000101000011101011010;
        end
        15291: begin
            cosine_reg0 <= 36'sb11101001110101101001110111000110101;
            sine_reg0   <= 36'sb110010111110011110100010101101010010;
        end
        15292: begin
            cosine_reg0 <= 36'sb11101001111000001101011100111100111;
            sine_reg0   <= 36'sb110010111111001100011101011101010100;
        end
        15293: begin
            cosine_reg0 <= 36'sb11101001111010110000111001110010001;
            sine_reg0   <= 36'sb110010111111111010011000101101011100;
        end
        15294: begin
            cosine_reg0 <= 36'sb11101001111101010100001101100110001;
            sine_reg0   <= 36'sb110011000000101000010100011101101001;
        end
        15295: begin
            cosine_reg0 <= 36'sb11101001111111110111011000011000111;
            sine_reg0   <= 36'sb110011000001010110010000101101111001;
        end
        15296: begin
            cosine_reg0 <= 36'sb11101010000010011010011010001010011;
            sine_reg0   <= 36'sb110011000010000100001101011110001011;
        end
        15297: begin
            cosine_reg0 <= 36'sb11101010000100111101010010111010010;
            sine_reg0   <= 36'sb110011000010110010001010101110011101;
        end
        15298: begin
            cosine_reg0 <= 36'sb11101010000111100000000010101000101;
            sine_reg0   <= 36'sb110011000011100000001000011110101101;
        end
        15299: begin
            cosine_reg0 <= 36'sb11101010001010000010101001010101011;
            sine_reg0   <= 36'sb110011000100001110000110101110111001;
        end
        15300: begin
            cosine_reg0 <= 36'sb11101010001100100101000111000000011;
            sine_reg0   <= 36'sb110011000100111100000101011110111111;
        end
        15301: begin
            cosine_reg0 <= 36'sb11101010001111000111011011101001100;
            sine_reg0   <= 36'sb110011000101101010000100101110111111;
        end
        15302: begin
            cosine_reg0 <= 36'sb11101010010001101001100111010000101;
            sine_reg0   <= 36'sb110011000110011000000100011110110101;
        end
        15303: begin
            cosine_reg0 <= 36'sb11101010010100001011101001110101110;
            sine_reg0   <= 36'sb110011000111000110000100101110100000;
        end
        15304: begin
            cosine_reg0 <= 36'sb11101010010110101101100011011000101;
            sine_reg0   <= 36'sb110011000111110100000101011101111111;
        end
        15305: begin
            cosine_reg0 <= 36'sb11101010011001001111010011111001011;
            sine_reg0   <= 36'sb110011001000100010000110101101001111;
        end
        15306: begin
            cosine_reg0 <= 36'sb11101010011011110000111011010111110;
            sine_reg0   <= 36'sb110011001001010000001000011100001111;
        end
        15307: begin
            cosine_reg0 <= 36'sb11101010011110010010011001110011101;
            sine_reg0   <= 36'sb110011001001111110001010101010111101;
        end
        15308: begin
            cosine_reg0 <= 36'sb11101010100000110011101111001101000;
            sine_reg0   <= 36'sb110011001010101100001101011001010111;
        end
        15309: begin
            cosine_reg0 <= 36'sb11101010100011010100111011100011110;
            sine_reg0   <= 36'sb110011001011011010010000100111011100;
        end
        15310: begin
            cosine_reg0 <= 36'sb11101010100101110101111110110111110;
            sine_reg0   <= 36'sb110011001100001000010100010101001010;
        end
        15311: begin
            cosine_reg0 <= 36'sb11101010101000010110111001001000111;
            sine_reg0   <= 36'sb110011001100110110011000100010011110;
        end
        15312: begin
            cosine_reg0 <= 36'sb11101010101010110111101010010111001;
            sine_reg0   <= 36'sb110011001101100100011101001111011000;
        end
        15313: begin
            cosine_reg0 <= 36'sb11101010101101011000010010100010011;
            sine_reg0   <= 36'sb110011001110010010100010011011110101;
        end
        15314: begin
            cosine_reg0 <= 36'sb11101010101111111000110001101010100;
            sine_reg0   <= 36'sb110011001111000000101000000111110100;
        end
        15315: begin
            cosine_reg0 <= 36'sb11101010110010011001000111101111011;
            sine_reg0   <= 36'sb110011001111101110101110010011010011;
        end
        15316: begin
            cosine_reg0 <= 36'sb11101010110100111001010100110001000;
            sine_reg0   <= 36'sb110011010000011100110100111110001111;
        end
        15317: begin
            cosine_reg0 <= 36'sb11101010110111011001011000101111001;
            sine_reg0   <= 36'sb110011010001001010111100001000101000;
        end
        15318: begin
            cosine_reg0 <= 36'sb11101010111001111001010011101001110;
            sine_reg0   <= 36'sb110011010001111001000011110010011100;
        end
        15319: begin
            cosine_reg0 <= 36'sb11101010111100011001000101100000110;
            sine_reg0   <= 36'sb110011010010100111001011111011101000;
        end
        15320: begin
            cosine_reg0 <= 36'sb11101010111110111000101110010100001;
            sine_reg0   <= 36'sb110011010011010101010100100100001011;
        end
        15321: begin
            cosine_reg0 <= 36'sb11101011000001011000001110000011110;
            sine_reg0   <= 36'sb110011010100000011011101101100000011;
        end
        15322: begin
            cosine_reg0 <= 36'sb11101011000011110111100100101111011;
            sine_reg0   <= 36'sb110011010100110001100111010011001111;
        end
        15323: begin
            cosine_reg0 <= 36'sb11101011000110010110110010010111000;
            sine_reg0   <= 36'sb110011010101011111110001011001101100;
        end
        15324: begin
            cosine_reg0 <= 36'sb11101011001000110101110110111010101;
            sine_reg0   <= 36'sb110011010110001101111011111111011001;
        end
        15325: begin
            cosine_reg0 <= 36'sb11101011001011010100110010011010000;
            sine_reg0   <= 36'sb110011010110111100000111000100010101;
        end
        15326: begin
            cosine_reg0 <= 36'sb11101011001101110011100100110101001;
            sine_reg0   <= 36'sb110011010111101010010010101000011100;
        end
        15327: begin
            cosine_reg0 <= 36'sb11101011010000010010001110001011111;
            sine_reg0   <= 36'sb110011011000011000011110101011101110;
        end
        15328: begin
            cosine_reg0 <= 36'sb11101011010010110000101110011110010;
            sine_reg0   <= 36'sb110011011001000110101011001110001001;
        end
        15329: begin
            cosine_reg0 <= 36'sb11101011010101001111000101101011111;
            sine_reg0   <= 36'sb110011011001110100111000001111101010;
        end
        15330: begin
            cosine_reg0 <= 36'sb11101011010111101101010011110101000;
            sine_reg0   <= 36'sb110011011010100011000101110000010001;
        end
        15331: begin
            cosine_reg0 <= 36'sb11101011011010001011011000111001010;
            sine_reg0   <= 36'sb110011011011010001010011101111111011;
        end
        15332: begin
            cosine_reg0 <= 36'sb11101011011100101001010100111000110;
            sine_reg0   <= 36'sb110011011011111111100010001110100111;
        end
        15333: begin
            cosine_reg0 <= 36'sb11101011011111000111000111110011010;
            sine_reg0   <= 36'sb110011011100101101110001001100010011;
        end
        15334: begin
            cosine_reg0 <= 36'sb11101011100001100100110001101000110;
            sine_reg0   <= 36'sb110011011101011100000000101000111100;
        end
        15335: begin
            cosine_reg0 <= 36'sb11101011100100000010010010011001001;
            sine_reg0   <= 36'sb110011011110001010010000100100100010;
        end
        15336: begin
            cosine_reg0 <= 36'sb11101011100110011111101010000100010;
            sine_reg0   <= 36'sb110011011110111000100000111111000010;
        end
        15337: begin
            cosine_reg0 <= 36'sb11101011101000111100111000101010000;
            sine_reg0   <= 36'sb110011011111100110110001111000011011;
        end
        15338: begin
            cosine_reg0 <= 36'sb11101011101011011001111110001010100;
            sine_reg0   <= 36'sb110011100000010101000011010000101011;
        end
        15339: begin
            cosine_reg0 <= 36'sb11101011101101110110111010100101011;
            sine_reg0   <= 36'sb110011100001000011010101000111110000;
        end
        15340: begin
            cosine_reg0 <= 36'sb11101011110000010011101101111010101;
            sine_reg0   <= 36'sb110011100001110001100111011101101001;
        end
        15341: begin
            cosine_reg0 <= 36'sb11101011110010110000011000001010001;
            sine_reg0   <= 36'sb110011100010011111111010010010010010;
        end
        15342: begin
            cosine_reg0 <= 36'sb11101011110101001100111001010011111;
            sine_reg0   <= 36'sb110011100011001110001101100101101100;
        end
        15343: begin
            cosine_reg0 <= 36'sb11101011110111101001010001010111110;
            sine_reg0   <= 36'sb110011100011111100100001010111110100;
        end
        15344: begin
            cosine_reg0 <= 36'sb11101011111010000101100000010101101;
            sine_reg0   <= 36'sb110011100100101010110101101000100111;
        end
        15345: begin
            cosine_reg0 <= 36'sb11101011111100100001100110001101100;
            sine_reg0   <= 36'sb110011100101011001001010011000000101;
        end
        15346: begin
            cosine_reg0 <= 36'sb11101011111110111101100010111111001;
            sine_reg0   <= 36'sb110011100110000111011111100110001100;
        end
        15347: begin
            cosine_reg0 <= 36'sb11101100000001011001010110101010100;
            sine_reg0   <= 36'sb110011100110110101110101010010111010;
        end
        15348: begin
            cosine_reg0 <= 36'sb11101100000011110101000001001111100;
            sine_reg0   <= 36'sb110011100111100100001011011110001100;
        end
        15349: begin
            cosine_reg0 <= 36'sb11101100000110010000100010101110000;
            sine_reg0   <= 36'sb110011101000010010100010001000000010;
        end
        15350: begin
            cosine_reg0 <= 36'sb11101100001000101011111011000110000;
            sine_reg0   <= 36'sb110011101001000000111001010000011010;
        end
        15351: begin
            cosine_reg0 <= 36'sb11101100001011000111001010010111011;
            sine_reg0   <= 36'sb110011101001101111010000110111010001;
        end
        15352: begin
            cosine_reg0 <= 36'sb11101100001101100010010000100010000;
            sine_reg0   <= 36'sb110011101010011101101000111100100110;
        end
        15353: begin
            cosine_reg0 <= 36'sb11101100001111111101001101100101111;
            sine_reg0   <= 36'sb110011101011001100000001100000010111;
        end
        15354: begin
            cosine_reg0 <= 36'sb11101100010010011000000001100010110;
            sine_reg0   <= 36'sb110011101011111010011010100010100010;
        end
        15355: begin
            cosine_reg0 <= 36'sb11101100010100110010101100011000101;
            sine_reg0   <= 36'sb110011101100101000110100000011000110;
        end
        15356: begin
            cosine_reg0 <= 36'sb11101100010111001101001110000111011;
            sine_reg0   <= 36'sb110011101101010111001110000010000001;
        end
        15357: begin
            cosine_reg0 <= 36'sb11101100011001100111100110101110111;
            sine_reg0   <= 36'sb110011101110000101101000011111010000;
        end
        15358: begin
            cosine_reg0 <= 36'sb11101100011100000001110110001111010;
            sine_reg0   <= 36'sb110011101110110100000011011010110011;
        end
        15359: begin
            cosine_reg0 <= 36'sb11101100011110011011111100101000001;
            sine_reg0   <= 36'sb110011101111100010011110110100100111;
        end
        15360: begin
            cosine_reg0 <= 36'sb11101100100000110101111001111001100;
            sine_reg0   <= 36'sb110011110000010000111010101100101011;
        end
        15361: begin
            cosine_reg0 <= 36'sb11101100100011001111101110000011010;
            sine_reg0   <= 36'sb110011110000111111010111000010111100;
        end
        15362: begin
            cosine_reg0 <= 36'sb11101100100101101001011001000101100;
            sine_reg0   <= 36'sb110011110001101101110011110111011001;
        end
        15363: begin
            cosine_reg0 <= 36'sb11101100101000000010111010111111111;
            sine_reg0   <= 36'sb110011110010011100010001001010000001;
        end
        15364: begin
            cosine_reg0 <= 36'sb11101100101010011100010011110010011;
            sine_reg0   <= 36'sb110011110011001010101110111010110001;
        end
        15365: begin
            cosine_reg0 <= 36'sb11101100101100110101100011011101000;
            sine_reg0   <= 36'sb110011110011111001001101001001101000;
        end
        15366: begin
            cosine_reg0 <= 36'sb11101100101111001110101001111111101;
            sine_reg0   <= 36'sb110011110100100111101011110110100011;
        end
        15367: begin
            cosine_reg0 <= 36'sb11101100110001100111100111011010000;
            sine_reg0   <= 36'sb110011110101010110001011000001100010;
        end
        15368: begin
            cosine_reg0 <= 36'sb11101100110100000000011011101100010;
            sine_reg0   <= 36'sb110011110110000100101010101010100010;
        end
        15369: begin
            cosine_reg0 <= 36'sb11101100110110011001000110110110001;
            sine_reg0   <= 36'sb110011110110110011001010110001100001;
        end
        15370: begin
            cosine_reg0 <= 36'sb11101100111000110001101000110111101;
            sine_reg0   <= 36'sb110011110111100001101011010110011110;
        end
        15371: begin
            cosine_reg0 <= 36'sb11101100111011001010000001110000101;
            sine_reg0   <= 36'sb110011111000010000001100011001010111;
        end
        15372: begin
            cosine_reg0 <= 36'sb11101100111101100010010001100001001;
            sine_reg0   <= 36'sb110011111000111110101101111010001010;
        end
        15373: begin
            cosine_reg0 <= 36'sb11101100111111111010011000001000111;
            sine_reg0   <= 36'sb110011111001101101001111111000110101;
        end
        15374: begin
            cosine_reg0 <= 36'sb11101101000010010010010101100111111;
            sine_reg0   <= 36'sb110011111010011011110010010101010111;
        end
        15375: begin
            cosine_reg0 <= 36'sb11101101000100101010001001111101111;
            sine_reg0   <= 36'sb110011111011001010010101001111101101;
        end
        15376: begin
            cosine_reg0 <= 36'sb11101101000111000001110101001011001;
            sine_reg0   <= 36'sb110011111011111000111000100111110111;
        end
        15377: begin
            cosine_reg0 <= 36'sb11101101001001011001010111001111010;
            sine_reg0   <= 36'sb110011111100100111011100011101110001;
        end
        15378: begin
            cosine_reg0 <= 36'sb11101101001011110000110000001010001;
            sine_reg0   <= 36'sb110011111101010110000000110001011011;
        end
        15379: begin
            cosine_reg0 <= 36'sb11101101001110000111111111111011111;
            sine_reg0   <= 36'sb110011111110000100100101100010110010;
        end
        15380: begin
            cosine_reg0 <= 36'sb11101101010000011111000110100100011;
            sine_reg0   <= 36'sb110011111110110011001010110001110101;
        end
        15381: begin
            cosine_reg0 <= 36'sb11101101010010110110000100000011011;
            sine_reg0   <= 36'sb110011111111100001110000011110100010;
        end
        15382: begin
            cosine_reg0 <= 36'sb11101101010101001100111000011000111;
            sine_reg0   <= 36'sb110100000000010000010110101000110111;
        end
        15383: begin
            cosine_reg0 <= 36'sb11101101010111100011100011100100111;
            sine_reg0   <= 36'sb110100000000111110111101010000110010;
        end
        15384: begin
            cosine_reg0 <= 36'sb11101101011001111010000101100111001;
            sine_reg0   <= 36'sb110100000001101101100100010110010010;
        end
        15385: begin
            cosine_reg0 <= 36'sb11101101011100010000011110011111101;
            sine_reg0   <= 36'sb110100000010011100001011111001010101;
        end
        15386: begin
            cosine_reg0 <= 36'sb11101101011110100110101110001110001;
            sine_reg0   <= 36'sb110100000011001010110011111001111000;
        end
        15387: begin
            cosine_reg0 <= 36'sb11101101100000111100110100110010111;
            sine_reg0   <= 36'sb110100000011111001011100010111111011;
        end
        15388: begin
            cosine_reg0 <= 36'sb11101101100011010010110010001101100;
            sine_reg0   <= 36'sb110100000100101000000101010011011011;
        end
        15389: begin
            cosine_reg0 <= 36'sb11101101100101101000100110011101111;
            sine_reg0   <= 36'sb110100000101010110101110101100010111;
        end
        15390: begin
            cosine_reg0 <= 36'sb11101101100111111110010001100100001;
            sine_reg0   <= 36'sb110100000110000101011000100010101100;
        end
        15391: begin
            cosine_reg0 <= 36'sb11101101101010010011110011100000001;
            sine_reg0   <= 36'sb110100000110110100000010110110011001;
        end
        15392: begin
            cosine_reg0 <= 36'sb11101101101100101001001100010001101;
            sine_reg0   <= 36'sb110100000111100010101101100111011101;
        end
        15393: begin
            cosine_reg0 <= 36'sb11101101101110111110011011111000110;
            sine_reg0   <= 36'sb110100001000010001011000110101110100;
        end
        15394: begin
            cosine_reg0 <= 36'sb11101101110001010011100010010101001;
            sine_reg0   <= 36'sb110100001001000000000100100001011111;
        end
        15395: begin
            cosine_reg0 <= 36'sb11101101110011101000011111100110111;
            sine_reg0   <= 36'sb110100001001101110110000101010011010;
        end
        15396: begin
            cosine_reg0 <= 36'sb11101101110101111101010011101110000;
            sine_reg0   <= 36'sb110100001010011101011101010000100100;
        end
        15397: begin
            cosine_reg0 <= 36'sb11101101111000010001111110101010001;
            sine_reg0   <= 36'sb110100001011001100001010010011111011;
        end
        15398: begin
            cosine_reg0 <= 36'sb11101101111010100110100000011011011;
            sine_reg0   <= 36'sb110100001011111010110111110100011110;
        end
        15399: begin
            cosine_reg0 <= 36'sb11101101111100111010111001000001100;
            sine_reg0   <= 36'sb110100001100101001100101110010001010;
        end
        15400: begin
            cosine_reg0 <= 36'sb11101101111111001111001000011100100;
            sine_reg0   <= 36'sb110100001101011000010100001100111110;
        end
        15401: begin
            cosine_reg0 <= 36'sb11101110000001100011001110101100011;
            sine_reg0   <= 36'sb110100001110000111000011000100111000;
        end
        15402: begin
            cosine_reg0 <= 36'sb11101110000011110111001011110001000;
            sine_reg0   <= 36'sb110100001110110101110010011001110110;
        end
        15403: begin
            cosine_reg0 <= 36'sb11101110000110001010111111101010001;
            sine_reg0   <= 36'sb110100001111100100100010001011110110;
        end
        15404: begin
            cosine_reg0 <= 36'sb11101110001000011110101010010111110;
            sine_reg0   <= 36'sb110100010000010011010010011010110111;
        end
        15405: begin
            cosine_reg0 <= 36'sb11101110001010110010001011111001111;
            sine_reg0   <= 36'sb110100010001000010000011000110110111;
        end
        15406: begin
            cosine_reg0 <= 36'sb11101110001101000101100100010000011;
            sine_reg0   <= 36'sb110100010001110000110100001111110011;
        end
        15407: begin
            cosine_reg0 <= 36'sb11101110001111011000110011011011000;
            sine_reg0   <= 36'sb110100010010011111100101110101101011;
        end
        15408: begin
            cosine_reg0 <= 36'sb11101110010001101011111001011001111;
            sine_reg0   <= 36'sb110100010011001110010111111000011100;
        end
        15409: begin
            cosine_reg0 <= 36'sb11101110010011111110110110001100111;
            sine_reg0   <= 36'sb110100010011111101001010011000000100;
        end
        15410: begin
            cosine_reg0 <= 36'sb11101110010110010001101001110011110;
            sine_reg0   <= 36'sb110100010100101011111101010100100011;
        end
        15411: begin
            cosine_reg0 <= 36'sb11101110011000100100010100001110101;
            sine_reg0   <= 36'sb110100010101011010110000101101110101;
        end
        15412: begin
            cosine_reg0 <= 36'sb11101110011010110110110101011101010;
            sine_reg0   <= 36'sb110100010110001001100100100011111001;
        end
        15413: begin
            cosine_reg0 <= 36'sb11101110011101001001001101011111101;
            sine_reg0   <= 36'sb110100010110111000011000110110101110;
        end
        15414: begin
            cosine_reg0 <= 36'sb11101110011111011011011100010101101;
            sine_reg0   <= 36'sb110100010111100111001101100110010001;
        end
        15415: begin
            cosine_reg0 <= 36'sb11101110100001101101100001111111010;
            sine_reg0   <= 36'sb110100011000010110000010110010100001;
        end
        15416: begin
            cosine_reg0 <= 36'sb11101110100011111111011110011100010;
            sine_reg0   <= 36'sb110100011001000100111000011011011100;
        end
        15417: begin
            cosine_reg0 <= 36'sb11101110100110010001010001101100101;
            sine_reg0   <= 36'sb110100011001110011101110100000111111;
        end
        15418: begin
            cosine_reg0 <= 36'sb11101110101000100010111011110000010;
            sine_reg0   <= 36'sb110100011010100010100101000011001011;
        end
        15419: begin
            cosine_reg0 <= 36'sb11101110101010110100011100100111001;
            sine_reg0   <= 36'sb110100011011010001011100000001111011;
        end
        15420: begin
            cosine_reg0 <= 36'sb11101110101101000101110100010001001;
            sine_reg0   <= 36'sb110100011100000000010011011101001111;
        end
        15421: begin
            cosine_reg0 <= 36'sb11101110101111010111000010101110001;
            sine_reg0   <= 36'sb110100011100101111001011010101000110;
        end
        15422: begin
            cosine_reg0 <= 36'sb11101110110001101000000111111110000;
            sine_reg0   <= 36'sb110100011101011110000011101001011100;
        end
        15423: begin
            cosine_reg0 <= 36'sb11101110110011111001000100000000110;
            sine_reg0   <= 36'sb110100011110001100111100011010010000;
        end
        15424: begin
            cosine_reg0 <= 36'sb11101110110110001001110110110110010;
            sine_reg0   <= 36'sb110100011110111011110101100111100001;
        end
        15425: begin
            cosine_reg0 <= 36'sb11101110111000011010100000011110100;
            sine_reg0   <= 36'sb110100011111101010101111010001001101;
        end
        15426: begin
            cosine_reg0 <= 36'sb11101110111010101011000000111001010;
            sine_reg0   <= 36'sb110100100000011001101001010111010001;
        end
        15427: begin
            cosine_reg0 <= 36'sb11101110111100111011011000000110100;
            sine_reg0   <= 36'sb110100100001001000100011111001101100;
        end
        15428: begin
            cosine_reg0 <= 36'sb11101110111111001011100110000110010;
            sine_reg0   <= 36'sb110100100001110111011110111000011101;
        end
        15429: begin
            cosine_reg0 <= 36'sb11101111000001011011101010111000010;
            sine_reg0   <= 36'sb110100100010100110011010010011100001;
        end
        15430: begin
            cosine_reg0 <= 36'sb11101111000011101011100110011100100;
            sine_reg0   <= 36'sb110100100011010101010110001010110110;
        end
        15431: begin
            cosine_reg0 <= 36'sb11101111000101111011011000110010111;
            sine_reg0   <= 36'sb110100100100000100010010011110011100;
        end
        15432: begin
            cosine_reg0 <= 36'sb11101111001000001011000001111011010;
            sine_reg0   <= 36'sb110100100100110011001111001110001111;
        end
        15433: begin
            cosine_reg0 <= 36'sb11101111001010011010100001110101110;
            sine_reg0   <= 36'sb110100100101100010001100011010001111;
        end
        15434: begin
            cosine_reg0 <= 36'sb11101111001100101001111000100010000;
            sine_reg0   <= 36'sb110100100110010001001010000010011000;
        end
        15435: begin
            cosine_reg0 <= 36'sb11101111001110111001000110000000001;
            sine_reg0   <= 36'sb110100100111000000001000000110101011;
        end
        15436: begin
            cosine_reg0 <= 36'sb11101111010001001000001010010000000;
            sine_reg0   <= 36'sb110100100111101111000110100111000100;
        end
        15437: begin
            cosine_reg0 <= 36'sb11101111010011010111000101010001100;
            sine_reg0   <= 36'sb110100101000011110000101100011100010;
        end
        15438: begin
            cosine_reg0 <= 36'sb11101111010101100101110111000100100;
            sine_reg0   <= 36'sb110100101001001101000100111100000011;
        end
        15439: begin
            cosine_reg0 <= 36'sb11101111010111110100011111101001000;
            sine_reg0   <= 36'sb110100101001111100000100110000100110;
        end
        15440: begin
            cosine_reg0 <= 36'sb11101111011010000010111110111110111;
            sine_reg0   <= 36'sb110100101010101011000101000001000111;
        end
        15441: begin
            cosine_reg0 <= 36'sb11101111011100010001010101000110000;
            sine_reg0   <= 36'sb110100101011011010000101101101100111;
        end
        15442: begin
            cosine_reg0 <= 36'sb11101111011110011111100001111110010;
            sine_reg0   <= 36'sb110100101100001001000110110110000010;
        end
        15443: begin
            cosine_reg0 <= 36'sb11101111100000101101100101100111110;
            sine_reg0   <= 36'sb110100101100111000001000011010011000;
        end
        15444: begin
            cosine_reg0 <= 36'sb11101111100010111011100000000010010;
            sine_reg0   <= 36'sb110100101101100111001010011010100110;
        end
        15445: begin
            cosine_reg0 <= 36'sb11101111100101001001010001001101101;
            sine_reg0   <= 36'sb110100101110010110001100110110101010;
        end
        15446: begin
            cosine_reg0 <= 36'sb11101111100111010110111001001010000;
            sine_reg0   <= 36'sb110100101111000101001111101110100011;
        end
        15447: begin
            cosine_reg0 <= 36'sb11101111101001100100010111110111000;
            sine_reg0   <= 36'sb110100101111110100010011000010001110;
        end
        15448: begin
            cosine_reg0 <= 36'sb11101111101011110001101101010100110;
            sine_reg0   <= 36'sb110100110000100011010110110001101011;
        end
        15449: begin
            cosine_reg0 <= 36'sb11101111101101111110111001100011001;
            sine_reg0   <= 36'sb110100110001010010011010111100110110;
        end
        15450: begin
            cosine_reg0 <= 36'sb11101111110000001011111100100010000;
            sine_reg0   <= 36'sb110100110010000001011111100011101111;
        end
        15451: begin
            cosine_reg0 <= 36'sb11101111110010011000110110010001010;
            sine_reg0   <= 36'sb110100110010110000100100100110010100;
        end
        15452: begin
            cosine_reg0 <= 36'sb11101111110100100101100110110000111;
            sine_reg0   <= 36'sb110100110011011111101010000100100010;
        end
        15453: begin
            cosine_reg0 <= 36'sb11101111110110110010001110000000111;
            sine_reg0   <= 36'sb110100110100001110101111111110011001;
        end
        15454: begin
            cosine_reg0 <= 36'sb11101111111000111110101100000000111;
            sine_reg0   <= 36'sb110100110100111101110110010011110101;
        end
        15455: begin
            cosine_reg0 <= 36'sb11101111111011001011000000110001001;
            sine_reg0   <= 36'sb110100110101101100111101000100110101;
        end
        15456: begin
            cosine_reg0 <= 36'sb11101111111101010111001100010001010;
            sine_reg0   <= 36'sb110100110110011100000100010001011000;
        end
        15457: begin
            cosine_reg0 <= 36'sb11101111111111100011001110100001011;
            sine_reg0   <= 36'sb110100110111001011001011111001011100;
        end
        15458: begin
            cosine_reg0 <= 36'sb11110000000001101111000111100001011;
            sine_reg0   <= 36'sb110100110111111010010011111100111111;
        end
        15459: begin
            cosine_reg0 <= 36'sb11110000000011111010110111010001001;
            sine_reg0   <= 36'sb110100111000101001011100011011111110;
        end
        15460: begin
            cosine_reg0 <= 36'sb11110000000110000110011101110000100;
            sine_reg0   <= 36'sb110100111001011000100101010110011001;
        end
        15461: begin
            cosine_reg0 <= 36'sb11110000001000010001111010111111100;
            sine_reg0   <= 36'sb110100111010000111101110101100001101;
        end
        15462: begin
            cosine_reg0 <= 36'sb11110000001010011101001110111110000;
            sine_reg0   <= 36'sb110100111010110110111000011101011001;
        end
        15463: begin
            cosine_reg0 <= 36'sb11110000001100101000011001101011111;
            sine_reg0   <= 36'sb110100111011100110000010101001111010;
        end
        15464: begin
            cosine_reg0 <= 36'sb11110000001110110011011011001001001;
            sine_reg0   <= 36'sb110100111100010101001101010001101111;
        end
        15465: begin
            cosine_reg0 <= 36'sb11110000010000111110010011010101101;
            sine_reg0   <= 36'sb110100111101000100011000010100110111;
        end
        15466: begin
            cosine_reg0 <= 36'sb11110000010011001001000010010001010;
            sine_reg0   <= 36'sb110100111101110011100011110011001110;
        end
        15467: begin
            cosine_reg0 <= 36'sb11110000010101010011100111111100000;
            sine_reg0   <= 36'sb110100111110100010101111101100110100;
        end
        15468: begin
            cosine_reg0 <= 36'sb11110000010111011110000100010101110;
            sine_reg0   <= 36'sb110100111111010001111100000001100111;
        end
        15469: begin
            cosine_reg0 <= 36'sb11110000011001101000010111011110100;
            sine_reg0   <= 36'sb110101000000000001001000110001100101;
        end
        15470: begin
            cosine_reg0 <= 36'sb11110000011011110010100001010110000;
            sine_reg0   <= 36'sb110101000000110000010101111100101100;
        end
        15471: begin
            cosine_reg0 <= 36'sb11110000011101111100100001111100010;
            sine_reg0   <= 36'sb110101000001011111100011100010111001;
        end
        15472: begin
            cosine_reg0 <= 36'sb11110000100000000110011001010001001;
            sine_reg0   <= 36'sb110101000010001110110001100100001101;
        end
        15473: begin
            cosine_reg0 <= 36'sb11110000100010010000000111010100110;
            sine_reg0   <= 36'sb110101000010111110000000000000100011;
        end
        15474: begin
            cosine_reg0 <= 36'sb11110000100100011001101100000110110;
            sine_reg0   <= 36'sb110101000011101101001110110111111100;
        end
        15475: begin
            cosine_reg0 <= 36'sb11110000100110100011000111100111001;
            sine_reg0   <= 36'sb110101000100011100011110001010010100;
        end
        15476: begin
            cosine_reg0 <= 36'sb11110000101000101100011001110101111;
            sine_reg0   <= 36'sb110101000101001011101101110111101010;
        end
        15477: begin
            cosine_reg0 <= 36'sb11110000101010110101100010110011000;
            sine_reg0   <= 36'sb110101000101111010111101111111111101;
        end
        15478: begin
            cosine_reg0 <= 36'sb11110000101100111110100010011110001;
            sine_reg0   <= 36'sb110101000110101010001110100011001010;
        end
        15479: begin
            cosine_reg0 <= 36'sb11110000101111000111011000110111100;
            sine_reg0   <= 36'sb110101000111011001011111100001010000;
        end
        15480: begin
            cosine_reg0 <= 36'sb11110000110001010000000101111110110;
            sine_reg0   <= 36'sb110101001000001000110000111010001101;
        end
        15481: begin
            cosine_reg0 <= 36'sb11110000110011011000101001110100000;
            sine_reg0   <= 36'sb110101001000111000000010101101111110;
        end
        15482: begin
            cosine_reg0 <= 36'sb11110000110101100001000100010111001;
            sine_reg0   <= 36'sb110101001001100111010100111100100011;
        end
        15483: begin
            cosine_reg0 <= 36'sb11110000110111101001010101100111111;
            sine_reg0   <= 36'sb110101001010010110100111100101111001;
        end
        15484: begin
            cosine_reg0 <= 36'sb11110000111001110001011101100110011;
            sine_reg0   <= 36'sb110101001011000101111010101001111110;
        end
        15485: begin
            cosine_reg0 <= 36'sb11110000111011111001011100010010100;
            sine_reg0   <= 36'sb110101001011110101001110001000110010;
        end
        15486: begin
            cosine_reg0 <= 36'sb11110000111110000001010001101100001;
            sine_reg0   <= 36'sb110101001100100100100010000010010001;
        end
        15487: begin
            cosine_reg0 <= 36'sb11110001000000001000111101110011001;
            sine_reg0   <= 36'sb110101001101010011110110010110011010;
        end
        15488: begin
            cosine_reg0 <= 36'sb11110001000010010000100000100111101;
            sine_reg0   <= 36'sb110101001110000011001011000101001011;
        end
        15489: begin
            cosine_reg0 <= 36'sb11110001000100010111111010001001010;
            sine_reg0   <= 36'sb110101001110110010100000001110100011;
        end
        15490: begin
            cosine_reg0 <= 36'sb11110001000110011111001010011000001;
            sine_reg0   <= 36'sb110101001111100001110101110010011111;
        end
        15491: begin
            cosine_reg0 <= 36'sb11110001001000100110010001010100001;
            sine_reg0   <= 36'sb110101010000010001001011110000111110;
        end
        15492: begin
            cosine_reg0 <= 36'sb11110001001010101101001110111101001;
            sine_reg0   <= 36'sb110101010001000000100010001001111110;
        end
        15493: begin
            cosine_reg0 <= 36'sb11110001001100110100000011010011000;
            sine_reg0   <= 36'sb110101010001101111111000111101011101;
        end
        15494: begin
            cosine_reg0 <= 36'sb11110001001110111010101110010101110;
            sine_reg0   <= 36'sb110101010010011111010000001011011001;
        end
        15495: begin
            cosine_reg0 <= 36'sb11110001010001000001010000000101011;
            sine_reg0   <= 36'sb110101010011001110100111110011110001;
        end
        15496: begin
            cosine_reg0 <= 36'sb11110001010011000111101000100001101;
            sine_reg0   <= 36'sb110101010011111101111111110110100010;
        end
        15497: begin
            cosine_reg0 <= 36'sb11110001010101001101110111101010101;
            sine_reg0   <= 36'sb110101010100101101011000010011101011;
        end
        15498: begin
            cosine_reg0 <= 36'sb11110001010111010011111101100000000;
            sine_reg0   <= 36'sb110101010101011100110001001011001010;
        end
        15499: begin
            cosine_reg0 <= 36'sb11110001011001011001111010000001111;
            sine_reg0   <= 36'sb110101010110001100001010011100111101;
        end
        15500: begin
            cosine_reg0 <= 36'sb11110001011011011111101101010000001;
            sine_reg0   <= 36'sb110101010110111011100100001001000010;
        end
        15501: begin
            cosine_reg0 <= 36'sb11110001011101100101010111001010110;
            sine_reg0   <= 36'sb110101010111101010111110001111011000;
        end
        15502: begin
            cosine_reg0 <= 36'sb11110001011111101010110111110001100;
            sine_reg0   <= 36'sb110101011000011010011000101111111101;
        end
        15503: begin
            cosine_reg0 <= 36'sb11110001100001110000001111000100011;
            sine_reg0   <= 36'sb110101011001001001110011101010101110;
        end
        15504: begin
            cosine_reg0 <= 36'sb11110001100011110101011101000011011;
            sine_reg0   <= 36'sb110101011001111001001110111111101010;
        end
        15505: begin
            cosine_reg0 <= 36'sb11110001100101111010100001101110011;
            sine_reg0   <= 36'sb110101011010101000101010101110110000;
        end
        15506: begin
            cosine_reg0 <= 36'sb11110001100111111111011101000101010;
            sine_reg0   <= 36'sb110101011011011000000110110111111101;
        end
        15507: begin
            cosine_reg0 <= 36'sb11110001101010000100001111000111111;
            sine_reg0   <= 36'sb110101011100000111100011011011001111;
        end
        15508: begin
            cosine_reg0 <= 36'sb11110001101100001000110111110110010;
            sine_reg0   <= 36'sb110101011100110111000000011000100101;
        end
        15509: begin
            cosine_reg0 <= 36'sb11110001101110001101010111010000010;
            sine_reg0   <= 36'sb110101011101100110011101101111111101;
        end
        15510: begin
            cosine_reg0 <= 36'sb11110001110000010001101101010101111;
            sine_reg0   <= 36'sb110101011110010101111011100001010101;
        end
        15511: begin
            cosine_reg0 <= 36'sb11110001110010010101111010000111000;
            sine_reg0   <= 36'sb110101011111000101011001101100101011;
        end
        15512: begin
            cosine_reg0 <= 36'sb11110001110100011001111101100011101;
            sine_reg0   <= 36'sb110101011111110100111000010001111101;
        end
        15513: begin
            cosine_reg0 <= 36'sb11110001110110011101110111101011011;
            sine_reg0   <= 36'sb110101100000100100010111010001001010;
        end
        15514: begin
            cosine_reg0 <= 36'sb11110001111000100001101000011110100;
            sine_reg0   <= 36'sb110101100001010011110110101010010000;
        end
        15515: begin
            cosine_reg0 <= 36'sb11110001111010100101001111111100111;
            sine_reg0   <= 36'sb110101100010000011010110011101001100;
        end
        15516: begin
            cosine_reg0 <= 36'sb11110001111100101000101110000110010;
            sine_reg0   <= 36'sb110101100010110010110110101001111110;
        end
        15517: begin
            cosine_reg0 <= 36'sb11110001111110101100000010111010101;
            sine_reg0   <= 36'sb110101100011100010010111010000100010;
        end
        15518: begin
            cosine_reg0 <= 36'sb11110010000000101111001110011010000;
            sine_reg0   <= 36'sb110101100100010001111000010000111000;
        end
        15519: begin
            cosine_reg0 <= 36'sb11110010000010110010010000100100010;
            sine_reg0   <= 36'sb110101100101000001011001101010111110;
        end
        15520: begin
            cosine_reg0 <= 36'sb11110010000100110101001001011001010;
            sine_reg0   <= 36'sb110101100101110000111011011110110001;
        end
        15521: begin
            cosine_reg0 <= 36'sb11110010000110110111111000111001000;
            sine_reg0   <= 36'sb110101100110100000011101101100010000;
        end
        15522: begin
            cosine_reg0 <= 36'sb11110010001000111010011111000011010;
            sine_reg0   <= 36'sb110101100111010000000000010011011010;
        end
        15523: begin
            cosine_reg0 <= 36'sb11110010001010111100111011111000001;
            sine_reg0   <= 36'sb110101100111111111100011010100001011;
        end
        15524: begin
            cosine_reg0 <= 36'sb11110010001100111111001111010111100;
            sine_reg0   <= 36'sb110101101000101111000110101110100011;
        end
        15525: begin
            cosine_reg0 <= 36'sb11110010001111000001011001100001010;
            sine_reg0   <= 36'sb110101101001011110101010100010011111;
        end
        15526: begin
            cosine_reg0 <= 36'sb11110010010001000011011010010101010;
            sine_reg0   <= 36'sb110101101010001110001110101111111110;
        end
        15527: begin
            cosine_reg0 <= 36'sb11110010010011000101010001110011100;
            sine_reg0   <= 36'sb110101101010111101110011010110111110;
        end
        15528: begin
            cosine_reg0 <= 36'sb11110010010101000110111111111100000;
            sine_reg0   <= 36'sb110101101011101101011000010111011101;
        end
        15529: begin
            cosine_reg0 <= 36'sb11110010010111001000100100101110011;
            sine_reg0   <= 36'sb110101101100011100111101110001011001;
        end
        15530: begin
            cosine_reg0 <= 36'sb11110010011001001010000000001010111;
            sine_reg0   <= 36'sb110101101101001100100011100100110001;
        end
        15531: begin
            cosine_reg0 <= 36'sb11110010011011001011010010010001011;
            sine_reg0   <= 36'sb110101101101111100001001110001100010;
        end
        15532: begin
            cosine_reg0 <= 36'sb11110010011101001100011011000001101;
            sine_reg0   <= 36'sb110101101110101011110000010111101010;
        end
        15533: begin
            cosine_reg0 <= 36'sb11110010011111001101011010011011101;
            sine_reg0   <= 36'sb110101101111011011010111010111001001;
        end
        15534: begin
            cosine_reg0 <= 36'sb11110010100001001110010000011111010;
            sine_reg0   <= 36'sb110101110000001010111110101111111011;
        end
        15535: begin
            cosine_reg0 <= 36'sb11110010100011001110111101001100101;
            sine_reg0   <= 36'sb110101110000111010100110100010000000;
        end
        15536: begin
            cosine_reg0 <= 36'sb11110010100101001111100000100011100;
            sine_reg0   <= 36'sb110101110001101010001110101101010101;
        end
        15537: begin
            cosine_reg0 <= 36'sb11110010100111001111111010100011110;
            sine_reg0   <= 36'sb110101110010011001110111010001111001;
        end
        15538: begin
            cosine_reg0 <= 36'sb11110010101001010000001011001101011;
            sine_reg0   <= 36'sb110101110011001001100000001111101001;
        end
        15539: begin
            cosine_reg0 <= 36'sb11110010101011010000010010100000011;
            sine_reg0   <= 36'sb110101110011111001001001100110100101;
        end
        15540: begin
            cosine_reg0 <= 36'sb11110010101101010000010000011100101;
            sine_reg0   <= 36'sb110101110100101000110011010110101001;
        end
        15541: begin
            cosine_reg0 <= 36'sb11110010101111010000000101000001111;
            sine_reg0   <= 36'sb110101110101011000011101011111110100;
        end
        15542: begin
            cosine_reg0 <= 36'sb11110010110001001111110000010000011;
            sine_reg0   <= 36'sb110101110110001000001000000010000101;
        end
        15543: begin
            cosine_reg0 <= 36'sb11110010110011001111010010000111110;
            sine_reg0   <= 36'sb110101110110110111110010111101011001;
        end
        15544: begin
            cosine_reg0 <= 36'sb11110010110101001110101010101000000;
            sine_reg0   <= 36'sb110101110111100111011110010001101111;
        end
        15545: begin
            cosine_reg0 <= 36'sb11110010110111001101111001110001001;
            sine_reg0   <= 36'sb110101111000010111001001111111000101;
        end
        15546: begin
            cosine_reg0 <= 36'sb11110010111001001100111111100011001;
            sine_reg0   <= 36'sb110101111001000110110110000101011001;
        end
        15547: begin
            cosine_reg0 <= 36'sb11110010111011001011111011111101101;
            sine_reg0   <= 36'sb110101111001110110100010100100101000;
        end
        15548: begin
            cosine_reg0 <= 36'sb11110010111101001010101111000000111;
            sine_reg0   <= 36'sb110101111010100110001111011100110011;
        end
        15549: begin
            cosine_reg0 <= 36'sb11110010111111001001011000101100101;
            sine_reg0   <= 36'sb110101111011010101111100101101110101;
        end
        15550: begin
            cosine_reg0 <= 36'sb11110011000001000111111001000000110;
            sine_reg0   <= 36'sb110101111100000101101010010111101110;
        end
        15551: begin
            cosine_reg0 <= 36'sb11110011000011000110001111111101010;
            sine_reg0   <= 36'sb110101111100110101011000011010011100;
        end
        15552: begin
            cosine_reg0 <= 36'sb11110011000101000100011101100010001;
            sine_reg0   <= 36'sb110101111101100101000110110101111101;
        end
        15553: begin
            cosine_reg0 <= 36'sb11110011000111000010100001101111010;
            sine_reg0   <= 36'sb110101111110010100110101101010001111;
        end
        15554: begin
            cosine_reg0 <= 36'sb11110011001001000000011100100100100;
            sine_reg0   <= 36'sb110101111111000100100100110111010001;
        end
        15555: begin
            cosine_reg0 <= 36'sb11110011001010111110001110000001110;
            sine_reg0   <= 36'sb110101111111110100010100011101000000;
        end
        15556: begin
            cosine_reg0 <= 36'sb11110011001100111011110110000111001;
            sine_reg0   <= 36'sb110110000000100100000100011011011010;
        end
        15557: begin
            cosine_reg0 <= 36'sb11110011001110111001010100110100011;
            sine_reg0   <= 36'sb110110000001010011110100110010011110;
        end
        15558: begin
            cosine_reg0 <= 36'sb11110011010000110110101010001001011;
            sine_reg0   <= 36'sb110110000010000011100101100010001010;
        end
        15559: begin
            cosine_reg0 <= 36'sb11110011010010110011110110000110010;
            sine_reg0   <= 36'sb110110000010110011010110101010011100;
        end
        15560: begin
            cosine_reg0 <= 36'sb11110011010100110000111000101010110;
            sine_reg0   <= 36'sb110110000011100011001000001011010010;
        end
        15561: begin
            cosine_reg0 <= 36'sb11110011010110101101110001110111000;
            sine_reg0   <= 36'sb110110000100010010111010000100101011;
        end
        15562: begin
            cosine_reg0 <= 36'sb11110011011000101010100001101010101;
            sine_reg0   <= 36'sb110110000101000010101100010110100100;
        end
        15563: begin
            cosine_reg0 <= 36'sb11110011011010100111001000000101111;
            sine_reg0   <= 36'sb110110000101110010011111000000111100;
        end
        15564: begin
            cosine_reg0 <= 36'sb11110011011100100011100101001000100;
            sine_reg0   <= 36'sb110110000110100010010010000011110001;
        end
        15565: begin
            cosine_reg0 <= 36'sb11110011011110011111111000110010011;
            sine_reg0   <= 36'sb110110000111010010000101011111000001;
        end
        15566: begin
            cosine_reg0 <= 36'sb11110011100000011100000011000011100;
            sine_reg0   <= 36'sb110110001000000001111001010010101010;
        end
        15567: begin
            cosine_reg0 <= 36'sb11110011100010011000000011111011110;
            sine_reg0   <= 36'sb110110001000110001101101011110101010;
        end
        15568: begin
            cosine_reg0 <= 36'sb11110011100100010011111011011011010;
            sine_reg0   <= 36'sb110110001001100001100010000011000000;
        end
        15569: begin
            cosine_reg0 <= 36'sb11110011100110001111101001100001101;
            sine_reg0   <= 36'sb110110001010010001010110111111101001;
        end
        15570: begin
            cosine_reg0 <= 36'sb11110011101000001011001110001111000;
            sine_reg0   <= 36'sb110110001011000001001100010100100100;
        end
        15571: begin
            cosine_reg0 <= 36'sb11110011101010000110101001100011010;
            sine_reg0   <= 36'sb110110001011110001000010000001110000;
        end
        15572: begin
            cosine_reg0 <= 36'sb11110011101100000001111011011110011;
            sine_reg0   <= 36'sb110110001100100000111000000111001001;
        end
        15573: begin
            cosine_reg0 <= 36'sb11110011101101111101000100000000001;
            sine_reg0   <= 36'sb110110001101010000101110100100101110;
        end
        15574: begin
            cosine_reg0 <= 36'sb11110011101111111000000011001000100;
            sine_reg0   <= 36'sb110110001110000000100101011010011110;
        end
        15575: begin
            cosine_reg0 <= 36'sb11110011110001110010111000110111100;
            sine_reg0   <= 36'sb110110001110110000011100101000010111;
        end
        15576: begin
            cosine_reg0 <= 36'sb11110011110011101101100101001101000;
            sine_reg0   <= 36'sb110110001111100000010100001110010110;
        end
        15577: begin
            cosine_reg0 <= 36'sb11110011110101101000001000001001000;
            sine_reg0   <= 36'sb110110010000010000001100001100011010;
        end
        15578: begin
            cosine_reg0 <= 36'sb11110011110111100010100001101011010;
            sine_reg0   <= 36'sb110110010001000000000100100010100001;
        end
        15579: begin
            cosine_reg0 <= 36'sb11110011111001011100110001110011111;
            sine_reg0   <= 36'sb110110010001101111111101010000101001;
        end
        15580: begin
            cosine_reg0 <= 36'sb11110011111011010110111000100010101;
            sine_reg0   <= 36'sb110110010010011111110110010110110001;
        end
        15581: begin
            cosine_reg0 <= 36'sb11110011111101010000110101110111100;
            sine_reg0   <= 36'sb110110010011001111101111110100110110;
        end
        15582: begin
            cosine_reg0 <= 36'sb11110011111111001010101001110010100;
            sine_reg0   <= 36'sb110110010011111111101001101010110111;
        end
        15583: begin
            cosine_reg0 <= 36'sb11110100000001000100010100010011011;
            sine_reg0   <= 36'sb110110010100101111100011111000110010;
        end
        15584: begin
            cosine_reg0 <= 36'sb11110100000010111101110101011010010;
            sine_reg0   <= 36'sb110110010101011111011110011110100100;
        end
        15585: begin
            cosine_reg0 <= 36'sb11110100000100110111001101000111000;
            sine_reg0   <= 36'sb110110010110001111011001011100001101;
        end
        15586: begin
            cosine_reg0 <= 36'sb11110100000110110000011011011001100;
            sine_reg0   <= 36'sb110110010110111111010100110001101010;
        end
        15587: begin
            cosine_reg0 <= 36'sb11110100001000101001100000010001101;
            sine_reg0   <= 36'sb110110010111101111010000011110111001;
        end
        15588: begin
            cosine_reg0 <= 36'sb11110100001010100010011011101111011;
            sine_reg0   <= 36'sb110110011000011111001100100011111001;
        end
        15589: begin
            cosine_reg0 <= 36'sb11110100001100011011001101110010110;
            sine_reg0   <= 36'sb110110011001001111001001000000101000;
        end
        15590: begin
            cosine_reg0 <= 36'sb11110100001110010011110110011011100;
            sine_reg0   <= 36'sb110110011001111111000101110101000011;
        end
        15591: begin
            cosine_reg0 <= 36'sb11110100010000001100010101101001110;
            sine_reg0   <= 36'sb110110011010101111000011000001001010;
        end
        15592: begin
            cosine_reg0 <= 36'sb11110100010010000100101011011101010;
            sine_reg0   <= 36'sb110110011011011111000000100100111001;
        end
        15593: begin
            cosine_reg0 <= 36'sb11110100010011111100110111110110001;
            sine_reg0   <= 36'sb110110011100001110111110100000010000;
        end
        15594: begin
            cosine_reg0 <= 36'sb11110100010101110100111010110100001;
            sine_reg0   <= 36'sb110110011100111110111100110011001101;
        end
        15595: begin
            cosine_reg0 <= 36'sb11110100010111101100110100010111001;
            sine_reg0   <= 36'sb110110011101101110111011011101101101;
        end
        15596: begin
            cosine_reg0 <= 36'sb11110100011001100100100100011111010;
            sine_reg0   <= 36'sb110110011110011110111010011111101111;
        end
        15597: begin
            cosine_reg0 <= 36'sb11110100011011011100001011001100011;
            sine_reg0   <= 36'sb110110011111001110111001111001010000;
        end
        15598: begin
            cosine_reg0 <= 36'sb11110100011101010011101000011110011;
            sine_reg0   <= 36'sb110110011111111110111001101010010000;
        end
        15599: begin
            cosine_reg0 <= 36'sb11110100011111001010111100010101010;
            sine_reg0   <= 36'sb110110100000101110111001110010101100;
        end
        15600: begin
            cosine_reg0 <= 36'sb11110100100001000010000110110000111;
            sine_reg0   <= 36'sb110110100001011110111010010010100011;
        end
        15601: begin
            cosine_reg0 <= 36'sb11110100100010111001000111110001001;
            sine_reg0   <= 36'sb110110100010001110111011001001110010;
        end
        15602: begin
            cosine_reg0 <= 36'sb11110100100100101111111111010110000;
            sine_reg0   <= 36'sb110110100010111110111100011000010111;
        end
        15603: begin
            cosine_reg0 <= 36'sb11110100100110100110101101011111011;
            sine_reg0   <= 36'sb110110100011101110111101111110010010;
        end
        15604: begin
            cosine_reg0 <= 36'sb11110100101000011101010010001101010;
            sine_reg0   <= 36'sb110110100100011110111111111011011111;
        end
        15605: begin
            cosine_reg0 <= 36'sb11110100101010010011101101011111100;
            sine_reg0   <= 36'sb110110100101001111000010001111111110;
        end
        15606: begin
            cosine_reg0 <= 36'sb11110100101100001001111111010110001;
            sine_reg0   <= 36'sb110110100101111111000100111011101100;
        end
        15607: begin
            cosine_reg0 <= 36'sb11110100101110000000000111110000111;
            sine_reg0   <= 36'sb110110100110101111000111111110100111;
        end
        15608: begin
            cosine_reg0 <= 36'sb11110100101111110110000110101111111;
            sine_reg0   <= 36'sb110110100111011111001011011000101110;
        end
        15609: begin
            cosine_reg0 <= 36'sb11110100110001101011111100010011000;
            sine_reg0   <= 36'sb110110101000001111001111001001111110;
        end
        15610: begin
            cosine_reg0 <= 36'sb11110100110011100001101000011010010;
            sine_reg0   <= 36'sb110110101000111111010011010010010110;
        end
        15611: begin
            cosine_reg0 <= 36'sb11110100110101010111001011000101011;
            sine_reg0   <= 36'sb110110101001101111010111110001110101;
        end
        15612: begin
            cosine_reg0 <= 36'sb11110100110111001100100100010100011;
            sine_reg0   <= 36'sb110110101010011111011100101000010111;
        end
        15613: begin
            cosine_reg0 <= 36'sb11110100111001000001110100000111010;
            sine_reg0   <= 36'sb110110101011001111100001110101111100;
        end
        15614: begin
            cosine_reg0 <= 36'sb11110100111010110110111010011101111;
            sine_reg0   <= 36'sb110110101011111111100111011010100001;
        end
        15615: begin
            cosine_reg0 <= 36'sb11110100111100101011110111011000001;
            sine_reg0   <= 36'sb110110101100101111101101010110000101;
        end
        15616: begin
            cosine_reg0 <= 36'sb11110100111110100000101010110110001;
            sine_reg0   <= 36'sb110110101101011111110011101000100110;
        end
        15617: begin
            cosine_reg0 <= 36'sb11110101000000010101010100110111100;
            sine_reg0   <= 36'sb110110101110001111111010010010000001;
        end
        15618: begin
            cosine_reg0 <= 36'sb11110101000010001001110101011100100;
            sine_reg0   <= 36'sb110110101111000000000001010010010101;
        end
        15619: begin
            cosine_reg0 <= 36'sb11110101000011111110001100100100110;
            sine_reg0   <= 36'sb110110101111110000001000101001100001;
        end
        15620: begin
            cosine_reg0 <= 36'sb11110101000101110010011010010000100;
            sine_reg0   <= 36'sb110110110000100000010000010111100010;
        end
        15621: begin
            cosine_reg0 <= 36'sb11110101000111100110011110011111011;
            sine_reg0   <= 36'sb110110110001010000011000011100010110;
        end
        15622: begin
            cosine_reg0 <= 36'sb11110101001001011010011001010001100;
            sine_reg0   <= 36'sb110110110010000000100000110111111100;
        end
        15623: begin
            cosine_reg0 <= 36'sb11110101001011001110001010100110110;
            sine_reg0   <= 36'sb110110110010110000101001101010010010;
        end
        15624: begin
            cosine_reg0 <= 36'sb11110101001101000001110010011111001;
            sine_reg0   <= 36'sb110110110011100000110010110011010110;
        end
        15625: begin
            cosine_reg0 <= 36'sb11110101001110110101010000111010011;
            sine_reg0   <= 36'sb110110110100010000111100010011000101;
        end
        15626: begin
            cosine_reg0 <= 36'sb11110101010000101000100101111000101;
            sine_reg0   <= 36'sb110110110101000001000110001001011111;
        end
        15627: begin
            cosine_reg0 <= 36'sb11110101010010011011110001011001101;
            sine_reg0   <= 36'sb110110110101110001010000010110100001;
        end
        15628: begin
            cosine_reg0 <= 36'sb11110101010100001110110011011101100;
            sine_reg0   <= 36'sb110110110110100001011010111010001010;
        end
        15629: begin
            cosine_reg0 <= 36'sb11110101010110000001101100000100000;
            sine_reg0   <= 36'sb110110110111010001100101110100010111;
        end
        15630: begin
            cosine_reg0 <= 36'sb11110101010111110100011011001101001;
            sine_reg0   <= 36'sb110110111000000001110001000101000111;
        end
        15631: begin
            cosine_reg0 <= 36'sb11110101011001100111000000111000111;
            sine_reg0   <= 36'sb110110111000110001111100101100011000;
        end
        15632: begin
            cosine_reg0 <= 36'sb11110101011011011001011101000111001;
            sine_reg0   <= 36'sb110110111001100010001000101010001000;
        end
        15633: begin
            cosine_reg0 <= 36'sb11110101011101001011101111110111110;
            sine_reg0   <= 36'sb110110111010010010010100111110010101;
        end
        15634: begin
            cosine_reg0 <= 36'sb11110101011110111101111001001010111;
            sine_reg0   <= 36'sb110110111011000010100001101000111101;
        end
        15635: begin
            cosine_reg0 <= 36'sb11110101100000101111111001000000001;
            sine_reg0   <= 36'sb110110111011110010101110101001111111;
        end
        15636: begin
            cosine_reg0 <= 36'sb11110101100010100001101111010111101;
            sine_reg0   <= 36'sb110110111100100010111100000001011001;
        end
        15637: begin
            cosine_reg0 <= 36'sb11110101100100010011011100010001011;
            sine_reg0   <= 36'sb110110111101010011001001101111001000;
        end
        15638: begin
            cosine_reg0 <= 36'sb11110101100110000100111111101101001;
            sine_reg0   <= 36'sb110110111110000011010111110011001011;
        end
        15639: begin
            cosine_reg0 <= 36'sb11110101100111110110011001101011000;
            sine_reg0   <= 36'sb110110111110110011100110001101100000;
        end
        15640: begin
            cosine_reg0 <= 36'sb11110101101001100111101010001010110;
            sine_reg0   <= 36'sb110110111111100011110100111110000101;
        end
        15641: begin
            cosine_reg0 <= 36'sb11110101101011011000110001001100011;
            sine_reg0   <= 36'sb110111000000010100000100000100111001;
        end
        15642: begin
            cosine_reg0 <= 36'sb11110101101101001001101110101111111;
            sine_reg0   <= 36'sb110111000001000100010011100001111001;
        end
        15643: begin
            cosine_reg0 <= 36'sb11110101101110111010100010110101000;
            sine_reg0   <= 36'sb110111000001110100100011010101000100;
        end
        15644: begin
            cosine_reg0 <= 36'sb11110101110000101011001101011011111;
            sine_reg0   <= 36'sb110111000010100100110011011110010111;
        end
        15645: begin
            cosine_reg0 <= 36'sb11110101110010011011101110100100011;
            sine_reg0   <= 36'sb110111000011010101000011111101110001;
        end
        15646: begin
            cosine_reg0 <= 36'sb11110101110100001100000110001110011;
            sine_reg0   <= 36'sb110111000100000101010100110011010001;
        end
        15647: begin
            cosine_reg0 <= 36'sb11110101110101111100010100011010000;
            sine_reg0   <= 36'sb110111000100110101100101111110110011;
        end
        15648: begin
            cosine_reg0 <= 36'sb11110101110111101100011001000110111;
            sine_reg0   <= 36'sb110111000101100101110111100000010111;
        end
        15649: begin
            cosine_reg0 <= 36'sb11110101111001011100010100010101001;
            sine_reg0   <= 36'sb110111000110010110001001010111111010;
        end
        15650: begin
            cosine_reg0 <= 36'sb11110101111011001100000110000100101;
            sine_reg0   <= 36'sb110111000111000110011011100101011010;
        end
        15651: begin
            cosine_reg0 <= 36'sb11110101111100111011101110010101011;
            sine_reg0   <= 36'sb110111000111110110101110001000110111;
        end
        15652: begin
            cosine_reg0 <= 36'sb11110101111110101011001101000111010;
            sine_reg0   <= 36'sb110111001000100111000001000010001101;
        end
        15653: begin
            cosine_reg0 <= 36'sb11110110000000011010100010011010001;
            sine_reg0   <= 36'sb110111001001010111010100010001011011;
        end
        15654: begin
            cosine_reg0 <= 36'sb11110110000010001001101110001110001;
            sine_reg0   <= 36'sb110111001010000111100111110110100000;
        end
        15655: begin
            cosine_reg0 <= 36'sb11110110000011111000110000100011000;
            sine_reg0   <= 36'sb110111001010110111111011110001011000;
        end
        15656: begin
            cosine_reg0 <= 36'sb11110110000101100111101001011000110;
            sine_reg0   <= 36'sb110111001011101000010000000010000011;
        end
        15657: begin
            cosine_reg0 <= 36'sb11110110000111010110011000101111010;
            sine_reg0   <= 36'sb110111001100011000100100101000011111;
        end
        15658: begin
            cosine_reg0 <= 36'sb11110110001001000100111110100110100;
            sine_reg0   <= 36'sb110111001101001000111001100100101001;
        end
        15659: begin
            cosine_reg0 <= 36'sb11110110001010110011011010111110100;
            sine_reg0   <= 36'sb110111001101111001001110110110100000;
        end
        15660: begin
            cosine_reg0 <= 36'sb11110110001100100001101101110111001;
            sine_reg0   <= 36'sb110111001110101001100100011110000010;
        end
        15661: begin
            cosine_reg0 <= 36'sb11110110001110001111110111010000001;
            sine_reg0   <= 36'sb110111001111011001111010011011001101;
        end
        15662: begin
            cosine_reg0 <= 36'sb11110110001111111101110111001001110;
            sine_reg0   <= 36'sb110111010000001010010000101101111111;
        end
        15663: begin
            cosine_reg0 <= 36'sb11110110010001101011101101100011110;
            sine_reg0   <= 36'sb110111010000111010100111010110010110;
        end
        15664: begin
            cosine_reg0 <= 36'sb11110110010011011001011010011110000;
            sine_reg0   <= 36'sb110111010001101010111110010100010001;
        end
        15665: begin
            cosine_reg0 <= 36'sb11110110010101000110111101111000101;
            sine_reg0   <= 36'sb110111010010011011010101100111101110;
        end
        15666: begin
            cosine_reg0 <= 36'sb11110110010110110100010111110011011;
            sine_reg0   <= 36'sb110111010011001011101101010000101011;
        end
        15667: begin
            cosine_reg0 <= 36'sb11110110011000100001101000001110010;
            sine_reg0   <= 36'sb110111010011111100000101001111000101;
        end
        15668: begin
            cosine_reg0 <= 36'sb11110110011010001110101111001001010;
            sine_reg0   <= 36'sb110111010100101100011101100010111011;
        end
        15669: begin
            cosine_reg0 <= 36'sb11110110011011111011101100100100010;
            sine_reg0   <= 36'sb110111010101011100110110001100001100;
        end
        15670: begin
            cosine_reg0 <= 36'sb11110110011101101000100000011111010;
            sine_reg0   <= 36'sb110111010110001101001111001010110100;
        end
        15671: begin
            cosine_reg0 <= 36'sb11110110011111010101001010111010000;
            sine_reg0   <= 36'sb110111010110111101101000011110110100;
        end
        15672: begin
            cosine_reg0 <= 36'sb11110110100001000001101011110100101;
            sine_reg0   <= 36'sb110111010111101110000010001000000111;
        end
        15673: begin
            cosine_reg0 <= 36'sb11110110100010101110000011001111000;
            sine_reg0   <= 36'sb110111011000011110011100000110101110;
        end
        15674: begin
            cosine_reg0 <= 36'sb11110110100100011010010001001001001;
            sine_reg0   <= 36'sb110111011001001110110110011010100101;
        end
        15675: begin
            cosine_reg0 <= 36'sb11110110100110000110010101100010110;
            sine_reg0   <= 36'sb110111011001111111010001000011101100;
        end
        15676: begin
            cosine_reg0 <= 36'sb11110110100111110010010000011100000;
            sine_reg0   <= 36'sb110111011010101111101100000001111111;
        end
        15677: begin
            cosine_reg0 <= 36'sb11110110101001011110000001110100110;
            sine_reg0   <= 36'sb110111011011100000000111010101011101;
        end
        15678: begin
            cosine_reg0 <= 36'sb11110110101011001001101001101100111;
            sine_reg0   <= 36'sb110111011100010000100010111110000101;
        end
        15679: begin
            cosine_reg0 <= 36'sb11110110101100110101001000000100011;
            sine_reg0   <= 36'sb110111011101000000111110111011110101;
        end
        15680: begin
            cosine_reg0 <= 36'sb11110110101110100000011100111011001;
            sine_reg0   <= 36'sb110111011101110001011011001110101010;
        end
        15681: begin
            cosine_reg0 <= 36'sb11110110110000001011101000010001001;
            sine_reg0   <= 36'sb110111011110100001110111110110100011;
        end
        15682: begin
            cosine_reg0 <= 36'sb11110110110001110110101010000110011;
            sine_reg0   <= 36'sb110111011111010010010100110011011110;
        end
        15683: begin
            cosine_reg0 <= 36'sb11110110110011100001100010011010101;
            sine_reg0   <= 36'sb110111100000000010110010000101011000;
        end
        15684: begin
            cosine_reg0 <= 36'sb11110110110101001100010001001101111;
            sine_reg0   <= 36'sb110111100000110011001111101100010001;
        end
        15685: begin
            cosine_reg0 <= 36'sb11110110110110110110110110100000001;
            sine_reg0   <= 36'sb110111100001100011101101101000000111;
        end
        15686: begin
            cosine_reg0 <= 36'sb11110110111000100001010010010001011;
            sine_reg0   <= 36'sb110111100010010100001011111000110110;
        end
        15687: begin
            cosine_reg0 <= 36'sb11110110111010001011100100100001011;
            sine_reg0   <= 36'sb110111100011000100101010011110011110;
        end
        15688: begin
            cosine_reg0 <= 36'sb11110110111011110101101101010000001;
            sine_reg0   <= 36'sb110111100011110101001001011000111101;
        end
        15689: begin
            cosine_reg0 <= 36'sb11110110111101011111101100011101101;
            sine_reg0   <= 36'sb110111100100100101101000101000010001;
        end
        15690: begin
            cosine_reg0 <= 36'sb11110110111111001001100010001001110;
            sine_reg0   <= 36'sb110111100101010110001000001100011000;
        end
        15691: begin
            cosine_reg0 <= 36'sb11110111000000110011001110010100100;
            sine_reg0   <= 36'sb110111100110000110101000000101001111;
        end
        15692: begin
            cosine_reg0 <= 36'sb11110111000010011100110000111101110;
            sine_reg0   <= 36'sb110111100110110111001000010010110110;
        end
        15693: begin
            cosine_reg0 <= 36'sb11110111000100000110001010000101100;
            sine_reg0   <= 36'sb110111100111100111101000110101001011;
        end
        15694: begin
            cosine_reg0 <= 36'sb11110111000101101111011001101011101;
            sine_reg0   <= 36'sb110111101000011000001001101100001010;
        end
        15695: begin
            cosine_reg0 <= 36'sb11110111000111011000011111110000000;
            sine_reg0   <= 36'sb110111101001001000101010110111110100;
        end
        15696: begin
            cosine_reg0 <= 36'sb11110111001001000001011100010010110;
            sine_reg0   <= 36'sb110111101001111001001100011000000101;
        end
        15697: begin
            cosine_reg0 <= 36'sb11110111001010101010001111010011101;
            sine_reg0   <= 36'sb110111101010101001101110001100111100;
        end
        15698: begin
            cosine_reg0 <= 36'sb11110111001100010010111000110010101;
            sine_reg0   <= 36'sb110111101011011010010000010110010111;
        end
        15699: begin
            cosine_reg0 <= 36'sb11110111001101111011011000101111110;
            sine_reg0   <= 36'sb110111101100001010110010110100010100;
        end
        15700: begin
            cosine_reg0 <= 36'sb11110111001111100011101111001010111;
            sine_reg0   <= 36'sb110111101100111011010101100110110001;
        end
        15701: begin
            cosine_reg0 <= 36'sb11110111010001001011111100000100000;
            sine_reg0   <= 36'sb110111101101101011111000101101101100;
        end
        15702: begin
            cosine_reg0 <= 36'sb11110111010010110011111111011011000;
            sine_reg0   <= 36'sb110111101110011100011100001001000101;
        end
        15703: begin
            cosine_reg0 <= 36'sb11110111010100011011111001001111111;
            sine_reg0   <= 36'sb110111101111001100111111111000110111;
        end
        15704: begin
            cosine_reg0 <= 36'sb11110111010110000011101001100010011;
            sine_reg0   <= 36'sb110111101111111101100011111101000011;
        end
        15705: begin
            cosine_reg0 <= 36'sb11110111010111101011010000010010101;
            sine_reg0   <= 36'sb110111110000101110001000010101100101;
        end
        15706: begin
            cosine_reg0 <= 36'sb11110111011001010010101101100000101;
            sine_reg0   <= 36'sb110111110001011110101101000010011101;
        end
        15707: begin
            cosine_reg0 <= 36'sb11110111011010111010000001001100001;
            sine_reg0   <= 36'sb110111110010001111010010000011100111;
        end
        15708: begin
            cosine_reg0 <= 36'sb11110111011100100001001011010101001;
            sine_reg0   <= 36'sb110111110010111111110111011001000011;
        end
        15709: begin
            cosine_reg0 <= 36'sb11110111011110001000001011111011100;
            sine_reg0   <= 36'sb110111110011110000011101000010101110;
        end
        15710: begin
            cosine_reg0 <= 36'sb11110111011111101111000010111111011;
            sine_reg0   <= 36'sb110111110100100001000011000000100111;
        end
        15711: begin
            cosine_reg0 <= 36'sb11110111100001010101110000100000101;
            sine_reg0   <= 36'sb110111110101010001101001010010101011;
        end
        15712: begin
            cosine_reg0 <= 36'sb11110111100010111100010100011111000;
            sine_reg0   <= 36'sb110111110110000010001111111000111001;
        end
        15713: begin
            cosine_reg0 <= 36'sb11110111100100100010101110111010101;
            sine_reg0   <= 36'sb110111110110110010110110110011001111;
        end
        15714: begin
            cosine_reg0 <= 36'sb11110111100110001000111111110011100;
            sine_reg0   <= 36'sb110111110111100011011110000001101011;
        end
        15715: begin
            cosine_reg0 <= 36'sb11110111100111101111000111001001011;
            sine_reg0   <= 36'sb110111111000010100000101100100001011;
        end
        15716: begin
            cosine_reg0 <= 36'sb11110111101001010101000100111100010;
            sine_reg0   <= 36'sb110111111001000100101101011010101110;
        end
        15717: begin
            cosine_reg0 <= 36'sb11110111101010111010111001001100001;
            sine_reg0   <= 36'sb110111111001110101010101100101010001;
        end
        15718: begin
            cosine_reg0 <= 36'sb11110111101100100000100011111000111;
            sine_reg0   <= 36'sb110111111010100101111110000011110010;
        end
        15719: begin
            cosine_reg0 <= 36'sb11110111101110000110000101000010011;
            sine_reg0   <= 36'sb110111111011010110100110110110010000;
        end
        15720: begin
            cosine_reg0 <= 36'sb11110111101111101011011100101000110;
            sine_reg0   <= 36'sb110111111100000111001111111100101001;
        end
        15721: begin
            cosine_reg0 <= 36'sb11110111110001010000101010101011111;
            sine_reg0   <= 36'sb110111111100110111111001010110111011;
        end
        15722: begin
            cosine_reg0 <= 36'sb11110111110010110101101111001011101;
            sine_reg0   <= 36'sb110111111101101000100011000101000011;
        end
        15723: begin
            cosine_reg0 <= 36'sb11110111110100011010101010000111111;
            sine_reg0   <= 36'sb110111111110011001001101000111000001;
        end
        15724: begin
            cosine_reg0 <= 36'sb11110111110101111111011011100000110;
            sine_reg0   <= 36'sb110111111111001001110111011100110010;
        end
        15725: begin
            cosine_reg0 <= 36'sb11110111110111100100000011010110001;
            sine_reg0   <= 36'sb110111111111111010100010000110010101;
        end
        15726: begin
            cosine_reg0 <= 36'sb11110111111001001000100001100111110;
            sine_reg0   <= 36'sb111000000000101011001101000011100111;
        end
        15727: begin
            cosine_reg0 <= 36'sb11110111111010101100110110010101111;
            sine_reg0   <= 36'sb111000000001011011111000010100100111;
        end
        15728: begin
            cosine_reg0 <= 36'sb11110111111100010001000001100000010;
            sine_reg0   <= 36'sb111000000010001100100011111001010010;
        end
        15729: begin
            cosine_reg0 <= 36'sb11110111111101110101000011000110111;
            sine_reg0   <= 36'sb111000000010111101001111110001101000;
        end
        15730: begin
            cosine_reg0 <= 36'sb11110111111111011000111011001001101;
            sine_reg0   <= 36'sb111000000011101101111011111101100101;
        end
        15731: begin
            cosine_reg0 <= 36'sb11111000000000111100101001101000100;
            sine_reg0   <= 36'sb111000000100011110101000011101001001;
        end
        15732: begin
            cosine_reg0 <= 36'sb11111000000010100000001110100011011;
            sine_reg0   <= 36'sb111000000101001111010101010000010000;
        end
        15733: begin
            cosine_reg0 <= 36'sb11111000000100000011101001111010010;
            sine_reg0   <= 36'sb111000000110000000000010010110111010;
        end
        15734: begin
            cosine_reg0 <= 36'sb11111000000101100110111011101101001;
            sine_reg0   <= 36'sb111000000110110000101111110001000101;
        end
        15735: begin
            cosine_reg0 <= 36'sb11111000000111001010000011111011111;
            sine_reg0   <= 36'sb111000000111100001011101011110101110;
        end
        15736: begin
            cosine_reg0 <= 36'sb11111000001000101101000010100110011;
            sine_reg0   <= 36'sb111000001000010010001011011111110100;
        end
        15737: begin
            cosine_reg0 <= 36'sb11111000001010001111110111101100101;
            sine_reg0   <= 36'sb111000001001000010111001110100010101;
        end
        15738: begin
            cosine_reg0 <= 36'sb11111000001011110010100011001110101;
            sine_reg0   <= 36'sb111000001001110011101000011100001111;
        end
        15739: begin
            cosine_reg0 <= 36'sb11111000001101010101000101001100001;
            sine_reg0   <= 36'sb111000001010100100010111010111100000;
        end
        15740: begin
            cosine_reg0 <= 36'sb11111000001110110111011101100101011;
            sine_reg0   <= 36'sb111000001011010101000110100110000110;
        end
        15741: begin
            cosine_reg0 <= 36'sb11111000010000011001101100011010000;
            sine_reg0   <= 36'sb111000001100000101110110001000000000;
        end
        15742: begin
            cosine_reg0 <= 36'sb11111000010001111011110001101010001;
            sine_reg0   <= 36'sb111000001100110110100101111101001011;
        end
        15743: begin
            cosine_reg0 <= 36'sb11111000010011011101101101010101101;
            sine_reg0   <= 36'sb111000001101100111010110000101100110;
        end
        15744: begin
            cosine_reg0 <= 36'sb11111000010100111111011111011100100;
            sine_reg0   <= 36'sb111000001110011000000110100001001110;
        end
        15745: begin
            cosine_reg0 <= 36'sb11111000010110100001000111111110101;
            sine_reg0   <= 36'sb111000001111001000110111010000000010;
        end
        15746: begin
            cosine_reg0 <= 36'sb11111000011000000010100110111011111;
            sine_reg0   <= 36'sb111000001111111001101000010010000001;
        end
        15747: begin
            cosine_reg0 <= 36'sb11111000011001100011111100010100011;
            sine_reg0   <= 36'sb111000010000101010011001100111000111;
        end
        15748: begin
            cosine_reg0 <= 36'sb11111000011011000101001000001000000;
            sine_reg0   <= 36'sb111000010001011011001011001111010011;
        end
        15749: begin
            cosine_reg0 <= 36'sb11111000011100100110001010010110101;
            sine_reg0   <= 36'sb111000010010001011111101001010100100;
        end
        15750: begin
            cosine_reg0 <= 36'sb11111000011110000111000011000000010;
            sine_reg0   <= 36'sb111000010010111100101111011000110111;
        end
        15751: begin
            cosine_reg0 <= 36'sb11111000011111100111110010000100110;
            sine_reg0   <= 36'sb111000010011101101100001111010001011;
        end
        15752: begin
            cosine_reg0 <= 36'sb11111000100001001000010111100100001;
            sine_reg0   <= 36'sb111000010100011110010100101110011101;
        end
        15753: begin
            cosine_reg0 <= 36'sb11111000100010101000110011011110011;
            sine_reg0   <= 36'sb111000010101001111000111110101101101;
        end
        15754: begin
            cosine_reg0 <= 36'sb11111000100100001001000101110011011;
            sine_reg0   <= 36'sb111000010101111111111011001111110111;
        end
        15755: begin
            cosine_reg0 <= 36'sb11111000100101101001001110100011000;
            sine_reg0   <= 36'sb111000010110110000101110111100111010;
        end
        15756: begin
            cosine_reg0 <= 36'sb11111000100111001001001101101101010;
            sine_reg0   <= 36'sb111000010111100001100010111100110100;
        end
        15757: begin
            cosine_reg0 <= 36'sb11111000101000101001000011010010001;
            sine_reg0   <= 36'sb111000011000010010010111001111100100;
        end
        15758: begin
            cosine_reg0 <= 36'sb11111000101010001000101111010001100;
            sine_reg0   <= 36'sb111000011001000011001011110101000111;
        end
        15759: begin
            cosine_reg0 <= 36'sb11111000101011101000010001101011011;
            sine_reg0   <= 36'sb111000011001110100000000101101011011;
        end
        15760: begin
            cosine_reg0 <= 36'sb11111000101101000111101010011111101;
            sine_reg0   <= 36'sb111000011010100100110101111000011111;
        end
        15761: begin
            cosine_reg0 <= 36'sb11111000101110100110111001101110001;
            sine_reg0   <= 36'sb111000011011010101101011010110010001;
        end
        15762: begin
            cosine_reg0 <= 36'sb11111000110000000101111111010111000;
            sine_reg0   <= 36'sb111000011100000110100001000110101111;
        end
        15763: begin
            cosine_reg0 <= 36'sb11111000110001100100111011011010001;
            sine_reg0   <= 36'sb111000011100110111010111001001110110;
        end
        15764: begin
            cosine_reg0 <= 36'sb11111000110011000011101101110111100;
            sine_reg0   <= 36'sb111000011101101000001101011111100110;
        end
        15765: begin
            cosine_reg0 <= 36'sb11111000110100100010010110101110111;
            sine_reg0   <= 36'sb111000011110011001000100000111111100;
        end
        15766: begin
            cosine_reg0 <= 36'sb11111000110110000000110110000000010;
            sine_reg0   <= 36'sb111000011111001001111011000010110110;
        end
        15767: begin
            cosine_reg0 <= 36'sb11111000110111011111001011101011110;
            sine_reg0   <= 36'sb111000011111111010110010010000010011;
        end
        15768: begin
            cosine_reg0 <= 36'sb11111000111000111101010111110001001;
            sine_reg0   <= 36'sb111000100000101011101001110000010000;
        end
        15769: begin
            cosine_reg0 <= 36'sb11111000111010011011011010010000011;
            sine_reg0   <= 36'sb111000100001011100100001100010101100;
        end
        15770: begin
            cosine_reg0 <= 36'sb11111000111011111001010011001001100;
            sine_reg0   <= 36'sb111000100010001101011001100111100101;
        end
        15771: begin
            cosine_reg0 <= 36'sb11111000111101010111000010011100100;
            sine_reg0   <= 36'sb111000100010111110010001111110111000;
        end
        15772: begin
            cosine_reg0 <= 36'sb11111000111110110100101000001001000;
            sine_reg0   <= 36'sb111000100011101111001010101000100101;
        end
        15773: begin
            cosine_reg0 <= 36'sb11111001000000010010000100001111011;
            sine_reg0   <= 36'sb111000100100100000000011100100101001;
        end
        15774: begin
            cosine_reg0 <= 36'sb11111001000001101111010110101111010;
            sine_reg0   <= 36'sb111000100101010000111100110011000010;
        end
        15775: begin
            cosine_reg0 <= 36'sb11111001000011001100011111101000101;
            sine_reg0   <= 36'sb111000100110000001110110010011101110;
        end
        15776: begin
            cosine_reg0 <= 36'sb11111001000100101001011110111011101;
            sine_reg0   <= 36'sb111000100110110010110000000110101100;
        end
        15777: begin
            cosine_reg0 <= 36'sb11111001000110000110010100101000000;
            sine_reg0   <= 36'sb111000100111100011101010001011111001;
        end
        15778: begin
            cosine_reg0 <= 36'sb11111001000111100011000000101101101;
            sine_reg0   <= 36'sb111000101000010100100100100011010100;
        end
        15779: begin
            cosine_reg0 <= 36'sb11111001001000111111100011001100110;
            sine_reg0   <= 36'sb111000101001000101011111001100111011;
        end
        15780: begin
            cosine_reg0 <= 36'sb11111001001010011011111100000101001;
            sine_reg0   <= 36'sb111000101001110110011010001000101100;
        end
        15781: begin
            cosine_reg0 <= 36'sb11111001001011111000001011010110101;
            sine_reg0   <= 36'sb111000101010100111010101010110100101;
        end
        15782: begin
            cosine_reg0 <= 36'sb11111001001101010100010001000001011;
            sine_reg0   <= 36'sb111000101011011000010000110110100100;
        end
        15783: begin
            cosine_reg0 <= 36'sb11111001001110110000001101000101010;
            sine_reg0   <= 36'sb111000101100001001001100101000101000;
        end
        15784: begin
            cosine_reg0 <= 36'sb11111001010000001011111111100010001;
            sine_reg0   <= 36'sb111000101100111010001000101100101101;
        end
        15785: begin
            cosine_reg0 <= 36'sb11111001010001100111101000010111111;
            sine_reg0   <= 36'sb111000101101101011000101000010110100;
        end
        15786: begin
            cosine_reg0 <= 36'sb11111001010011000011000111100110110;
            sine_reg0   <= 36'sb111000101110011100000001101010111001;
        end
        15787: begin
            cosine_reg0 <= 36'sb11111001010100011110011101001110011;
            sine_reg0   <= 36'sb111000101111001100111110100100111010;
        end
        15788: begin
            cosine_reg0 <= 36'sb11111001010101111001101001001110111;
            sine_reg0   <= 36'sb111000101111111101111011110000110111;
        end
        15789: begin
            cosine_reg0 <= 36'sb11111001010111010100101011101000010;
            sine_reg0   <= 36'sb111000110000101110111001001110101100;
        end
        15790: begin
            cosine_reg0 <= 36'sb11111001011000101111100100011010010;
            sine_reg0   <= 36'sb111000110001011111110110111110011000;
        end
        15791: begin
            cosine_reg0 <= 36'sb11111001011010001010010011100100111;
            sine_reg0   <= 36'sb111000110010010000110100111111111010;
        end
        15792: begin
            cosine_reg0 <= 36'sb11111001011011100100111001001000001;
            sine_reg0   <= 36'sb111000110011000001110011010011001111;
        end
        15793: begin
            cosine_reg0 <= 36'sb11111001011100111111010101000100000;
            sine_reg0   <= 36'sb111000110011110010110001111000010101;
        end
        15794: begin
            cosine_reg0 <= 36'sb11111001011110011001100111011000010;
            sine_reg0   <= 36'sb111000110100100011110000101111001011;
        end
        15795: begin
            cosine_reg0 <= 36'sb11111001011111110011110000000101001;
            sine_reg0   <= 36'sb111000110101010100101111110111101111;
        end
        15796: begin
            cosine_reg0 <= 36'sb11111001100001001101101111001010010;
            sine_reg0   <= 36'sb111000110110000101101111010001111110;
        end
        15797: begin
            cosine_reg0 <= 36'sb11111001100010100111100100100111110;
            sine_reg0   <= 36'sb111000110110110110101110111101110111;
        end
        15798: begin
            cosine_reg0 <= 36'sb11111001100100000001010000011101100;
            sine_reg0   <= 36'sb111000110111100111101110111011011000;
        end
        15799: begin
            cosine_reg0 <= 36'sb11111001100101011010110010101011100;
            sine_reg0   <= 36'sb111000111000011000101111001010011111;
        end
        15800: begin
            cosine_reg0 <= 36'sb11111001100110110100001011010001110;
            sine_reg0   <= 36'sb111000111001001001101111101011001010;
        end
        15801: begin
            cosine_reg0 <= 36'sb11111001101000001101011010010000000;
            sine_reg0   <= 36'sb111000111001111010110000011101011000;
        end
        15802: begin
            cosine_reg0 <= 36'sb11111001101001100110011111100110011;
            sine_reg0   <= 36'sb111000111010101011110001100001000110;
        end
        15803: begin
            cosine_reg0 <= 36'sb11111001101010111111011011010100110;
            sine_reg0   <= 36'sb111000111011011100110010110110010010;
        end
        15804: begin
            cosine_reg0 <= 36'sb11111001101100011000001101011011001;
            sine_reg0   <= 36'sb111000111100001101110100011100111011;
        end
        15805: begin
            cosine_reg0 <= 36'sb11111001101101110000110101111001011;
            sine_reg0   <= 36'sb111000111100111110110110010100111111;
        end
        15806: begin
            cosine_reg0 <= 36'sb11111001101111001001010100101111100;
            sine_reg0   <= 36'sb111000111101101111111000011110011100;
        end
        15807: begin
            cosine_reg0 <= 36'sb11111001110000100001101001111101011;
            sine_reg0   <= 36'sb111000111110100000111010111001010000;
        end
        15808: begin
            cosine_reg0 <= 36'sb11111001110001111001110101100011000;
            sine_reg0   <= 36'sb111000111111010001111101100101011000;
        end
        15809: begin
            cosine_reg0 <= 36'sb11111001110011010001110111100000011;
            sine_reg0   <= 36'sb111001000000000011000000100010110100;
        end
        15810: begin
            cosine_reg0 <= 36'sb11111001110100101001101111110101011;
            sine_reg0   <= 36'sb111001000000110100000011110001100001;
        end
        15811: begin
            cosine_reg0 <= 36'sb11111001110110000001011110100001111;
            sine_reg0   <= 36'sb111001000001100101000111010001011110;
        end
        15812: begin
            cosine_reg0 <= 36'sb11111001110111011001000011100110000;
            sine_reg0   <= 36'sb111001000010010110001011000010101000;
        end
        15813: begin
            cosine_reg0 <= 36'sb11111001111000110000011111000001101;
            sine_reg0   <= 36'sb111001000011000111001111000100111110;
        end
        15814: begin
            cosine_reg0 <= 36'sb11111001111010000111110000110100101;
            sine_reg0   <= 36'sb111001000011111000010011011000011101;
        end
        15815: begin
            cosine_reg0 <= 36'sb11111001111011011110111000111111000;
            sine_reg0   <= 36'sb111001000100101001010111111101000100;
        end
        15816: begin
            cosine_reg0 <= 36'sb11111001111100110101110111100000110;
            sine_reg0   <= 36'sb111001000101011010011100110010110001;
        end
        15817: begin
            cosine_reg0 <= 36'sb11111001111110001100101100011001110;
            sine_reg0   <= 36'sb111001000110001011100001111001100010;
        end
        15818: begin
            cosine_reg0 <= 36'sb11111001111111100011010111101010000;
            sine_reg0   <= 36'sb111001000110111100100111010001010110;
        end
        15819: begin
            cosine_reg0 <= 36'sb11111010000000111001111001010001011;
            sine_reg0   <= 36'sb111001000111101101101100111010001001;
        end
        15820: begin
            cosine_reg0 <= 36'sb11111010000010010000010001001111110;
            sine_reg0   <= 36'sb111001001000011110110010110011111011;
        end
        15821: begin
            cosine_reg0 <= 36'sb11111010000011100110011111100101011;
            sine_reg0   <= 36'sb111001001001001111111000111110101001;
        end
        15822: begin
            cosine_reg0 <= 36'sb11111010000100111100100100010001111;
            sine_reg0   <= 36'sb111001001010000000111111011010010010;
        end
        15823: begin
            cosine_reg0 <= 36'sb11111010000110010010011111010101011;
            sine_reg0   <= 36'sb111001001010110010000110000110110100;
        end
        15824: begin
            cosine_reg0 <= 36'sb11111010000111101000010000101111111;
            sine_reg0   <= 36'sb111001001011100011001101000100001100;
        end
        15825: begin
            cosine_reg0 <= 36'sb11111010001000111101111000100001001;
            sine_reg0   <= 36'sb111001001100010100010100010010011010;
        end
        15826: begin
            cosine_reg0 <= 36'sb11111010001010010011010110101001010;
            sine_reg0   <= 36'sb111001001101000101011011110001011010;
        end
        15827: begin
            cosine_reg0 <= 36'sb11111010001011101000101011001000001;
            sine_reg0   <= 36'sb111001001101110110100011100001001011;
        end
        15828: begin
            cosine_reg0 <= 36'sb11111010001100111101110101111101101;
            sine_reg0   <= 36'sb111001001110100111101011100001101100;
        end
        15829: begin
            cosine_reg0 <= 36'sb11111010001110010010110111001001110;
            sine_reg0   <= 36'sb111001001111011000110011110010111010;
        end
        15830: begin
            cosine_reg0 <= 36'sb11111010001111100111101110101100101;
            sine_reg0   <= 36'sb111001010000001001111100010100110011;
        end
        15831: begin
            cosine_reg0 <= 36'sb11111010010000111100011100100110000;
            sine_reg0   <= 36'sb111001010000111011000101000111010110;
        end
        15832: begin
            cosine_reg0 <= 36'sb11111010010010010001000000110101110;
            sine_reg0   <= 36'sb111001010001101100001110001010100001;
        end
        15833: begin
            cosine_reg0 <= 36'sb11111010010011100101011011011100000;
            sine_reg0   <= 36'sb111001010010011101010111011110010001;
        end
        15834: begin
            cosine_reg0 <= 36'sb11111010010100111001101100011000110;
            sine_reg0   <= 36'sb111001010011001110100001000010100101;
        end
        15835: begin
            cosine_reg0 <= 36'sb11111010010110001101110011101011110;
            sine_reg0   <= 36'sb111001010011111111101010110111011100;
        end
        15836: begin
            cosine_reg0 <= 36'sb11111010010111100001110001010101000;
            sine_reg0   <= 36'sb111001010100110000110100111100110010;
        end
        15837: begin
            cosine_reg0 <= 36'sb11111010011000110101100101010100101;
            sine_reg0   <= 36'sb111001010101100001111111010010100110;
        end
        15838: begin
            cosine_reg0 <= 36'sb11111010011010001001001111101010011;
            sine_reg0   <= 36'sb111001010110010011001001111000110111;
        end
        15839: begin
            cosine_reg0 <= 36'sb11111010011011011100110000010110010;
            sine_reg0   <= 36'sb111001010111000100010100101111100010;
        end
        15840: begin
            cosine_reg0 <= 36'sb11111010011100110000000111011000010;
            sine_reg0   <= 36'sb111001010111110101011111110110100101;
        end
        15841: begin
            cosine_reg0 <= 36'sb11111010011110000011010100110000010;
            sine_reg0   <= 36'sb111001011000100110101011001101111111;
        end
        15842: begin
            cosine_reg0 <= 36'sb11111010011111010110011000011110010;
            sine_reg0   <= 36'sb111001011001010111110110110101101110;
        end
        15843: begin
            cosine_reg0 <= 36'sb11111010100000101001010010100010010;
            sine_reg0   <= 36'sb111001011010001001000010101101110000;
        end
        15844: begin
            cosine_reg0 <= 36'sb11111010100001111100000010111100000;
            sine_reg0   <= 36'sb111001011010111010001110110110000010;
        end
        15845: begin
            cosine_reg0 <= 36'sb11111010100011001110101001101011110;
            sine_reg0   <= 36'sb111001011011101011011011001110100011;
        end
        15846: begin
            cosine_reg0 <= 36'sb11111010100100100001000110110001010;
            sine_reg0   <= 36'sb111001011100011100100111110111010010;
        end
        15847: begin
            cosine_reg0 <= 36'sb11111010100101110011011010001100100;
            sine_reg0   <= 36'sb111001011101001101110100110000001100;
        end
        15848: begin
            cosine_reg0 <= 36'sb11111010100111000101100011111101011;
            sine_reg0   <= 36'sb111001011101111111000001111001001111;
        end
        15849: begin
            cosine_reg0 <= 36'sb11111010101000010111100100000011111;
            sine_reg0   <= 36'sb111001011110110000001111010010011001;
        end
        15850: begin
            cosine_reg0 <= 36'sb11111010101001101001011010100000000;
            sine_reg0   <= 36'sb111001011111100001011100111011101001;
        end
        15851: begin
            cosine_reg0 <= 36'sb11111010101010111011000111010001110;
            sine_reg0   <= 36'sb111001100000010010101010110100111101;
        end
        15852: begin
            cosine_reg0 <= 36'sb11111010101100001100101010011000111;
            sine_reg0   <= 36'sb111001100001000011111000111110010010;
        end
        15853: begin
            cosine_reg0 <= 36'sb11111010101101011110000011110101101;
            sine_reg0   <= 36'sb111001100001110101000111010111100111;
        end
        15854: begin
            cosine_reg0 <= 36'sb11111010101110101111010011100111101;
            sine_reg0   <= 36'sb111001100010100110010110000000111010;
        end
        15855: begin
            cosine_reg0 <= 36'sb11111010110000000000011001101111000;
            sine_reg0   <= 36'sb111001100011010111100100111010001001;
        end
        15856: begin
            cosine_reg0 <= 36'sb11111010110001010001010110001011101;
            sine_reg0   <= 36'sb111001100100001000110100000011010010;
        end
        15857: begin
            cosine_reg0 <= 36'sb11111010110010100010001000111101101;
            sine_reg0   <= 36'sb111001100100111010000011011100010100;
        end
        15858: begin
            cosine_reg0 <= 36'sb11111010110011110010110010000100110;
            sine_reg0   <= 36'sb111001100101101011010011000101001100;
        end
        15859: begin
            cosine_reg0 <= 36'sb11111010110101000011010001100001000;
            sine_reg0   <= 36'sb111001100110011100100010111101111000;
        end
        15860: begin
            cosine_reg0 <= 36'sb11111010110110010011100111010010011;
            sine_reg0   <= 36'sb111001100111001101110011000110010111;
        end
        15861: begin
            cosine_reg0 <= 36'sb11111010110111100011110011011000110;
            sine_reg0   <= 36'sb111001100111111111000011011110100110;
        end
        15862: begin
            cosine_reg0 <= 36'sb11111010111000110011110101110100010;
            sine_reg0   <= 36'sb111001101000110000010100000110100100;
        end
        15863: begin
            cosine_reg0 <= 36'sb11111010111010000011101110100100101;
            sine_reg0   <= 36'sb111001101001100001100100111110001111;
        end
        15864: begin
            cosine_reg0 <= 36'sb11111010111011010011011101101010000;
            sine_reg0   <= 36'sb111001101010010010110110000101100101;
        end
        15865: begin
            cosine_reg0 <= 36'sb11111010111100100011000011000100001;
            sine_reg0   <= 36'sb111001101011000100000111011100100100;
        end
        15866: begin
            cosine_reg0 <= 36'sb11111010111101110010011110110011001;
            sine_reg0   <= 36'sb111001101011110101011001000011001010;
        end
        15867: begin
            cosine_reg0 <= 36'sb11111010111111000001110000110110111;
            sine_reg0   <= 36'sb111001101100100110101010111001010101;
        end
        15868: begin
            cosine_reg0 <= 36'sb11111011000000010000111001001111011;
            sine_reg0   <= 36'sb111001101101010111111100111111000100;
        end
        15869: begin
            cosine_reg0 <= 36'sb11111011000001011111110111111100101;
            sine_reg0   <= 36'sb111001101110001001001111010100010100;
        end
        15870: begin
            cosine_reg0 <= 36'sb11111011000010101110101100111110011;
            sine_reg0   <= 36'sb111001101110111010100001111001000011;
        end
        15871: begin
            cosine_reg0 <= 36'sb11111011000011111101011000010100110;
            sine_reg0   <= 36'sb111001101111101011110100101101010001;
        end
        15872: begin
            cosine_reg0 <= 36'sb11111011000101001011111001111111101;
            sine_reg0   <= 36'sb111001110000011101000111110000111010;
        end
        15873: begin
            cosine_reg0 <= 36'sb11111011000110011010010001111111000;
            sine_reg0   <= 36'sb111001110001001110011011000011111100;
        end
        15874: begin
            cosine_reg0 <= 36'sb11111011000111101000100000010010110;
            sine_reg0   <= 36'sb111001110001111111101110100110010111;
        end
        15875: begin
            cosine_reg0 <= 36'sb11111011001000110110100100111011000;
            sine_reg0   <= 36'sb111001110010110001000010011000001000;
        end
        15876: begin
            cosine_reg0 <= 36'sb11111011001010000100011111110111100;
            sine_reg0   <= 36'sb111001110011100010010110011001001101;
        end
        15877: begin
            cosine_reg0 <= 36'sb11111011001011010010010001001000011;
            sine_reg0   <= 36'sb111001110100010011101010101001100100;
        end
        15878: begin
            cosine_reg0 <= 36'sb11111011001100011111111000101101011;
            sine_reg0   <= 36'sb111001110101000100111111001001001100;
        end
        15879: begin
            cosine_reg0 <= 36'sb11111011001101101101010110100110110;
            sine_reg0   <= 36'sb111001110101110110010011111000000001;
        end
        15880: begin
            cosine_reg0 <= 36'sb11111011001110111010101010110100001;
            sine_reg0   <= 36'sb111001110110100111101000110110000100;
        end
        15881: begin
            cosine_reg0 <= 36'sb11111011010000000111110101010101101;
            sine_reg0   <= 36'sb111001110111011000111110000011010001;
        end
        15882: begin
            cosine_reg0 <= 36'sb11111011010001010100110110001011010;
            sine_reg0   <= 36'sb111001111000001010010011011111100111;
        end
        15883: begin
            cosine_reg0 <= 36'sb11111011010010100001101101010100111;
            sine_reg0   <= 36'sb111001111000111011101001001011000011;
        end
        15884: begin
            cosine_reg0 <= 36'sb11111011010011101110011010110010100;
            sine_reg0   <= 36'sb111001111001101100111111000101100101;
        end
        15885: begin
            cosine_reg0 <= 36'sb11111011010100111010111110100100000;
            sine_reg0   <= 36'sb111001111010011110010101001111001010;
        end
        15886: begin
            cosine_reg0 <= 36'sb11111011010110000111011000101001011;
            sine_reg0   <= 36'sb111001111011001111101011100111101111;
        end
        15887: begin
            cosine_reg0 <= 36'sb11111011010111010011101001000010101;
            sine_reg0   <= 36'sb111001111100000001000010001111010100;
        end
        15888: begin
            cosine_reg0 <= 36'sb11111011011000011111101111101111100;
            sine_reg0   <= 36'sb111001111100110010011001000101110110;
        end
        15889: begin
            cosine_reg0 <= 36'sb11111011011001101011101100110000010;
            sine_reg0   <= 36'sb111001111101100011110000001011010100;
        end
        15890: begin
            cosine_reg0 <= 36'sb11111011011010110111100000000100110;
            sine_reg0   <= 36'sb111001111110010101000111011111101011;
        end
        15891: begin
            cosine_reg0 <= 36'sb11111011011100000011001001101100110;
            sine_reg0   <= 36'sb111001111111000110011111000010111010;
        end
        15892: begin
            cosine_reg0 <= 36'sb11111011011101001110101001101000100;
            sine_reg0   <= 36'sb111001111111110111110110110100111110;
        end
        15893: begin
            cosine_reg0 <= 36'sb11111011011110011001111111110111101;
            sine_reg0   <= 36'sb111010000000101001001110110101110111;
        end
        15894: begin
            cosine_reg0 <= 36'sb11111011011111100101001100011010011;
            sine_reg0   <= 36'sb111010000001011010100111000101100001;
        end
        15895: begin
            cosine_reg0 <= 36'sb11111011100000110000001111010000101;
            sine_reg0   <= 36'sb111010000010001011111111100011111011;
        end
        15896: begin
            cosine_reg0 <= 36'sb11111011100001111011001000011010010;
            sine_reg0   <= 36'sb111010000010111101011000010001000011;
        end
        15897: begin
            cosine_reg0 <= 36'sb11111011100011000101110111110111010;
            sine_reg0   <= 36'sb111010000011101110110001001100110111;
        end
        15898: begin
            cosine_reg0 <= 36'sb11111011100100010000011101100111100;
            sine_reg0   <= 36'sb111010000100100000001010010111010110;
        end
        15899: begin
            cosine_reg0 <= 36'sb11111011100101011010111001101011001;
            sine_reg0   <= 36'sb111010000101010001100011110000011101;
        end
        15900: begin
            cosine_reg0 <= 36'sb11111011100110100101001100000010000;
            sine_reg0   <= 36'sb111010000110000010111101011000001011;
        end
        15901: begin
            cosine_reg0 <= 36'sb11111011100111101111010100101100000;
            sine_reg0   <= 36'sb111010000110110100010111001110011101;
        end
        15902: begin
            cosine_reg0 <= 36'sb11111011101000111001010011101001010;
            sine_reg0   <= 36'sb111010000111100101110001010011010001;
        end
        15903: begin
            cosine_reg0 <= 36'sb11111011101010000011001000111001100;
            sine_reg0   <= 36'sb111010001000010111001011100110100111;
        end
        15904: begin
            cosine_reg0 <= 36'sb11111011101011001100110100011100111;
            sine_reg0   <= 36'sb111010001001001000100110001000011011;
        end
        15905: begin
            cosine_reg0 <= 36'sb11111011101100010110010110010011010;
            sine_reg0   <= 36'sb111010001001111010000000111000101100;
        end
        15906: begin
            cosine_reg0 <= 36'sb11111011101101011111101110011100101;
            sine_reg0   <= 36'sb111010001010101011011011110111011001;
        end
        15907: begin
            cosine_reg0 <= 36'sb11111011101110101000111100111000111;
            sine_reg0   <= 36'sb111010001011011100110111000100011110;
        end
        15908: begin
            cosine_reg0 <= 36'sb11111011101111110010000001101000001;
            sine_reg0   <= 36'sb111010001100001110010010011111111011;
        end
        15909: begin
            cosine_reg0 <= 36'sb11111011110000111010111100101010001;
            sine_reg0   <= 36'sb111010001100111111101110001001101101;
        end
        15910: begin
            cosine_reg0 <= 36'sb11111011110010000011101101111110111;
            sine_reg0   <= 36'sb111010001101110001001010000001110010;
        end
        15911: begin
            cosine_reg0 <= 36'sb11111011110011001100010101100110011;
            sine_reg0   <= 36'sb111010001110100010100110001000001001;
        end
        15912: begin
            cosine_reg0 <= 36'sb11111011110100010100110011100000110;
            sine_reg0   <= 36'sb111010001111010100000010011100110000;
        end
        15913: begin
            cosine_reg0 <= 36'sb11111011110101011101000111101101101;
            sine_reg0   <= 36'sb111010010000000101011110111111100100;
        end
        15914: begin
            cosine_reg0 <= 36'sb11111011110110100101010010001101001;
            sine_reg0   <= 36'sb111010010000110110111011110000100100;
        end
        15915: begin
            cosine_reg0 <= 36'sb11111011110111101101010010111111010;
            sine_reg0   <= 36'sb111010010001101000011000101111101110;
        end
        15916: begin
            cosine_reg0 <= 36'sb11111011111000110101001010000100000;
            sine_reg0   <= 36'sb111010010010011001110101111101000000;
        end
        15917: begin
            cosine_reg0 <= 36'sb11111011111001111100110111011011001;
            sine_reg0   <= 36'sb111010010011001011010011011000011000;
        end
        15918: begin
            cosine_reg0 <= 36'sb11111011111011000100011011000100110;
            sine_reg0   <= 36'sb111010010011111100110001000001110100;
        end
        15919: begin
            cosine_reg0 <= 36'sb11111011111100001011110101000000110;
            sine_reg0   <= 36'sb111010010100101110001110111001010010;
        end
        15920: begin
            cosine_reg0 <= 36'sb11111011111101010011000101001111001;
            sine_reg0   <= 36'sb111010010101011111101100111110110001;
        end
        15921: begin
            cosine_reg0 <= 36'sb11111011111110011010001011101111110;
            sine_reg0   <= 36'sb111010010110010001001011010010001110;
        end
        15922: begin
            cosine_reg0 <= 36'sb11111011111111100001001000100010110;
            sine_reg0   <= 36'sb111010010111000010101001110011101000;
        end
        15923: begin
            cosine_reg0 <= 36'sb11111100000000100111111011100111111;
            sine_reg0   <= 36'sb111010010111110100001000100010111100;
        end
        15924: begin
            cosine_reg0 <= 36'sb11111100000001101110100100111111010;
            sine_reg0   <= 36'sb111010011000100101100111100000001001;
        end
        15925: begin
            cosine_reg0 <= 36'sb11111100000010110101000100101000111;
            sine_reg0   <= 36'sb111010011001010111000110101011001101;
        end
        15926: begin
            cosine_reg0 <= 36'sb11111100000011111011011010100100100;
            sine_reg0   <= 36'sb111010011010001000100110000100000110;
        end
        15927: begin
            cosine_reg0 <= 36'sb11111100000101000001100110110010001;
            sine_reg0   <= 36'sb111010011010111010000101101010110001;
        end
        15928: begin
            cosine_reg0 <= 36'sb11111100000110000111101001010001111;
            sine_reg0   <= 36'sb111010011011101011100101011111001110;
        end
        15929: begin
            cosine_reg0 <= 36'sb11111100000111001101100010000011101;
            sine_reg0   <= 36'sb111010011100011101000101100001011010;
        end
        15930: begin
            cosine_reg0 <= 36'sb11111100001000010011010001000111010;
            sine_reg0   <= 36'sb111010011101001110100101110001010100;
        end
        15931: begin
            cosine_reg0 <= 36'sb11111100001001011000110110011100110;
            sine_reg0   <= 36'sb111010011110000000000110001110111000;
        end
        15932: begin
            cosine_reg0 <= 36'sb11111100001010011110010010000100001;
            sine_reg0   <= 36'sb111010011110110001100110111010000111;
        end
        15933: begin
            cosine_reg0 <= 36'sb11111100001011100011100011111101011;
            sine_reg0   <= 36'sb111010011111100011000111110010111100;
        end
        15934: begin
            cosine_reg0 <= 36'sb11111100001100101000101100001000011;
            sine_reg0   <= 36'sb111010100000010100101000111001011000;
        end
        15935: begin
            cosine_reg0 <= 36'sb11111100001101101101101010100101000;
            sine_reg0   <= 36'sb111010100001000110001010001101010111;
        end
        15936: begin
            cosine_reg0 <= 36'sb11111100001110110010011111010011011;
            sine_reg0   <= 36'sb111010100001110111101011101110110111;
        end
        15937: begin
            cosine_reg0 <= 36'sb11111100001111110111001010010011100;
            sine_reg0   <= 36'sb111010100010101001001101011101111000;
        end
        15938: begin
            cosine_reg0 <= 36'sb11111100010000111011101011100101001;
            sine_reg0   <= 36'sb111010100011011010101111011010010111;
        end
        15939: begin
            cosine_reg0 <= 36'sb11111100010010000000000011001000010;
            sine_reg0   <= 36'sb111010100100001100010001100100010010;
        end
        15940: begin
            cosine_reg0 <= 36'sb11111100010011000100010000111101000;
            sine_reg0   <= 36'sb111010100100111101110011111011100111;
        end
        15941: begin
            cosine_reg0 <= 36'sb11111100010100001000010101000011001;
            sine_reg0   <= 36'sb111010100101101111010110100000010100;
        end
        15942: begin
            cosine_reg0 <= 36'sb11111100010101001100001111011010110;
            sine_reg0   <= 36'sb111010100110100000111001010010011000;
        end
        15943: begin
            cosine_reg0 <= 36'sb11111100010110010000000000000011111;
            sine_reg0   <= 36'sb111010100111010010011100010001110000;
        end
        15944: begin
            cosine_reg0 <= 36'sb11111100010111010011100110111110010;
            sine_reg0   <= 36'sb111010101000000011111111011110011011;
        end
        15945: begin
            cosine_reg0 <= 36'sb11111100011000010111000100001001111;
            sine_reg0   <= 36'sb111010101000110101100010111000010110;
        end
        15946: begin
            cosine_reg0 <= 36'sb11111100011001011010010111100110111;
            sine_reg0   <= 36'sb111010101001100111000110011111100000;
        end
        15947: begin
            cosine_reg0 <= 36'sb11111100011010011101100001010101001;
            sine_reg0   <= 36'sb111010101010011000101010010011110111;
        end
        15948: begin
            cosine_reg0 <= 36'sb11111100011011100000100001010100100;
            sine_reg0   <= 36'sb111010101011001010001110010101011001;
        end
        15949: begin
            cosine_reg0 <= 36'sb11111100011100100011010111100101001;
            sine_reg0   <= 36'sb111010101011111011110010100100000100;
        end
        15950: begin
            cosine_reg0 <= 36'sb11111100011101100110000100000110110;
            sine_reg0   <= 36'sb111010101100101101010110111111110101;
        end
        15951: begin
            cosine_reg0 <= 36'sb11111100011110101000100110111001100;
            sine_reg0   <= 36'sb111010101101011110111011101000101100;
        end
        15952: begin
            cosine_reg0 <= 36'sb11111100011111101010111111111101011;
            sine_reg0   <= 36'sb111010101110010000100000011110100111;
        end
        15953: begin
            cosine_reg0 <= 36'sb11111100100000101101001111010010001;
            sine_reg0   <= 36'sb111010101111000010000101100001100010;
        end
        15954: begin
            cosine_reg0 <= 36'sb11111100100001101111010100110111111;
            sine_reg0   <= 36'sb111010101111110011101010110001011101;
        end
        15955: begin
            cosine_reg0 <= 36'sb11111100100010110001010000101110100;
            sine_reg0   <= 36'sb111010110000100101010000001110010110;
        end
        15956: begin
            cosine_reg0 <= 36'sb11111100100011110011000010110110000;
            sine_reg0   <= 36'sb111010110001010110110101111000001010;
        end
        15957: begin
            cosine_reg0 <= 36'sb11111100100100110100101011001110011;
            sine_reg0   <= 36'sb111010110010001000011011101110111000;
        end
        15958: begin
            cosine_reg0 <= 36'sb11111100100101110110001001110111100;
            sine_reg0   <= 36'sb111010110010111010000001110010011110;
        end
        15959: begin
            cosine_reg0 <= 36'sb11111100100110110111011110110001011;
            sine_reg0   <= 36'sb111010110011101011101000000010111001;
        end
        15960: begin
            cosine_reg0 <= 36'sb11111100100111111000101001111100000;
            sine_reg0   <= 36'sb111010110100011101001110100000001001;
        end
        15961: begin
            cosine_reg0 <= 36'sb11111100101000111001101011010111011;
            sine_reg0   <= 36'sb111010110101001110110101001010001010;
        end
        15962: begin
            cosine_reg0 <= 36'sb11111100101001111010100011000011010;
            sine_reg0   <= 36'sb111010110110000000011100000000111100;
        end
        15963: begin
            cosine_reg0 <= 36'sb11111100101010111011010000111111111;
            sine_reg0   <= 36'sb111010110110110010000011000100011100;
        end
        15964: begin
            cosine_reg0 <= 36'sb11111100101011111011110101001100111;
            sine_reg0   <= 36'sb111010110111100011101010010100101000;
        end
        15965: begin
            cosine_reg0 <= 36'sb11111100101100111100001111101010100;
            sine_reg0   <= 36'sb111010111000010101010001110001011110;
        end
        15966: begin
            cosine_reg0 <= 36'sb11111100101101111100100000011000101;
            sine_reg0   <= 36'sb111010111001000110111001011010111110;
        end
        15967: begin
            cosine_reg0 <= 36'sb11111100101110111100100111010111010;
            sine_reg0   <= 36'sb111010111001111000100001010001000011;
        end
        15968: begin
            cosine_reg0 <= 36'sb11111100101111111100100100100110001;
            sine_reg0   <= 36'sb111010111010101010001001010011101110;
        end
        15969: begin
            cosine_reg0 <= 36'sb11111100110000111100011000000101100;
            sine_reg0   <= 36'sb111010111011011011110001100010111011;
        end
        15970: begin
            cosine_reg0 <= 36'sb11111100110001111100000001110101001;
            sine_reg0   <= 36'sb111010111100001101011001111110101001;
        end
        15971: begin
            cosine_reg0 <= 36'sb11111100110010111011100001110101000;
            sine_reg0   <= 36'sb111010111100111111000010100110110101;
        end
        15972: begin
            cosine_reg0 <= 36'sb11111100110011111010111000000101010;
            sine_reg0   <= 36'sb111010111101110000101011011011011111;
        end
        15973: begin
            cosine_reg0 <= 36'sb11111100110100111010000100100101101;
            sine_reg0   <= 36'sb111010111110100010010100011100100100;
        end
        15974: begin
            cosine_reg0 <= 36'sb11111100110101111001000111010110010;
            sine_reg0   <= 36'sb111010111111010011111101101010000010;
        end
        15975: begin
            cosine_reg0 <= 36'sb11111100110110111000000000010110111;
            sine_reg0   <= 36'sb111011000000000101100111000011111000;
        end
        15976: begin
            cosine_reg0 <= 36'sb11111100110111110110101111100111110;
            sine_reg0   <= 36'sb111011000000110111010000101010000010;
        end
        15977: begin
            cosine_reg0 <= 36'sb11111100111000110101010101001000101;
            sine_reg0   <= 36'sb111011000001101000111010011100100001;
        end
        15978: begin
            cosine_reg0 <= 36'sb11111100111001110011110000111001100;
            sine_reg0   <= 36'sb111011000010011010100100011011010000;
        end
        15979: begin
            cosine_reg0 <= 36'sb11111100111010110010000010111010011;
            sine_reg0   <= 36'sb111011000011001100001110100110010000;
        end
        15980: begin
            cosine_reg0 <= 36'sb11111100111011110000001011001011010;
            sine_reg0   <= 36'sb111011000011111101111000111101011101;
        end
        15981: begin
            cosine_reg0 <= 36'sb11111100111100101110001001101100000;
            sine_reg0   <= 36'sb111011000100101111100011100000110101;
        end
        15982: begin
            cosine_reg0 <= 36'sb11111100111101101011111110011100101;
            sine_reg0   <= 36'sb111011000101100001001110010000011000;
        end
        15983: begin
            cosine_reg0 <= 36'sb11111100111110101001101001011101000;
            sine_reg0   <= 36'sb111011000110010010111001001100000011;
        end
        15984: begin
            cosine_reg0 <= 36'sb11111100111111100111001010101101010;
            sine_reg0   <= 36'sb111011000111000100100100010011110011;
        end
        15985: begin
            cosine_reg0 <= 36'sb11111101000000100100100010001101011;
            sine_reg0   <= 36'sb111011000111110110001111100111101000;
        end
        15986: begin
            cosine_reg0 <= 36'sb11111101000001100001101111111101001;
            sine_reg0   <= 36'sb111011001000100111111011000111011111;
        end
        15987: begin
            cosine_reg0 <= 36'sb11111101000010011110110011111100100;
            sine_reg0   <= 36'sb111011001001011001100110110011010110;
        end
        15988: begin
            cosine_reg0 <= 36'sb11111101000011011011101110001011101;
            sine_reg0   <= 36'sb111011001010001011010010101011001100;
        end
        15989: begin
            cosine_reg0 <= 36'sb11111101000100011000011110101010010;
            sine_reg0   <= 36'sb111011001010111100111110101110111110;
        end
        15990: begin
            cosine_reg0 <= 36'sb11111101000101010101000101011000100;
            sine_reg0   <= 36'sb111011001011101110101010111110101011;
        end
        15991: begin
            cosine_reg0 <= 36'sb11111101000110010001100010010110011;
            sine_reg0   <= 36'sb111011001100100000010111011010010000;
        end
        15992: begin
            cosine_reg0 <= 36'sb11111101000111001101110101100011110;
            sine_reg0   <= 36'sb111011001101010010000100000001101100;
        end
        15993: begin
            cosine_reg0 <= 36'sb11111101001000001001111111000000100;
            sine_reg0   <= 36'sb111011001110000011110000110100111101;
        end
        15994: begin
            cosine_reg0 <= 36'sb11111101001001000101111110101100110;
            sine_reg0   <= 36'sb111011001110110101011101110100000000;
        end
        15995: begin
            cosine_reg0 <= 36'sb11111101001010000001110100101000011;
            sine_reg0   <= 36'sb111011001111100111001010111110110101;
        end
        15996: begin
            cosine_reg0 <= 36'sb11111101001010111101100000110011011;
            sine_reg0   <= 36'sb111011010000011000111000010101011000;
        end
        15997: begin
            cosine_reg0 <= 36'sb11111101001011111001000011001101101;
            sine_reg0   <= 36'sb111011010001001010100101110111101001;
        end
        15998: begin
            cosine_reg0 <= 36'sb11111101001100110100011011110111010;
            sine_reg0   <= 36'sb111011010001111100010011100101100101;
        end
        15999: begin
            cosine_reg0 <= 36'sb11111101001101101111101010110000001;
            sine_reg0   <= 36'sb111011010010101110000001011111001011;
        end
        16000: begin
            cosine_reg0 <= 36'sb11111101001110101010101111111000001;
            sine_reg0   <= 36'sb111011010011011111101111100100010111;
        end
        16001: begin
            cosine_reg0 <= 36'sb11111101001111100101101011001111011;
            sine_reg0   <= 36'sb111011010100010001011101110101001001;
        end
        16002: begin
            cosine_reg0 <= 36'sb11111101010000100000011100110101110;
            sine_reg0   <= 36'sb111011010101000011001100010001011111;
        end
        16003: begin
            cosine_reg0 <= 36'sb11111101010001011011000100101011010;
            sine_reg0   <= 36'sb111011010101110100111010111001010110;
        end
        16004: begin
            cosine_reg0 <= 36'sb11111101010010010101100010101111111;
            sine_reg0   <= 36'sb111011010110100110101001101100101101;
        end
        16005: begin
            cosine_reg0 <= 36'sb11111101010011001111110111000011100;
            sine_reg0   <= 36'sb111011010111011000011000101011100010;
        end
        16006: begin
            cosine_reg0 <= 36'sb11111101010100001010000001100110001;
            sine_reg0   <= 36'sb111011011000001010000111110101110011;
        end
        16007: begin
            cosine_reg0 <= 36'sb11111101010101000100000010010111110;
            sine_reg0   <= 36'sb111011011000111011110111001011011110;
        end
        16008: begin
            cosine_reg0 <= 36'sb11111101010101111101111001011000010;
            sine_reg0   <= 36'sb111011011001101101100110101100100000;
        end
        16009: begin
            cosine_reg0 <= 36'sb11111101010110110111100110100111110;
            sine_reg0   <= 36'sb111011011010011111010110011000111001;
        end
        16010: begin
            cosine_reg0 <= 36'sb11111101010111110001001010000110000;
            sine_reg0   <= 36'sb111011011011010001000110010000100110;
        end
        16011: begin
            cosine_reg0 <= 36'sb11111101011000101010100011110011001;
            sine_reg0   <= 36'sb111011011100000010110110010011100110;
        end
        16012: begin
            cosine_reg0 <= 36'sb11111101011001100011110011101111001;
            sine_reg0   <= 36'sb111011011100110100100110100001110101;
        end
        16013: begin
            cosine_reg0 <= 36'sb11111101011010011100111001111001110;
            sine_reg0   <= 36'sb111011011101100110010110111011010011;
        end
        16014: begin
            cosine_reg0 <= 36'sb11111101011011010101110110010011010;
            sine_reg0   <= 36'sb111011011110011000000111011111111110;
        end
        16015: begin
            cosine_reg0 <= 36'sb11111101011100001110101000111011011;
            sine_reg0   <= 36'sb111011011111001001111000001111110011;
        end
        16016: begin
            cosine_reg0 <= 36'sb11111101011101000111010001110010001;
            sine_reg0   <= 36'sb111011011111111011101001001010110001;
        end
        16017: begin
            cosine_reg0 <= 36'sb11111101011101111111110000110111100;
            sine_reg0   <= 36'sb111011100000101101011010010000110110;
        end
        16018: begin
            cosine_reg0 <= 36'sb11111101011110111000000110001011100;
            sine_reg0   <= 36'sb111011100001011111001011100010000000;
        end
        16019: begin
            cosine_reg0 <= 36'sb11111101011111110000010001101110000;
            sine_reg0   <= 36'sb111011100010010000111100111110001100;
        end
        16020: begin
            cosine_reg0 <= 36'sb11111101100000101000010011011111001;
            sine_reg0   <= 36'sb111011100011000010101110100101011010;
        end
        16021: begin
            cosine_reg0 <= 36'sb11111101100001100000001011011110101;
            sine_reg0   <= 36'sb111011100011110100100000010111100111;
        end
        16022: begin
            cosine_reg0 <= 36'sb11111101100010010111111001101100101;
            sine_reg0   <= 36'sb111011100100100110010010010100110001;
        end
        16023: begin
            cosine_reg0 <= 36'sb11111101100011001111011110001001001;
            sine_reg0   <= 36'sb111011100101011000000100011100110110;
        end
        16024: begin
            cosine_reg0 <= 36'sb11111101100100000110111000110011111;
            sine_reg0   <= 36'sb111011100110001001110110101111110100;
        end
        16025: begin
            cosine_reg0 <= 36'sb11111101100100111110001001101101001;
            sine_reg0   <= 36'sb111011100110111011101001001101101010;
        end
        16026: begin
            cosine_reg0 <= 36'sb11111101100101110101010000110100101;
            sine_reg0   <= 36'sb111011100111101101011011110110010110;
        end
        16027: begin
            cosine_reg0 <= 36'sb11111101100110101100001110001010011;
            sine_reg0   <= 36'sb111011101000011111001110101001110101;
        end
        16028: begin
            cosine_reg0 <= 36'sb11111101100111100011000001101110100;
            sine_reg0   <= 36'sb111011101001010001000001101000000101;
        end
        16029: begin
            cosine_reg0 <= 36'sb11111101101000011001101011100000110;
            sine_reg0   <= 36'sb111011101010000010110100110001000110;
        end
        16030: begin
            cosine_reg0 <= 36'sb11111101101001010000001011100001010;
            sine_reg0   <= 36'sb111011101010110100101000000100110100;
        end
        16031: begin
            cosine_reg0 <= 36'sb11111101101010000110100001101111111;
            sine_reg0   <= 36'sb111011101011100110011011100011001110;
        end
        16032: begin
            cosine_reg0 <= 36'sb11111101101010111100101110001100100;
            sine_reg0   <= 36'sb111011101100011000001111001100010010;
        end
        16033: begin
            cosine_reg0 <= 36'sb11111101101011110010110000110111011;
            sine_reg0   <= 36'sb111011101101001010000010111111111111;
        end
        16034: begin
            cosine_reg0 <= 36'sb11111101101100101000101001110000010;
            sine_reg0   <= 36'sb111011101101111011110110111110010001;
        end
        16035: begin
            cosine_reg0 <= 36'sb11111101101101011110011000110111010;
            sine_reg0   <= 36'sb111011101110101101101011000111001000;
        end
        16036: begin
            cosine_reg0 <= 36'sb11111101101110010011111110001100001;
            sine_reg0   <= 36'sb111011101111011111011111011010100001;
        end
        16037: begin
            cosine_reg0 <= 36'sb11111101101111001001011001101111000;
            sine_reg0   <= 36'sb111011110000010001010011111000011010;
        end
        16038: begin
            cosine_reg0 <= 36'sb11111101101111111110101011011111110;
            sine_reg0   <= 36'sb111011110001000011001000100000110010;
        end
        16039: begin
            cosine_reg0 <= 36'sb11111101110000110011110011011110100;
            sine_reg0   <= 36'sb111011110001110100111101010011100110;
        end
        16040: begin
            cosine_reg0 <= 36'sb11111101110001101000110001101011001;
            sine_reg0   <= 36'sb111011110010100110110010010000110101;
        end
        16041: begin
            cosine_reg0 <= 36'sb11111101110010011101100110000101100;
            sine_reg0   <= 36'sb111011110011011000100111011000011101;
        end
        16042: begin
            cosine_reg0 <= 36'sb11111101110011010010010000101101110;
            sine_reg0   <= 36'sb111011110100001010011100101010011011;
        end
        16043: begin
            cosine_reg0 <= 36'sb11111101110100000110110001100011101;
            sine_reg0   <= 36'sb111011110100111100010010000110101110;
        end
        16044: begin
            cosine_reg0 <= 36'sb11111101110100111011001000100111011;
            sine_reg0   <= 36'sb111011110101101110000111101101010101;
        end
        16045: begin
            cosine_reg0 <= 36'sb11111101110101101111010101111000110;
            sine_reg0   <= 36'sb111011110110011111111101011110001100;
        end
        16046: begin
            cosine_reg0 <= 36'sb11111101110110100011011001010111111;
            sine_reg0   <= 36'sb111011110111010001110011011001010010;
        end
        16047: begin
            cosine_reg0 <= 36'sb11111101110111010111010011000100101;
            sine_reg0   <= 36'sb111011111000000011101001011110100110;
        end
        16048: begin
            cosine_reg0 <= 36'sb11111101111000001011000010111111000;
            sine_reg0   <= 36'sb111011111000110101011111101110000100;
        end
        16049: begin
            cosine_reg0 <= 36'sb11111101111000111110101001000111000;
            sine_reg0   <= 36'sb111011111001100111010110000111101101;
        end
        16050: begin
            cosine_reg0 <= 36'sb11111101111001110010000101011100011;
            sine_reg0   <= 36'sb111011111010011001001100101011011100;
        end
        16051: begin
            cosine_reg0 <= 36'sb11111101111010100101010111111111100;
            sine_reg0   <= 36'sb111011111011001011000011011001010001;
        end
        16052: begin
            cosine_reg0 <= 36'sb11111101111011011000100000110000000;
            sine_reg0   <= 36'sb111011111011111100111010010001001010;
        end
        16053: begin
            cosine_reg0 <= 36'sb11111101111100001011011111101101111;
            sine_reg0   <= 36'sb111011111100101110110001010011000100;
        end
        16054: begin
            cosine_reg0 <= 36'sb11111101111100111110010100111001010;
            sine_reg0   <= 36'sb111011111101100000101000011110111110;
        end
        16055: begin
            cosine_reg0 <= 36'sb11111101111101110001000000010010000;
            sine_reg0   <= 36'sb111011111110010010011111110100110110;
        end
        16056: begin
            cosine_reg0 <= 36'sb11111101111110100011100001111000010;
            sine_reg0   <= 36'sb111011111111000100010111010100101001;
        end
        16057: begin
            cosine_reg0 <= 36'sb11111101111111010101111001101011110;
            sine_reg0   <= 36'sb111011111111110110001110111110010111;
        end
        16058: begin
            cosine_reg0 <= 36'sb11111110000000001000000111101100100;
            sine_reg0   <= 36'sb111100000000101000000110110001111100;
        end
        16059: begin
            cosine_reg0 <= 36'sb11111110000000111010001011111010100;
            sine_reg0   <= 36'sb111100000001011001111110101111011000;
        end
        16060: begin
            cosine_reg0 <= 36'sb11111110000001101100000110010101111;
            sine_reg0   <= 36'sb111100000010001011110110110110101000;
        end
        16061: begin
            cosine_reg0 <= 36'sb11111110000010011101110110111110011;
            sine_reg0   <= 36'sb111100000010111101101111000111101010;
        end
        16062: begin
            cosine_reg0 <= 36'sb11111110000011001111011101110100001;
            sine_reg0   <= 36'sb111100000011101111100111100010011101;
        end
        16063: begin
            cosine_reg0 <= 36'sb11111110000100000000111010110111000;
            sine_reg0   <= 36'sb111100000100100001100000000110111101;
        end
        16064: begin
            cosine_reg0 <= 36'sb11111110000100110010001110000110111;
            sine_reg0   <= 36'sb111100000101010011011000110101001011;
        end
        16065: begin
            cosine_reg0 <= 36'sb11111110000101100011010111100100000;
            sine_reg0   <= 36'sb111100000110000101010001101101000011;
        end
        16066: begin
            cosine_reg0 <= 36'sb11111110000110010100010111001110001;
            sine_reg0   <= 36'sb111100000110110111001010101110100011;
        end
        16067: begin
            cosine_reg0 <= 36'sb11111110000111000101001101000101011;
            sine_reg0   <= 36'sb111100000111101001000011111001101011;
        end
        16068: begin
            cosine_reg0 <= 36'sb11111110000111110101111001001001100;
            sine_reg0   <= 36'sb111100001000011010111101001110010111;
        end
        16069: begin
            cosine_reg0 <= 36'sb11111110001000100110011011011010110;
            sine_reg0   <= 36'sb111100001001001100110110101100100110;
        end
        16070: begin
            cosine_reg0 <= 36'sb11111110001001010110110011111000111;
            sine_reg0   <= 36'sb111100001001111110110000010100010110;
        end
        16071: begin
            cosine_reg0 <= 36'sb11111110001010000111000010100011111;
            sine_reg0   <= 36'sb111100001010110000101010000101100101;
        end
        16072: begin
            cosine_reg0 <= 36'sb11111110001010110111000111011011110;
            sine_reg0   <= 36'sb111100001011100010100100000000010001;
        end
        16073: begin
            cosine_reg0 <= 36'sb11111110001011100111000010100000101;
            sine_reg0   <= 36'sb111100001100010100011110000100011000;
        end
        16074: begin
            cosine_reg0 <= 36'sb11111110001100010110110011110010010;
            sine_reg0   <= 36'sb111100001101000110011000010001111001;
        end
        16075: begin
            cosine_reg0 <= 36'sb11111110001101000110011011010000101;
            sine_reg0   <= 36'sb111100001101111000010010101000110001;
        end
        16076: begin
            cosine_reg0 <= 36'sb11111110001101110101111000111011111;
            sine_reg0   <= 36'sb111100001110101010001101001000111110;
        end
        16077: begin
            cosine_reg0 <= 36'sb11111110001110100101001100110011110;
            sine_reg0   <= 36'sb111100001111011100000111110010011111;
        end
        16078: begin
            cosine_reg0 <= 36'sb11111110001111010100010110111000100;
            sine_reg0   <= 36'sb111100010000001110000010100101010001;
        end
        16079: begin
            cosine_reg0 <= 36'sb11111110010000000011010111001001111;
            sine_reg0   <= 36'sb111100010000111111111101100001010011;
        end
        16080: begin
            cosine_reg0 <= 36'sb11111110010000110010001101100111111;
            sine_reg0   <= 36'sb111100010001110001111000100110100011;
        end
        16081: begin
            cosine_reg0 <= 36'sb11111110010001100000111010010010100;
            sine_reg0   <= 36'sb111100010010100011110011110100111110;
        end
        16082: begin
            cosine_reg0 <= 36'sb11111110010010001111011101001001110;
            sine_reg0   <= 36'sb111100010011010101101111001100100011;
        end
        16083: begin
            cosine_reg0 <= 36'sb11111110010010111101110110001101101;
            sine_reg0   <= 36'sb111100010100000111101010101101010001;
        end
        16084: begin
            cosine_reg0 <= 36'sb11111110010011101100000101011110000;
            sine_reg0   <= 36'sb111100010100111001100110010111000100;
        end
        16085: begin
            cosine_reg0 <= 36'sb11111110010100011010001010111010111;
            sine_reg0   <= 36'sb111100010101101011100010001001111011;
        end
        16086: begin
            cosine_reg0 <= 36'sb11111110010101001000000110100100010;
            sine_reg0   <= 36'sb111100010110011101011110000101110101;
        end
        16087: begin
            cosine_reg0 <= 36'sb11111110010101110101111000011010001;
            sine_reg0   <= 36'sb111100010111001111011010001010101111;
        end
        16088: begin
            cosine_reg0 <= 36'sb11111110010110100011100000011100011;
            sine_reg0   <= 36'sb111100011000000001010110011000100111;
        end
        16089: begin
            cosine_reg0 <= 36'sb11111110010111010000111110101011001;
            sine_reg0   <= 36'sb111100011000110011010010101111011011;
        end
        16090: begin
            cosine_reg0 <= 36'sb11111110010111111110010011000110010;
            sine_reg0   <= 36'sb111100011001100101001111001111001010;
        end
        16091: begin
            cosine_reg0 <= 36'sb11111110011000101011011101101101101;
            sine_reg0   <= 36'sb111100011010010111001011110111110001;
        end
        16092: begin
            cosine_reg0 <= 36'sb11111110011001011000011110100001100;
            sine_reg0   <= 36'sb111100011011001001001000101001001111;
        end
        16093: begin
            cosine_reg0 <= 36'sb11111110011010000101010101100001100;
            sine_reg0   <= 36'sb111100011011111011000101100011100010;
        end
        16094: begin
            cosine_reg0 <= 36'sb11111110011010110010000010101101111;
            sine_reg0   <= 36'sb111100011100101101000010100110101000;
        end
        16095: begin
            cosine_reg0 <= 36'sb11111110011011011110100110000110100;
            sine_reg0   <= 36'sb111100011101011110111111110010011110;
        end
        16096: begin
            cosine_reg0 <= 36'sb11111110011100001010111111101011010;
            sine_reg0   <= 36'sb111100011110010000111101000111000011;
        end
        16097: begin
            cosine_reg0 <= 36'sb11111110011100110111001111011100011;
            sine_reg0   <= 36'sb111100011111000010111010100100010101;
        end
        16098: begin
            cosine_reg0 <= 36'sb11111110011101100011010101011001100;
            sine_reg0   <= 36'sb111100011111110100111000001010010011;
        end
        16099: begin
            cosine_reg0 <= 36'sb11111110011110001111010001100010111;
            sine_reg0   <= 36'sb111100100000100110110101111000111001;
        end
        16100: begin
            cosine_reg0 <= 36'sb11111110011110111011000011111000010;
            sine_reg0   <= 36'sb111100100001011000110011110000000111;
        end
        16101: begin
            cosine_reg0 <= 36'sb11111110011111100110101100011001110;
            sine_reg0   <= 36'sb111100100010001010110001101111111001;
        end
        16102: begin
            cosine_reg0 <= 36'sb11111110100000010010001011000111011;
            sine_reg0   <= 36'sb111100100010111100101111111000010000;
        end
        16103: begin
            cosine_reg0 <= 36'sb11111110100000111101100000000001000;
            sine_reg0   <= 36'sb111100100011101110101110001001000111;
        end
        16104: begin
            cosine_reg0 <= 36'sb11111110100001101000101011000110101;
            sine_reg0   <= 36'sb111100100100100000101100100010011110;
        end
        16105: begin
            cosine_reg0 <= 36'sb11111110100010010011101100011000010;
            sine_reg0   <= 36'sb111100100101010010101011000100010011;
        end
        16106: begin
            cosine_reg0 <= 36'sb11111110100010111110100011110101111;
            sine_reg0   <= 36'sb111100100110000100101001101110100011;
        end
        16107: begin
            cosine_reg0 <= 36'sb11111110100011101001010001011111011;
            sine_reg0   <= 36'sb111100100110110110101000100001001101;
        end
        16108: begin
            cosine_reg0 <= 36'sb11111110100100010011110101010100110;
            sine_reg0   <= 36'sb111100100111101000100111011100001111;
        end
        16109: begin
            cosine_reg0 <= 36'sb11111110100100111110001111010110000;
            sine_reg0   <= 36'sb111100101000011010100110011111100111;
        end
        16110: begin
            cosine_reg0 <= 36'sb11111110100101101000011111100011001;
            sine_reg0   <= 36'sb111100101001001100100101101011010010;
        end
        16111: begin
            cosine_reg0 <= 36'sb11111110100110010010100101111100001;
            sine_reg0   <= 36'sb111100101001111110100100111111010000;
        end
        16112: begin
            cosine_reg0 <= 36'sb11111110100110111100100010100001000;
            sine_reg0   <= 36'sb111100101010110000100100011011011110;
        end
        16113: begin
            cosine_reg0 <= 36'sb11111110100111100110010101010001100;
            sine_reg0   <= 36'sb111100101011100010100011111111111010;
        end
        16114: begin
            cosine_reg0 <= 36'sb11111110101000001111111110001101110;
            sine_reg0   <= 36'sb111100101100010100100011101100100010;
        end
        16115: begin
            cosine_reg0 <= 36'sb11111110101000111001011101010101111;
            sine_reg0   <= 36'sb111100101101000110100011100001010100;
        end
        16116: begin
            cosine_reg0 <= 36'sb11111110101001100010110010101001101;
            sine_reg0   <= 36'sb111100101101111000100011011110001111;
        end
        16117: begin
            cosine_reg0 <= 36'sb11111110101010001011111110001001000;
            sine_reg0   <= 36'sb111100101110101010100011100011010000;
        end
        16118: begin
            cosine_reg0 <= 36'sb11111110101010110100111111110100001;
            sine_reg0   <= 36'sb111100101111011100100011110000010110;
        end
        16119: begin
            cosine_reg0 <= 36'sb11111110101011011101110111101010110;
            sine_reg0   <= 36'sb111100110000001110100100000101011110;
        end
        16120: begin
            cosine_reg0 <= 36'sb11111110101100000110100101101101001;
            sine_reg0   <= 36'sb111100110001000000100100100010100111;
        end
        16121: begin
            cosine_reg0 <= 36'sb11111110101100101111001001111011000;
            sine_reg0   <= 36'sb111100110001110010100101000111101111;
        end
        16122: begin
            cosine_reg0 <= 36'sb11111110101101010111100100010100100;
            sine_reg0   <= 36'sb111100110010100100100101110100110011;
        end
        16123: begin
            cosine_reg0 <= 36'sb11111110101101111111110100111001011;
            sine_reg0   <= 36'sb111100110011010110100110101001110010;
        end
        16124: begin
            cosine_reg0 <= 36'sb11111110101110100111111011101001111;
            sine_reg0   <= 36'sb111100110100001000100111100110101011;
        end
        16125: begin
            cosine_reg0 <= 36'sb11111110101111001111111000100101111;
            sine_reg0   <= 36'sb111100110100111010101000101011011010;
        end
        16126: begin
            cosine_reg0 <= 36'sb11111110101111110111101011101101010;
            sine_reg0   <= 36'sb111100110101101100101001110111111110;
        end
        16127: begin
            cosine_reg0 <= 36'sb11111110110000011111010101000000001;
            sine_reg0   <= 36'sb111100110110011110101011001100010110;
        end
        16128: begin
            cosine_reg0 <= 36'sb11111110110001000110110100011110011;
            sine_reg0   <= 36'sb111100110111010000101100101000011111;
        end
        16129: begin
            cosine_reg0 <= 36'sb11111110110001101110001010001000001;
            sine_reg0   <= 36'sb111100111000000010101110001100010111;
        end
        16130: begin
            cosine_reg0 <= 36'sb11111110110010010101010101111101001;
            sine_reg0   <= 36'sb111100111000110100101111110111111100;
        end
        16131: begin
            cosine_reg0 <= 36'sb11111110110010111100010111111101100;
            sine_reg0   <= 36'sb111100111001100110110001101011001101;
        end
        16132: begin
            cosine_reg0 <= 36'sb11111110110011100011010000001001001;
            sine_reg0   <= 36'sb111100111010011000110011100110001000;
        end
        16133: begin
            cosine_reg0 <= 36'sb11111110110100001001111110100000001;
            sine_reg0   <= 36'sb111100111011001010110101101000101010;
        end
        16134: begin
            cosine_reg0 <= 36'sb11111110110100110000100011000010011;
            sine_reg0   <= 36'sb111100111011111100110111110010110001;
        end
        16135: begin
            cosine_reg0 <= 36'sb11111110110101010110111101101111110;
            sine_reg0   <= 36'sb111100111100101110111010000100011101;
        end
        16136: begin
            cosine_reg0 <= 36'sb11111110110101111101001110101000100;
            sine_reg0   <= 36'sb111100111101100000111100011101101010;
        end
        16137: begin
            cosine_reg0 <= 36'sb11111110110110100011010101101100011;
            sine_reg0   <= 36'sb111100111110010010111110111110010111;
        end
        16138: begin
            cosine_reg0 <= 36'sb11111110110111001001010010111011100;
            sine_reg0   <= 36'sb111100111111000101000001100110100010;
        end
        16139: begin
            cosine_reg0 <= 36'sb11111110110111101111000110010101110;
            sine_reg0   <= 36'sb111100111111110111000100010110001001;
        end
        16140: begin
            cosine_reg0 <= 36'sb11111110111000010100101111111011001;
            sine_reg0   <= 36'sb111101000000101001000111001101001010;
        end
        16141: begin
            cosine_reg0 <= 36'sb11111110111000111010001111101011101;
            sine_reg0   <= 36'sb111101000001011011001010001011100100;
        end
        16142: begin
            cosine_reg0 <= 36'sb11111110111001011111100101100111001;
            sine_reg0   <= 36'sb111101000010001101001101010001010011;
        end
        16143: begin
            cosine_reg0 <= 36'sb11111110111010000100110001101101110;
            sine_reg0   <= 36'sb111101000010111111010000011110010111;
        end
        16144: begin
            cosine_reg0 <= 36'sb11111110111010101001110011111111011;
            sine_reg0   <= 36'sb111101000011110001010011110010101101;
        end
        16145: begin
            cosine_reg0 <= 36'sb11111110111011001110101100011100001;
            sine_reg0   <= 36'sb111101000100100011010111001110010100;
        end
        16146: begin
            cosine_reg0 <= 36'sb11111110111011110011011011000011110;
            sine_reg0   <= 36'sb111101000101010101011010110001001001;
        end
        16147: begin
            cosine_reg0 <= 36'sb11111110111100010111111111110110100;
            sine_reg0   <= 36'sb111101000110000111011110011011001011;
        end
        16148: begin
            cosine_reg0 <= 36'sb11111110111100111100011010110100001;
            sine_reg0   <= 36'sb111101000110111001100010001100010111;
        end
        16149: begin
            cosine_reg0 <= 36'sb11111110111101100000101011111100101;
            sine_reg0   <= 36'sb111101000111101011100110000100101100;
        end
        16150: begin
            cosine_reg0 <= 36'sb11111110111110000100110011010000001;
            sine_reg0   <= 36'sb111101001000011101101010000100001000;
        end
        16151: begin
            cosine_reg0 <= 36'sb11111110111110101000110000101110011;
            sine_reg0   <= 36'sb111101001001001111101110001010101001;
        end
        16152: begin
            cosine_reg0 <= 36'sb11111110111111001100100100010111101;
            sine_reg0   <= 36'sb111101001010000001110010011000001100;
        end
        16153: begin
            cosine_reg0 <= 36'sb11111110111111110000001110001011101;
            sine_reg0   <= 36'sb111101001010110011110110101100110001;
        end
        16154: begin
            cosine_reg0 <= 36'sb11111111000000010011101110001010100;
            sine_reg0   <= 36'sb111101001011100101111011001000010101;
        end
        16155: begin
            cosine_reg0 <= 36'sb11111111000000110111000100010100001;
            sine_reg0   <= 36'sb111101001100010111111111101010110101;
        end
        16156: begin
            cosine_reg0 <= 36'sb11111111000001011010010000101000101;
            sine_reg0   <= 36'sb111101001101001010000100010100010010;
        end
        16157: begin
            cosine_reg0 <= 36'sb11111111000001111101010011000111111;
            sine_reg0   <= 36'sb111101001101111100001001000100100111;
        end
        16158: begin
            cosine_reg0 <= 36'sb11111111000010100000001011110001110;
            sine_reg0   <= 36'sb111101001110101110001101111011110100;
        end
        16159: begin
            cosine_reg0 <= 36'sb11111111000011000010111010100110100;
            sine_reg0   <= 36'sb111101001111100000010010111001110110;
        end
        16160: begin
            cosine_reg0 <= 36'sb11111111000011100101011111100101110;
            sine_reg0   <= 36'sb111101010000010010010111111110101011;
        end
        16161: begin
            cosine_reg0 <= 36'sb11111111000100000111111010101111111;
            sine_reg0   <= 36'sb111101010001000100011101001010010010;
        end
        16162: begin
            cosine_reg0 <= 36'sb11111111000100101010001100000100100;
            sine_reg0   <= 36'sb111101010001110110100010011100101001;
        end
        16163: begin
            cosine_reg0 <= 36'sb11111111000101001100010011100011111;
            sine_reg0   <= 36'sb111101010010101000100111110101101110;
        end
        16164: begin
            cosine_reg0 <= 36'sb11111111000101101110010001001101110;
            sine_reg0   <= 36'sb111101010011011010101101010101011110;
        end
        16165: begin
            cosine_reg0 <= 36'sb11111111000110010000000101000010010;
            sine_reg0   <= 36'sb111101010100001100110010111011111000;
        end
        16166: begin
            cosine_reg0 <= 36'sb11111111000110110001101111000001011;
            sine_reg0   <= 36'sb111101010100111110111000101000111010;
        end
        16167: begin
            cosine_reg0 <= 36'sb11111111000111010011001111001011000;
            sine_reg0   <= 36'sb111101010101110000111110011100100010;
        end
        16168: begin
            cosine_reg0 <= 36'sb11111111000111110100100101011111001;
            sine_reg0   <= 36'sb111101010110100011000100010110101110;
        end
        16169: begin
            cosine_reg0 <= 36'sb11111111001000010101110001111101111;
            sine_reg0   <= 36'sb111101010111010101001010010111011100;
        end
        16170: begin
            cosine_reg0 <= 36'sb11111111001000110110110100100111000;
            sine_reg0   <= 36'sb111101011000000111010000011110101010;
        end
        16171: begin
            cosine_reg0 <= 36'sb11111111001001010111101101011010110;
            sine_reg0   <= 36'sb111101011000111001010110101100010110;
        end
        16172: begin
            cosine_reg0 <= 36'sb11111111001001111000011100011000110;
            sine_reg0   <= 36'sb111101011001101011011101000000011111;
        end
        16173: begin
            cosine_reg0 <= 36'sb11111111001010011001000001100001011;
            sine_reg0   <= 36'sb111101011010011101100011011011000010;
        end
        16174: begin
            cosine_reg0 <= 36'sb11111111001010111001011100110100010;
            sine_reg0   <= 36'sb111101011011001111101001111011111110;
        end
        16175: begin
            cosine_reg0 <= 36'sb11111111001011011001101110010001101;
            sine_reg0   <= 36'sb111101011100000001110000100011010000;
        end
        16176: begin
            cosine_reg0 <= 36'sb11111111001011111001110101111001011;
            sine_reg0   <= 36'sb111101011100110011110111010000110111;
        end
        16177: begin
            cosine_reg0 <= 36'sb11111111001100011001110011101011011;
            sine_reg0   <= 36'sb111101011101100101111110000100110000;
        end
        16178: begin
            cosine_reg0 <= 36'sb11111111001100111001100111100111110;
            sine_reg0   <= 36'sb111101011110011000000100111110111010;
        end
        16179: begin
            cosine_reg0 <= 36'sb11111111001101011001010001101110100;
            sine_reg0   <= 36'sb111101011111001010001011111111010011;
        end
        16180: begin
            cosine_reg0 <= 36'sb11111111001101111000110001111111100;
            sine_reg0   <= 36'sb111101011111111100010011000101111001;
        end
        16181: begin
            cosine_reg0 <= 36'sb11111111001110011000001000011010110;
            sine_reg0   <= 36'sb111101100000101110011010010010101010;
        end
        16182: begin
            cosine_reg0 <= 36'sb11111111001110110111010101000000011;
            sine_reg0   <= 36'sb111101100001100000100001100101100011;
        end
        16183: begin
            cosine_reg0 <= 36'sb11111111001111010110010111110000001;
            sine_reg0   <= 36'sb111101100010010010101000111110100100;
        end
        16184: begin
            cosine_reg0 <= 36'sb11111111001111110101010000101010001;
            sine_reg0   <= 36'sb111101100011000100110000011101101010;
        end
        16185: begin
            cosine_reg0 <= 36'sb11111111010000010011111111101110011;
            sine_reg0   <= 36'sb111101100011110110111000000010110011;
        end
        16186: begin
            cosine_reg0 <= 36'sb11111111010000110010100100111100110;
            sine_reg0   <= 36'sb111101100100101000111111101101111101;
        end
        16187: begin
            cosine_reg0 <= 36'sb11111111010001010001000000010101010;
            sine_reg0   <= 36'sb111101100101011011000111011111000111;
        end
        16188: begin
            cosine_reg0 <= 36'sb11111111010001101111010001111000000;
            sine_reg0   <= 36'sb111101100110001101001111010110001110;
        end
        16189: begin
            cosine_reg0 <= 36'sb11111111010010001101011001100100111;
            sine_reg0   <= 36'sb111101100110111111010111010011010001;
        end
        16190: begin
            cosine_reg0 <= 36'sb11111111010010101011010111011011110;
            sine_reg0   <= 36'sb111101100111110001011111010110001101;
        end
        16191: begin
            cosine_reg0 <= 36'sb11111111010011001001001011011100110;
            sine_reg0   <= 36'sb111101101000100011100111011111000000;
        end
        16192: begin
            cosine_reg0 <= 36'sb11111111010011100110110101100111111;
            sine_reg0   <= 36'sb111101101001010101101111101101101010;
        end
        16193: begin
            cosine_reg0 <= 36'sb11111111010100000100010101111101001;
            sine_reg0   <= 36'sb111101101010000111111000000010000111;
        end
        16194: begin
            cosine_reg0 <= 36'sb11111111010100100001101100011100010;
            sine_reg0   <= 36'sb111101101010111010000000011100010110;
        end
        16195: begin
            cosine_reg0 <= 36'sb11111111010100111110111001000101100;
            sine_reg0   <= 36'sb111101101011101100001000111100010100;
        end
        16196: begin
            cosine_reg0 <= 36'sb11111111010101011011111011111000110;
            sine_reg0   <= 36'sb111101101100011110010001100010000001;
        end
        16197: begin
            cosine_reg0 <= 36'sb11111111010101111000110100110110000;
            sine_reg0   <= 36'sb111101101101010000011010001101011010;
        end
        16198: begin
            cosine_reg0 <= 36'sb11111111010110010101100011111101001;
            sine_reg0   <= 36'sb111101101110000010100010111110011101;
        end
        16199: begin
            cosine_reg0 <= 36'sb11111111010110110010001001001110010;
            sine_reg0   <= 36'sb111101101110110100101011110101001000;
        end
        16200: begin
            cosine_reg0 <= 36'sb11111111010111001110100100101001011;
            sine_reg0   <= 36'sb111101101111100110110100110001011001;
        end
        16201: begin
            cosine_reg0 <= 36'sb11111111010111101010110110001110011;
            sine_reg0   <= 36'sb111101110000011000111101110011001110;
        end
        16202: begin
            cosine_reg0 <= 36'sb11111111011000000110111101111101010;
            sine_reg0   <= 36'sb111101110001001011000110111010100110;
        end
        16203: begin
            cosine_reg0 <= 36'sb11111111011000100010111011110110000;
            sine_reg0   <= 36'sb111101110001111101010000000111011110;
        end
        16204: begin
            cosine_reg0 <= 36'sb11111111011000111110101111111000101;
            sine_reg0   <= 36'sb111101110010101111011001011001110101;
        end
        16205: begin
            cosine_reg0 <= 36'sb11111111011001011010011010000101001;
            sine_reg0   <= 36'sb111101110011100001100010110001101000;
        end
        16206: begin
            cosine_reg0 <= 36'sb11111111011001110101111010011011100;
            sine_reg0   <= 36'sb111101110100010011101100001110110110;
        end
        16207: begin
            cosine_reg0 <= 36'sb11111111011010010001010000111011101;
            sine_reg0   <= 36'sb111101110101000101110101110001011100;
        end
        16208: begin
            cosine_reg0 <= 36'sb11111111011010101100011101100101101;
            sine_reg0   <= 36'sb111101110101110111111111011001011001;
        end
        16209: begin
            cosine_reg0 <= 36'sb11111111011011000111100000011001010;
            sine_reg0   <= 36'sb111101110110101010001001000110101011;
        end
        16210: begin
            cosine_reg0 <= 36'sb11111111011011100010011001010110110;
            sine_reg0   <= 36'sb111101110111011100010010111001010000;
        end
        16211: begin
            cosine_reg0 <= 36'sb11111111011011111101001000011110000;
            sine_reg0   <= 36'sb111101111000001110011100110001000110;
        end
        16212: begin
            cosine_reg0 <= 36'sb11111111011100010111101101101111000;
            sine_reg0   <= 36'sb111101111001000000100110101110001011;
        end
        16213: begin
            cosine_reg0 <= 36'sb11111111011100110010001001001001110;
            sine_reg0   <= 36'sb111101111001110010110000110000011101;
        end
        16214: begin
            cosine_reg0 <= 36'sb11111111011101001100011010101110001;
            sine_reg0   <= 36'sb111101111010100100111010110111111010;
        end
        16215: begin
            cosine_reg0 <= 36'sb11111111011101100110100010011100010;
            sine_reg0   <= 36'sb111101111011010111000101000100100000;
        end
        16216: begin
            cosine_reg0 <= 36'sb11111111011110000000100000010100000;
            sine_reg0   <= 36'sb111101111100001001001111010110001110;
        end
        16217: begin
            cosine_reg0 <= 36'sb11111111011110011010010100010101011;
            sine_reg0   <= 36'sb111101111100111011011001101101000001;
        end
        16218: begin
            cosine_reg0 <= 36'sb11111111011110110011111110100000011;
            sine_reg0   <= 36'sb111101111101101101100100001000110111;
        end
        16219: begin
            cosine_reg0 <= 36'sb11111111011111001101011110110101001;
            sine_reg0   <= 36'sb111101111110011111101110101001101111;
        end
        16220: begin
            cosine_reg0 <= 36'sb11111111011111100110110101010011011;
            sine_reg0   <= 36'sb111101111111010001111001001111100110;
        end
        16221: begin
            cosine_reg0 <= 36'sb11111111100000000000000001111011010;
            sine_reg0   <= 36'sb111110000000000100000011111010011011;
        end
        16222: begin
            cosine_reg0 <= 36'sb11111111100000011001000100101100110;
            sine_reg0   <= 36'sb111110000000110110001110101010001100;
        end
        16223: begin
            cosine_reg0 <= 36'sb11111111100000110001111101100111110;
            sine_reg0   <= 36'sb111110000001101000011001011110110110;
        end
        16224: begin
            cosine_reg0 <= 36'sb11111111100001001010101100101100011;
            sine_reg0   <= 36'sb111110000010011010100100011000011000;
        end
        16225: begin
            cosine_reg0 <= 36'sb11111111100001100011010001111010011;
            sine_reg0   <= 36'sb111110000011001100101111010110110000;
        end
        16226: begin
            cosine_reg0 <= 36'sb11111111100001111011101101010010000;
            sine_reg0   <= 36'sb111110000011111110111010011001111100;
        end
        16227: begin
            cosine_reg0 <= 36'sb11111111100010010011111110110011010;
            sine_reg0   <= 36'sb111110000100110001000101100001111010;
        end
        16228: begin
            cosine_reg0 <= 36'sb11111111100010101100000110011101111;
            sine_reg0   <= 36'sb111110000101100011010000101110101000;
        end
        16229: begin
            cosine_reg0 <= 36'sb11111111100011000100000100010001111;
            sine_reg0   <= 36'sb111110000110010101011100000000000100;
        end
        16230: begin
            cosine_reg0 <= 36'sb11111111100011011011111000001111100;
            sine_reg0   <= 36'sb111110000111000111100111010110001101;
        end
        16231: begin
            cosine_reg0 <= 36'sb11111111100011110011100010010110100;
            sine_reg0   <= 36'sb111110000111111001110010110000111111;
        end
        16232: begin
            cosine_reg0 <= 36'sb11111111100100001011000010100110111;
            sine_reg0   <= 36'sb111110001000101011111110010000011010;
        end
        16233: begin
            cosine_reg0 <= 36'sb11111111100100100010011001000000110;
            sine_reg0   <= 36'sb111110001001011110001001110100011011;
        end
        16234: begin
            cosine_reg0 <= 36'sb11111111100100111001100101100100000;
            sine_reg0   <= 36'sb111110001010010000010101011101000001;
        end
        16235: begin
            cosine_reg0 <= 36'sb11111111100101010000101000010000101;
            sine_reg0   <= 36'sb111110001011000010100001001010001001;
        end
        16236: begin
            cosine_reg0 <= 36'sb11111111100101100111100001000110110;
            sine_reg0   <= 36'sb111110001011110100101100111011110010;
        end
        16237: begin
            cosine_reg0 <= 36'sb11111111100101111110010000000110001;
            sine_reg0   <= 36'sb111110001100100110111000110001111010;
        end
        16238: begin
            cosine_reg0 <= 36'sb11111111100110010100110101001110111;
            sine_reg0   <= 36'sb111110001101011001000100101100011110;
        end
        16239: begin
            cosine_reg0 <= 36'sb11111111100110101011010000100000111;
            sine_reg0   <= 36'sb111110001110001011010000101011011101;
        end
        16240: begin
            cosine_reg0 <= 36'sb11111111100111000001100001111100010;
            sine_reg0   <= 36'sb111110001110111101011100101110110101;
        end
        16241: begin
            cosine_reg0 <= 36'sb11111111100111010111101001100001000;
            sine_reg0   <= 36'sb111110001111101111101000110110100100;
        end
        16242: begin
            cosine_reg0 <= 36'sb11111111100111101101100111001111000;
            sine_reg0   <= 36'sb111110010000100001110101000010101000;
        end
        16243: begin
            cosine_reg0 <= 36'sb11111111101000000011011011000110010;
            sine_reg0   <= 36'sb111110010001010100000001010010111110;
        end
        16244: begin
            cosine_reg0 <= 36'sb11111111101000011001000101000110111;
            sine_reg0   <= 36'sb111110010010000110001101100111100110;
        end
        16245: begin
            cosine_reg0 <= 36'sb11111111101000101110100101010000101;
            sine_reg0   <= 36'sb111110010010111000011010000000011110;
        end
        16246: begin
            cosine_reg0 <= 36'sb11111111101001000011111011100011101;
            sine_reg0   <= 36'sb111110010011101010100110011101100010;
        end
        16247: begin
            cosine_reg0 <= 36'sb11111111101001011001001000000000000;
            sine_reg0   <= 36'sb111110010100011100110010111110110010;
        end
        16248: begin
            cosine_reg0 <= 36'sb11111111101001101110001010100101011;
            sine_reg0   <= 36'sb111110010101001110111111100100001011;
        end
        16249: begin
            cosine_reg0 <= 36'sb11111111101010000011000011010100001;
            sine_reg0   <= 36'sb111110010110000001001100001101101011;
        end
        16250: begin
            cosine_reg0 <= 36'sb11111111101010010111110010001100000;
            sine_reg0   <= 36'sb111110010110110011011000111011010001;
        end
        16251: begin
            cosine_reg0 <= 36'sb11111111101010101100010111001101001;
            sine_reg0   <= 36'sb111110010111100101100101101100111011;
        end
        16252: begin
            cosine_reg0 <= 36'sb11111111101011000000110010010111011;
            sine_reg0   <= 36'sb111110011000010111110010100010100110;
        end
        16253: begin
            cosine_reg0 <= 36'sb11111111101011010101000011101010110;
            sine_reg0   <= 36'sb111110011001001001111111011100010001;
        end
        16254: begin
            cosine_reg0 <= 36'sb11111111101011101001001011000111010;
            sine_reg0   <= 36'sb111110011001111100001100011001111001;
        end
        16255: begin
            cosine_reg0 <= 36'sb11111111101011111101001000101100111;
            sine_reg0   <= 36'sb111110011010101110011001011011011110;
        end
        16256: begin
            cosine_reg0 <= 36'sb11111111101100010000111100011011101;
            sine_reg0   <= 36'sb111110011011100000100110100000111100;
        end
        16257: begin
            cosine_reg0 <= 36'sb11111111101100100100100110010011100;
            sine_reg0   <= 36'sb111110011100010010110011101010010010;
        end
        16258: begin
            cosine_reg0 <= 36'sb11111111101100111000000110010100100;
            sine_reg0   <= 36'sb111110011101000101000000110111011110;
        end
        16259: begin
            cosine_reg0 <= 36'sb11111111101101001011011100011110101;
            sine_reg0   <= 36'sb111110011101110111001110001000011111;
        end
        16260: begin
            cosine_reg0 <= 36'sb11111111101101011110101000110001110;
            sine_reg0   <= 36'sb111110011110101001011011011101010001;
        end
        16261: begin
            cosine_reg0 <= 36'sb11111111101101110001101011001101111;
            sine_reg0   <= 36'sb111110011111011011101000110101110100;
        end
        16262: begin
            cosine_reg0 <= 36'sb11111111101110000100100011110011001;
            sine_reg0   <= 36'sb111110100000001101110110010010000101;
        end
        16263: begin
            cosine_reg0 <= 36'sb11111111101110010111010010100001011;
            sine_reg0   <= 36'sb111110100001000000000011110010000010;
        end
        16264: begin
            cosine_reg0 <= 36'sb11111111101110101001110111011000110;
            sine_reg0   <= 36'sb111110100001110010010001010101101010;
        end
        16265: begin
            cosine_reg0 <= 36'sb11111111101110111100010010011001000;
            sine_reg0   <= 36'sb111110100010100100011110111100111010;
        end
        16266: begin
            cosine_reg0 <= 36'sb11111111101111001110100011100010011;
            sine_reg0   <= 36'sb111110100011010110101100100111110001;
        end
        16267: begin
            cosine_reg0 <= 36'sb11111111101111100000101010110100101;
            sine_reg0   <= 36'sb111110100100001000111010010110001100;
        end
        16268: begin
            cosine_reg0 <= 36'sb11111111101111110010101000010000000;
            sine_reg0   <= 36'sb111110100100111011001000001000001010;
        end
        16269: begin
            cosine_reg0 <= 36'sb11111111110000000100011011110100010;
            sine_reg0   <= 36'sb111110100101101101010101111101101001;
        end
        16270: begin
            cosine_reg0 <= 36'sb11111111110000010110000101100001100;
            sine_reg0   <= 36'sb111110100110011111100011110110100110;
        end
        16271: begin
            cosine_reg0 <= 36'sb11111111110000100111100101010111101;
            sine_reg0   <= 36'sb111110100111010001110001110011000001;
        end
        16272: begin
            cosine_reg0 <= 36'sb11111111110000111000111011010110110;
            sine_reg0   <= 36'sb111110101000000011111111110010110110;
        end
        16273: begin
            cosine_reg0 <= 36'sb11111111110001001010000111011110110;
            sine_reg0   <= 36'sb111110101000110110001101110110000100;
        end
        16274: begin
            cosine_reg0 <= 36'sb11111111110001011011001001101111110;
            sine_reg0   <= 36'sb111110101001101000011011111100101001;
        end
        16275: begin
            cosine_reg0 <= 36'sb11111111110001101100000010001001101;
            sine_reg0   <= 36'sb111110101010011010101010000110100100;
        end
        16276: begin
            cosine_reg0 <= 36'sb11111111110001111100110000101100011;
            sine_reg0   <= 36'sb111110101011001100111000010011110001;
        end
        16277: begin
            cosine_reg0 <= 36'sb11111111110010001101010101011000000;
            sine_reg0   <= 36'sb111110101011111111000110100100010000;
        end
        16278: begin
            cosine_reg0 <= 36'sb11111111110010011101110000001100100;
            sine_reg0   <= 36'sb111110101100110001010100110111111110;
        end
        16279: begin
            cosine_reg0 <= 36'sb11111111110010101110000001001001111;
            sine_reg0   <= 36'sb111110101101100011100011001110111001;
        end
        16280: begin
            cosine_reg0 <= 36'sb11111111110010111110001000010000001;
            sine_reg0   <= 36'sb111110101110010101110001101001000000;
        end
        16281: begin
            cosine_reg0 <= 36'sb11111111110011001110000101011111010;
            sine_reg0   <= 36'sb111110101111001000000000000110010000;
        end
        16282: begin
            cosine_reg0 <= 36'sb11111111110011011101111000110111001;
            sine_reg0   <= 36'sb111110101111111010001110100110101000;
        end
        16283: begin
            cosine_reg0 <= 36'sb11111111110011101101100010010111111;
            sine_reg0   <= 36'sb111110110000101100011101001010000110;
        end
        16284: begin
            cosine_reg0 <= 36'sb11111111110011111101000010000001100;
            sine_reg0   <= 36'sb111110110001011110101011110000100111;
        end
        16285: begin
            cosine_reg0 <= 36'sb11111111110100001100010111110011111;
            sine_reg0   <= 36'sb111110110010010000111010011010001010;
        end
        16286: begin
            cosine_reg0 <= 36'sb11111111110100011011100011101111001;
            sine_reg0   <= 36'sb111110110011000011001001000110101101;
        end
        16287: begin
            cosine_reg0 <= 36'sb11111111110100101010100101110011001;
            sine_reg0   <= 36'sb111110110011110101010111110110001101;
        end
        16288: begin
            cosine_reg0 <= 36'sb11111111110100111001011101111111111;
            sine_reg0   <= 36'sb111110110100100111100110101000101010;
        end
        16289: begin
            cosine_reg0 <= 36'sb11111111110101001000001100010101011;
            sine_reg0   <= 36'sb111110110101011001110101011110000000;
        end
        16290: begin
            cosine_reg0 <= 36'sb11111111110101010110110000110011101;
            sine_reg0   <= 36'sb111110110110001100000100010110001111;
        end
        16291: begin
            cosine_reg0 <= 36'sb11111111110101100101001011011010110;
            sine_reg0   <= 36'sb111110110110111110010011010001010011;
        end
        16292: begin
            cosine_reg0 <= 36'sb11111111110101110011011100001010100;
            sine_reg0   <= 36'sb111110110111110000100010001111001100;
        end
        16293: begin
            cosine_reg0 <= 36'sb11111111110110000001100011000011001;
            sine_reg0   <= 36'sb111110111000100010110001001111110111;
        end
        16294: begin
            cosine_reg0 <= 36'sb11111111110110001111100000000100011;
            sine_reg0   <= 36'sb111110111001010101000000010011010011;
        end
        16295: begin
            cosine_reg0 <= 36'sb11111111110110011101010011001110011;
            sine_reg0   <= 36'sb111110111010000111001111011001011101;
        end
        16296: begin
            cosine_reg0 <= 36'sb11111111110110101010111100100001000;
            sine_reg0   <= 36'sb111110111010111001011110100010010011;
        end
        16297: begin
            cosine_reg0 <= 36'sb11111111110110111000011011111100100;
            sine_reg0   <= 36'sb111110111011101011101101101101110100;
        end
        16298: begin
            cosine_reg0 <= 36'sb11111111110111000101110001100000101;
            sine_reg0   <= 36'sb111110111100011101111100111011111101;
        end
        16299: begin
            cosine_reg0 <= 36'sb11111111110111010010111101001101011;
            sine_reg0   <= 36'sb111110111101010000001100001100101101;
        end
        16300: begin
            cosine_reg0 <= 36'sb11111111110111011111111111000010111;
            sine_reg0   <= 36'sb111110111110000010011011100000000010;
        end
        16301: begin
            cosine_reg0 <= 36'sb11111111110111101100110111000001000;
            sine_reg0   <= 36'sb111110111110110100101010110101111001;
        end
        16302: begin
            cosine_reg0 <= 36'sb11111111110111111001100101000111111;
            sine_reg0   <= 36'sb111110111111100110111010001110010001;
        end
        16303: begin
            cosine_reg0 <= 36'sb11111111111000000110001001010111010;
            sine_reg0   <= 36'sb111111000000011001001001101001001000;
        end
        16304: begin
            cosine_reg0 <= 36'sb11111111111000010010100011101111011;
            sine_reg0   <= 36'sb111111000001001011011001000110011100;
        end
        16305: begin
            cosine_reg0 <= 36'sb11111111111000011110110100010000010;
            sine_reg0   <= 36'sb111111000001111101101000100110001011;
        end
        16306: begin
            cosine_reg0 <= 36'sb11111111111000101010111010111001101;
            sine_reg0   <= 36'sb111111000010101111111000001000010100;
        end
        16307: begin
            cosine_reg0 <= 36'sb11111111111000110110110111101011101;
            sine_reg0   <= 36'sb111111000011100010000111101100110011;
        end
        16308: begin
            cosine_reg0 <= 36'sb11111111111001000010101010100110010;
            sine_reg0   <= 36'sb111111000100010100010111010011100111;
        end
        16309: begin
            cosine_reg0 <= 36'sb11111111111001001110010011101001100;
            sine_reg0   <= 36'sb111111000101000110100110111100101111;
        end
        16310: begin
            cosine_reg0 <= 36'sb11111111111001011001110010110101011;
            sine_reg0   <= 36'sb111111000101111000110110101000001000;
        end
        16311: begin
            cosine_reg0 <= 36'sb11111111111001100101001000001001111;
            sine_reg0   <= 36'sb111111000110101011000110010101110000;
        end
        16312: begin
            cosine_reg0 <= 36'sb11111111111001110000010011100111000;
            sine_reg0   <= 36'sb111111000111011101010110000101100110;
        end
        16313: begin
            cosine_reg0 <= 36'sb11111111111001111011010101001100101;
            sine_reg0   <= 36'sb111111001000001111100101110111101000;
        end
        16314: begin
            cosine_reg0 <= 36'sb11111111111010000110001100111010111;
            sine_reg0   <= 36'sb111111001001000001110101101011110011;
        end
        16315: begin
            cosine_reg0 <= 36'sb11111111111010010000111010110001101;
            sine_reg0   <= 36'sb111111001001110100000101100010000101;
        end
        16316: begin
            cosine_reg0 <= 36'sb11111111111010011011011110110001000;
            sine_reg0   <= 36'sb111111001010100110010101011010011101;
        end
        16317: begin
            cosine_reg0 <= 36'sb11111111111010100101111000111001000;
            sine_reg0   <= 36'sb111111001011011000100101010100111001;
        end
        16318: begin
            cosine_reg0 <= 36'sb11111111111010110000001001001001011;
            sine_reg0   <= 36'sb111111001100001010110101010001010111;
        end
        16319: begin
            cosine_reg0 <= 36'sb11111111111010111010001111100010100;
            sine_reg0   <= 36'sb111111001100111101000101001111110101;
        end
        16320: begin
            cosine_reg0 <= 36'sb11111111111011000100001100000100000;
            sine_reg0   <= 36'sb111111001101101111010101010000010001;
        end
        16321: begin
            cosine_reg0 <= 36'sb11111111111011001101111110101110001;
            sine_reg0   <= 36'sb111111001110100001100101010010101000;
        end
        16322: begin
            cosine_reg0 <= 36'sb11111111111011010111100111100000110;
            sine_reg0   <= 36'sb111111001111010011110101010110111010;
        end
        16323: begin
            cosine_reg0 <= 36'sb11111111111011100001000110011011111;
            sine_reg0   <= 36'sb111111010000000110000101011101000100;
        end
        16324: begin
            cosine_reg0 <= 36'sb11111111111011101010011011011111101;
            sine_reg0   <= 36'sb111111010000111000010101100101000100;
        end
        16325: begin
            cosine_reg0 <= 36'sb11111111111011110011100110101011110;
            sine_reg0   <= 36'sb111111010001101010100101101110111001;
        end
        16326: begin
            cosine_reg0 <= 36'sb11111111111011111100101000000000100;
            sine_reg0   <= 36'sb111111010010011100110101111010011111;
        end
        16327: begin
            cosine_reg0 <= 36'sb11111111111100000101011111011101110;
            sine_reg0   <= 36'sb111111010011001111000110000111110111;
        end
        16328: begin
            cosine_reg0 <= 36'sb11111111111100001110001101000011011;
            sine_reg0   <= 36'sb111111010100000001010110010110111100;
        end
        16329: begin
            cosine_reg0 <= 36'sb11111111111100010110110000110001101;
            sine_reg0   <= 36'sb111111010100110011100110100111101110;
        end
        16330: begin
            cosine_reg0 <= 36'sb11111111111100011111001010101000010;
            sine_reg0   <= 36'sb111111010101100101110110111010001011;
        end
        16331: begin
            cosine_reg0 <= 36'sb11111111111100100111011010100111011;
            sine_reg0   <= 36'sb111111010110011000000111001110010000;
        end
        16332: begin
            cosine_reg0 <= 36'sb11111111111100101111100000101111000;
            sine_reg0   <= 36'sb111111010111001010010111100011111100;
        end
        16333: begin
            cosine_reg0 <= 36'sb11111111111100110111011100111111001;
            sine_reg0   <= 36'sb111111010111111100100111111011001101;
        end
        16334: begin
            cosine_reg0 <= 36'sb11111111111100111111001111010111110;
            sine_reg0   <= 36'sb111111011000101110111000010100000000;
        end
        16335: begin
            cosine_reg0 <= 36'sb11111111111101000110110111111000110;
            sine_reg0   <= 36'sb111111011001100001001000101110010101;
        end
        16336: begin
            cosine_reg0 <= 36'sb11111111111101001110010110100010010;
            sine_reg0   <= 36'sb111111011010010011011001001010001000;
        end
        16337: begin
            cosine_reg0 <= 36'sb11111111111101010101101011010100001;
            sine_reg0   <= 36'sb111111011011000101101001100111011001;
        end
        16338: begin
            cosine_reg0 <= 36'sb11111111111101011100110110001110100;
            sine_reg0   <= 36'sb111111011011110111111010000110000100;
        end
        16339: begin
            cosine_reg0 <= 36'sb11111111111101100011110111010001011;
            sine_reg0   <= 36'sb111111011100101010001010100110001001;
        end
        16340: begin
            cosine_reg0 <= 36'sb11111111111101101010101110011100101;
            sine_reg0   <= 36'sb111111011101011100011011000111100101;
        end
        16341: begin
            cosine_reg0 <= 36'sb11111111111101110001011011110000011;
            sine_reg0   <= 36'sb111111011110001110101011101010010110;
        end
        16342: begin
            cosine_reg0 <= 36'sb11111111111101110111111111001100100;
            sine_reg0   <= 36'sb111111011111000000111100001110011010;
        end
        16343: begin
            cosine_reg0 <= 36'sb11111111111101111110011000110001000;
            sine_reg0   <= 36'sb111111011111110011001100110011110000;
        end
        16344: begin
            cosine_reg0 <= 36'sb11111111111110000100101000011110000;
            sine_reg0   <= 36'sb111111100000100101011101011010010101;
        end
        16345: begin
            cosine_reg0 <= 36'sb11111111111110001010101110010011100;
            sine_reg0   <= 36'sb111111100001010111101110000010001000;
        end
        16346: begin
            cosine_reg0 <= 36'sb11111111111110010000101010010001010;
            sine_reg0   <= 36'sb111111100010001001111110101011000110;
        end
        16347: begin
            cosine_reg0 <= 36'sb11111111111110010110011100010111100;
            sine_reg0   <= 36'sb111111100010111100001111010101001110;
        end
        16348: begin
            cosine_reg0 <= 36'sb11111111111110011100000100100110001;
            sine_reg0   <= 36'sb111111100011101110100000000000011110;
        end
        16349: begin
            cosine_reg0 <= 36'sb11111111111110100001100010111101010;
            sine_reg0   <= 36'sb111111100100100000110000101100110100;
        end
        16350: begin
            cosine_reg0 <= 36'sb11111111111110100110110111011100101;
            sine_reg0   <= 36'sb111111100101010011000001011010001101;
        end
        16351: begin
            cosine_reg0 <= 36'sb11111111111110101100000010000100100;
            sine_reg0   <= 36'sb111111100110000101010010001000101000;
        end
        16352: begin
            cosine_reg0 <= 36'sb11111111111110110001000010110100110;
            sine_reg0   <= 36'sb111111100110110111100010111000000011;
        end
        16353: begin
            cosine_reg0 <= 36'sb11111111111110110101111001101101011;
            sine_reg0   <= 36'sb111111100111101001110011101000011100;
        end
        16354: begin
            cosine_reg0 <= 36'sb11111111111110111010100110101110011;
            sine_reg0   <= 36'sb111111101000011100000100011001110001;
        end
        16355: begin
            cosine_reg0 <= 36'sb11111111111110111111001001110111111;
            sine_reg0   <= 36'sb111111101001001110010101001100000001;
        end
        16356: begin
            cosine_reg0 <= 36'sb11111111111111000011100011001001101;
            sine_reg0   <= 36'sb111111101010000000100101111111001000;
        end
        16357: begin
            cosine_reg0 <= 36'sb11111111111111000111110010100011110;
            sine_reg0   <= 36'sb111111101010110010110110110011000110;
        end
        16358: begin
            cosine_reg0 <= 36'sb11111111111111001011111000000110011;
            sine_reg0   <= 36'sb111111101011100101000111100111111000;
        end
        16359: begin
            cosine_reg0 <= 36'sb11111111111111001111110011110001010;
            sine_reg0   <= 36'sb111111101100010111011000011101011101;
        end
        16360: begin
            cosine_reg0 <= 36'sb11111111111111010011100101100100101;
            sine_reg0   <= 36'sb111111101101001001101001010011110010;
        end
        16361: begin
            cosine_reg0 <= 36'sb11111111111111010111001101100000010;
            sine_reg0   <= 36'sb111111101101111011111010001010110101;
        end
        16362: begin
            cosine_reg0 <= 36'sb11111111111111011010101011100100011;
            sine_reg0   <= 36'sb111111101110101110001011000010100101;
        end
        16363: begin
            cosine_reg0 <= 36'sb11111111111111011101111111110000110;
            sine_reg0   <= 36'sb111111101111100000011011111011000000;
        end
        16364: begin
            cosine_reg0 <= 36'sb11111111111111100001001010000101100;
            sine_reg0   <= 36'sb111111110000010010101100110100000011;
        end
        16365: begin
            cosine_reg0 <= 36'sb11111111111111100100001010100010110;
            sine_reg0   <= 36'sb111111110001000100111101101101101101;
        end
        16366: begin
            cosine_reg0 <= 36'sb11111111111111100111000001001000010;
            sine_reg0   <= 36'sb111111110001110111001110100111111100;
        end
        16367: begin
            cosine_reg0 <= 36'sb11111111111111101001101101110110001;
            sine_reg0   <= 36'sb111111110010101001011111100010101110;
        end
        16368: begin
            cosine_reg0 <= 36'sb11111111111111101100010000101100011;
            sine_reg0   <= 36'sb111111110011011011110000011110000001;
        end
        16369: begin
            cosine_reg0 <= 36'sb11111111111111101110101001101010111;
            sine_reg0   <= 36'sb111111110100001110000001011001110011;
        end
        16370: begin
            cosine_reg0 <= 36'sb11111111111111110000111000110001111;
            sine_reg0   <= 36'sb111111110101000000010010010110000001;
        end
        16371: begin
            cosine_reg0 <= 36'sb11111111111111110010111110000001001;
            sine_reg0   <= 36'sb111111110101110010100011010010101011;
        end
        16372: begin
            cosine_reg0 <= 36'sb11111111111111110100111001011000111;
            sine_reg0   <= 36'sb111111110110100100110100001111101111;
        end
        16373: begin
            cosine_reg0 <= 36'sb11111111111111110110101010111000111;
            sine_reg0   <= 36'sb111111110111010111000101001101001001;
        end
        16374: begin
            cosine_reg0 <= 36'sb11111111111111111000010010100001001;
            sine_reg0   <= 36'sb111111111000001001010110001010111001;
        end
        16375: begin
            cosine_reg0 <= 36'sb11111111111111111001110000010001111;
            sine_reg0   <= 36'sb111111111000111011100111001000111100;
        end
        16376: begin
            cosine_reg0 <= 36'sb11111111111111111011000100001011000;
            sine_reg0   <= 36'sb111111111001101101111000000111010000;
        end
        16377: begin
            cosine_reg0 <= 36'sb11111111111111111100001110001100011;
            sine_reg0   <= 36'sb111111111010100000001001000101110100;
        end
        16378: begin
            cosine_reg0 <= 36'sb11111111111111111101001110010110001;
            sine_reg0   <= 36'sb111111111011010010011010000100100110;
        end
        16379: begin
            cosine_reg0 <= 36'sb11111111111111111110000100101000010;
            sine_reg0   <= 36'sb111111111100000100101011000011100011;
        end
        16380: begin
            cosine_reg0 <= 36'sb11111111111111111110110001000010101;
            sine_reg0   <= 36'sb111111111100110110111100000010101010;
        end
        16381: begin
            cosine_reg0 <= 36'sb11111111111111111111010011100101011;
            sine_reg0   <= 36'sb111111111101101001001101000001111001;
        end
        16382: begin
            cosine_reg0 <= 36'sb11111111111111111111101100010000101;
            sine_reg0   <= 36'sb111111111110011011011110000001001101;
        end
        default: begin
            cosine_reg0 <= 36'sb11111111111111111111111011000100000;
            sine_reg0   <= 36'sb111111111111001101101111000000100110;
        end
        endcase
        // Compute residual (value not obtained from table * 2*pi) // unsigned mult okay
        // residual_reg0 <= phase_accum[32-14-1:0] * 16'b1100100100001111;
    end
end

// Perform Correction
logic signed [WIDTH-1:0]                cosine_reg1;
logic signed [WIDTH-1:0]                sine_reg1;
// logic signed [RESIDUAL_WIDTH-1:0]       residual_reg1;

logic signed [WIDTH-1:0]                cosine_reg2;
logic signed [WIDTH-1:0]                sine_reg2;

always_ff @ (posedge i_clock) begin
    if (i_ready == 1'b1) begin
        // Pipeline Stage 1
        cosine_reg1 <= cosine_reg0;
        sine_reg1 <= sine_reg0;
        // residual_reg1 <= (residual_reg0[14+RESIDUAL_WIDTH-1:13] + 1'b1) >> 1;
        // Pipeline Stage 2
        cosine_reg2 <= cosine_reg1;
        sine_reg2 <= sine_reg1;

        // Pipeline Stage 3
        o_cosine_data <= cosine_reg2;
        o_sine_data <= sine_reg2;
    end
end

endmodule: dds

`default_nettype wire
