`timescale 10ps / 10ps

`default_nettype none

module skid #(
    parameter WIDTH = 16
) (
    input wire logic                i_clock,
    input wire logic                i_reset,
    // Upstream signaling
    input wire logic [WIDTH-1:0]    i_in_data,
    input wire logic                i_in_valid,
    output     logic                o_in_ready,
    // Downstream signaling
    output     logic [WIDTH-1:0]    o_out_data,
    output     logic                o_out_valid,
    input wire logic                i_out_ready);

// Reserve a place for out stored data, and a
// signal to indicate whether or not it is full.
logic [WIDTH-1:0] skid_reg;
logic             skid_reg_full;

// enum {
//     ST_START,
//     ST_IDLE,
//     ST_PASSTHRU,
//     ST_HALT
// } curr_state, next_state;
localparam ST_START    = 2'b00;
localparam ST_IDLE     = 2'b01;
localparam ST_PASSTHRU = 2'b10;
localparam ST_HALT     = 2'b11;
logic [1:0] curr_state;
logic [1:0] next_state;

// Combinatorial outputs of FSM
logic next_out_data;
logic next_out_valid;
logic next_skid_reg;
logic next_skid_reg_full;
logic next_in_ready;

// Register containing same data as output
logic [WIDTH-1:0] out_data_reg;

always @(posedge i_clock) begin
    if (i_reset == 1'b1) begin
        curr_state <= ST_START;
        o_out_data <= 0;
        o_out_valid <= 1'b0;
        out_data_reg <= 0;
        skid_reg <= 0;
        skid_reg_full <= 1'b0;
        o_in_ready <= 1'b0;
    end else begin
        // Update state machine
        curr_state <= next_state;
        // Update output interface signals
        o_out_data <= next_out_data;
        out_data_reg <= next_out_data;
        o_out_valid <= next_out_valid;
        // Update skid buffer signals
        skid_reg <= next_skid_reg;
        skid_reg_full <= next_skid_reg_full;
        // Update input interface signals
        o_in_ready <= next_in_ready;
    end
end

always @(*) begin
    case (curr_state)
    ST_IDLE: begin
        next_out_data = i_in_data;
        next_out_valid = i_in_valid;
        next_skid_reg = 0;
        next_skid_reg_full = 1'b0;
        next_in_ready = 1'b1;
        next_state = i_in_valid ? ST_PASSTHRU : ST_IDLE;
    end
    ST_PASSTHRU: begin
        next_out_data = i_out_ready ? i_in_data : out_data_reg;
        next_out_valid = ~(i_out_ready & (~i_in_valid));
        next_skid_reg = i_in_data;
        next_skid_reg_full = ~i_out_ready;
        next_in_ready = i_out_ready | ((~i_out_ready) & (~i_in_valid));
        case ({i_out_ready, i_in_valid})
        2'b11: next_state = ST_PASSTHRU;
        2'b10: next_state = ST_IDLE;
        2'b01: next_state = ST_HALT;
        2'b00: next_state = ST_PASSTHRU;
        default: $display("Error: Reached the unreachable state!");
        endcase
    end
    ST_HALT: begin
        next_out_data = i_out_ready ? skid_reg : out_data_reg;
        next_out_valid = 1'b1;
        next_skid_reg = skid_reg;
        next_skid_reg_full = ~i_out_ready;
        next_in_ready = i_out_ready;
        next_state = i_out_ready ? ST_PASSTHRU : ST_HALT;
    end
    default: begin
        next_out_data = 0;
        next_out_valid = 1'b0;
        next_skid_reg = 0;
        next_skid_reg_full = 1'b0;
        next_in_ready = 1'b1;
        next_state = ST_IDLE;
    end
    endcase
end

endmodule: skid

`default_nettype wire
