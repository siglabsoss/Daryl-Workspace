// Generated from template on 01/10/2017.
`timescale 1ps / 1ps

`default_nettype none

module sparse_mult_by_A #(
    parameter integer IN_WIDTH = 8,  // SHOULD BE A POWER OF 2
    parameter integer OUT_WIDTH = 96  // SHOULD BE A POWER OF 2
) (
    input  wire logic [IN_WIDTH-1:0]    i_input_data,
    input  wire logic                   i_input_valid,
    output      logic                   o_input_ready,
    output      logic [OUT_WIDTH-1:0]   o_output_data,
    output      logic                   o_output_valid,
    input  wire logic                   i_output_ready,
    input  wire logic                   i_clock,
    input  wire logic                   i_reset
);

localparam integer INPUT_LENGTH = 144;
localparam integer OUTPUT_LENGTH = 11;

// Track which buffers are full on current clock cycle
logic ping_is_full;
logic pong_is_full;

typedef enum {
    ST_INIT,
    ST_PING,
    ST_PONG,
    ST_WAIT_FOR_PING,
    ST_WAIT_FOR_PONG
} states_t;

states_t fillup_state;
states_t next_fillup_state;
states_t readout_state;
states_t next_readout_state;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        fillup_state <= ST_INIT;
        readout_state <= ST_INIT;
    end else begin
        fillup_state <= next_fillup_state;
        readout_state <= next_readout_state;
    end
end

logic [$clog2(INPUT_LENGTH)-1:0] input_count;
logic [$clog2(OUTPUT_LENGTH)-1:0] output_count;
always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        input_count <= '0;
        output_count <= '0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (input_count >= INPUT_LENGTH - 1) begin
                input_count <= '0;
            end else begin
                input_count <= input_count + 1;
            end
        end
        if ((o_output_valid & i_output_ready) == 1'b1) begin
            if (output_count >= OUTPUT_LENGTH - 1) begin
                output_count <= '0;
            end else begin
                output_count <= output_count + 1;
            end
        end

    end
end

// Used for the case structure in the next always block
logic [5:0] ping_pong_test;
logic       last_cycle_in;
logic       last_cycle_out;
// A transition to ST_PING or ST_PONG indicates that
// the bit accumulators should be reset to 1'b0...
logic       fillup_transition;
assign ping_pong_test = {
    last_cycle_in, last_cycle_out,
    i_input_valid, o_input_ready,
    o_output_valid, i_output_ready
};
always_ff @(posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_is_full <= 1'b0;
        pong_is_full <= 1'b0;
        fillup_transition <= 1'b0;
    end else begin
        // Calculate when we are on the last cycle of input
        if ((i_input_valid == 1'b1)
                && ((fillup_state == ST_PING)
                    || (fillup_state == ST_PONG))) begin
            last_cycle_in <= input_count == INPUT_LENGTH-2;
        end else begin
            last_cycle_in <= 1'b0;
        end
        // Calculate when we are on the last cycle of output
        if ((i_output_ready == 1'b1)
                && ((readout_state == ST_PING)
                    || (readout_state == ST_PONG))) begin
            last_cycle_out <= output_count == OUTPUT_LENGTH-2;
        end else begin
            last_cycle_out <= 1'b0;
        end
        // Incdicate when the ping and/or pong buffer is full to FSM
        case (ping_pong_test)
        6'b101100, 6'b101101, 6'b101110, 6'b101111, 6'b111100, 6'b111101, 6'b111110: begin
            if (fillup_state == ST_PING) begin
                ping_is_full <= 1'b1;
            end else begin
                pong_is_full <= 1'b1;
            end
        end
        6'b010011, 6'b010111, 6'b011011, 6'b011111, 6'b110011, 6'b110111, 6'b111011: begin
            if (readout_state == ST_PING) begin
                ping_is_full <= 1'b0;
            end else begin
                pong_is_full <= 1'b0;
            end
        end
        6'b111111:
            if (readout_state == ST_PING) begin
                ping_is_full <= 1'b0;
                pong_is_full <= 1'b1;
            end else begin
                ping_is_full <= 1'b1;
                pong_is_full <= 1'b0;
            end
        default: begin
            ping_is_full <= ping_is_full;
            pong_is_full <= pong_is_full;
        end
        endcase
        // Indicate a clock cycle when a transition occurs.
        if (((next_fillup_state == ST_PING) && (fillup_state != ST_PING))
                || ((next_fillup_state == ST_PONG) && (fillup_state != ST_PONG))) begin
            fillup_transition <= 1'b1;
        end else begin
            fillup_transition <= 1'b0;
        end
    end
end

always_comb begin
    case (fillup_state)
    ST_PING: begin
        if ((input_count == INPUT_LENGTH - 1)
                && (i_input_valid == 1'b1)) begin
            next_fillup_state = pong_is_full ? ST_WAIT_FOR_PONG : ST_PONG;
        end else begin
            next_fillup_state = ST_PING;
        end
        o_input_ready = 1'b1;
    end
    ST_PONG: begin
        if ((input_count == INPUT_LENGTH - 1)
                && (i_input_valid == 1'b1)) begin
            next_fillup_state = ping_is_full ? ST_WAIT_FOR_PING : ST_PING;
        end else begin
            next_fillup_state = ST_PONG;
        end
        o_input_ready = 1'b1;
    end
    ST_WAIT_FOR_PING: begin
        if (ping_is_full == 1'b0) begin
            next_fillup_state = ST_PING;
        end else begin
            next_fillup_state = ST_WAIT_FOR_PING;
        end
        o_input_ready = 1'b0;
    end
    ST_WAIT_FOR_PONG: begin
        if (pong_is_full == 1'b0) begin
            next_fillup_state = ST_PONG;
        end else begin
            next_fillup_state = ST_WAIT_FOR_PONG;
        end
        o_input_ready = 1'b0;
    end
    default: begin // ST_INIT
        next_fillup_state = ST_PING;
        o_input_ready = 1'b0;
    end
    endcase
end

always_comb begin
    case (readout_state)
    ST_PING: begin
        if ((output_count == OUTPUT_LENGTH - 1)
                && (i_output_ready == 1'b1)) begin
            next_readout_state = pong_is_full ? ST_PONG : ST_WAIT_FOR_PONG;
        end else begin
            next_readout_state = ST_PING;
        end
        case (output_count)
        0: o_output_data = {
            ping_storage_data_95,
            ping_storage_data_94,
            ping_storage_data_93,
            ping_storage_data_92,
            ping_storage_data_91,
            ping_storage_data_90,
            ping_storage_data_89,
            ping_storage_data_88,
            ping_storage_data_87,
            ping_storage_data_86,
            ping_storage_data_85,
            ping_storage_data_84,
            ping_storage_data_83,
            ping_storage_data_82,
            ping_storage_data_81,
            ping_storage_data_80,
            ping_storage_data_79,
            ping_storage_data_78,
            ping_storage_data_77,
            ping_storage_data_76,
            ping_storage_data_75,
            ping_storage_data_74,
            ping_storage_data_73,
            ping_storage_data_72,
            ping_storage_data_71,
            ping_storage_data_70,
            ping_storage_data_69,
            ping_storage_data_68,
            ping_storage_data_67,
            ping_storage_data_66,
            ping_storage_data_65,
            ping_storage_data_64,
            ping_storage_data_63,
            ping_storage_data_62,
            ping_storage_data_61,
            ping_storage_data_60,
            ping_storage_data_59,
            ping_storage_data_58,
            ping_storage_data_57,
            ping_storage_data_56,
            ping_storage_data_55,
            ping_storage_data_54,
            ping_storage_data_53,
            ping_storage_data_52,
            ping_storage_data_51,
            ping_storage_data_50,
            ping_storage_data_49,
            ping_storage_data_48,
            ping_storage_data_47,
            ping_storage_data_46,
            ping_storage_data_45,
            ping_storage_data_44,
            ping_storage_data_43,
            ping_storage_data_42,
            ping_storage_data_41,
            ping_storage_data_40,
            ping_storage_data_39,
            ping_storage_data_38,
            ping_storage_data_37,
            ping_storage_data_36,
            ping_storage_data_35,
            ping_storage_data_34,
            ping_storage_data_33,
            ping_storage_data_32,
            ping_storage_data_31,
            ping_storage_data_30,
            ping_storage_data_29,
            ping_storage_data_28,
            ping_storage_data_27,
            ping_storage_data_26,
            ping_storage_data_25,
            ping_storage_data_24,
            ping_storage_data_23,
            ping_storage_data_22,
            ping_storage_data_21,
            ping_storage_data_20,
            ping_storage_data_19,
            ping_storage_data_18,
            ping_storage_data_17,
            ping_storage_data_16,
            ping_storage_data_15,
            ping_storage_data_14,
            ping_storage_data_13,
            ping_storage_data_12,
            ping_storage_data_11,
            ping_storage_data_10,
            ping_storage_data_9,
            ping_storage_data_8,
            ping_storage_data_7,
            ping_storage_data_6,
            ping_storage_data_5,
            ping_storage_data_4,
            ping_storage_data_3,
            ping_storage_data_2,
            ping_storage_data_1,
            ping_storage_data_0
        };
        1: o_output_data = {
            ping_storage_data_191,
            ping_storage_data_190,
            ping_storage_data_189,
            ping_storage_data_188,
            ping_storage_data_187,
            ping_storage_data_186,
            ping_storage_data_185,
            ping_storage_data_184,
            ping_storage_data_183,
            ping_storage_data_182,
            ping_storage_data_181,
            ping_storage_data_180,
            ping_storage_data_179,
            ping_storage_data_178,
            ping_storage_data_177,
            ping_storage_data_176,
            ping_storage_data_175,
            ping_storage_data_174,
            ping_storage_data_173,
            ping_storage_data_172,
            ping_storage_data_171,
            ping_storage_data_170,
            ping_storage_data_169,
            ping_storage_data_168,
            ping_storage_data_167,
            ping_storage_data_166,
            ping_storage_data_165,
            ping_storage_data_164,
            ping_storage_data_163,
            ping_storage_data_162,
            ping_storage_data_161,
            ping_storage_data_160,
            ping_storage_data_159,
            ping_storage_data_158,
            ping_storage_data_157,
            ping_storage_data_156,
            ping_storage_data_155,
            ping_storage_data_154,
            ping_storage_data_153,
            ping_storage_data_152,
            ping_storage_data_151,
            ping_storage_data_150,
            ping_storage_data_149,
            ping_storage_data_148,
            ping_storage_data_147,
            ping_storage_data_146,
            ping_storage_data_145,
            ping_storage_data_144,
            ping_storage_data_143,
            ping_storage_data_142,
            ping_storage_data_141,
            ping_storage_data_140,
            ping_storage_data_139,
            ping_storage_data_138,
            ping_storage_data_137,
            ping_storage_data_136,
            ping_storage_data_135,
            ping_storage_data_134,
            ping_storage_data_133,
            ping_storage_data_132,
            ping_storage_data_131,
            ping_storage_data_130,
            ping_storage_data_129,
            ping_storage_data_128,
            ping_storage_data_127,
            ping_storage_data_126,
            ping_storage_data_125,
            ping_storage_data_124,
            ping_storage_data_123,
            ping_storage_data_122,
            ping_storage_data_121,
            ping_storage_data_120,
            ping_storage_data_119,
            ping_storage_data_118,
            ping_storage_data_117,
            ping_storage_data_116,
            ping_storage_data_115,
            ping_storage_data_114,
            ping_storage_data_113,
            ping_storage_data_112,
            ping_storage_data_111,
            ping_storage_data_110,
            ping_storage_data_109,
            ping_storage_data_108,
            ping_storage_data_107,
            ping_storage_data_106,
            ping_storage_data_105,
            ping_storage_data_104,
            ping_storage_data_103,
            ping_storage_data_102,
            ping_storage_data_101,
            ping_storage_data_100,
            ping_storage_data_99,
            ping_storage_data_98,
            ping_storage_data_97,
            ping_storage_data_96
        };
        2: o_output_data = {
            ping_storage_data_287,
            ping_storage_data_286,
            ping_storage_data_285,
            ping_storage_data_284,
            ping_storage_data_283,
            ping_storage_data_282,
            ping_storage_data_281,
            ping_storage_data_280,
            ping_storage_data_279,
            ping_storage_data_278,
            ping_storage_data_277,
            ping_storage_data_276,
            ping_storage_data_275,
            ping_storage_data_274,
            ping_storage_data_273,
            ping_storage_data_272,
            ping_storage_data_271,
            ping_storage_data_270,
            ping_storage_data_269,
            ping_storage_data_268,
            ping_storage_data_267,
            ping_storage_data_266,
            ping_storage_data_265,
            ping_storage_data_264,
            ping_storage_data_263,
            ping_storage_data_262,
            ping_storage_data_261,
            ping_storage_data_260,
            ping_storage_data_259,
            ping_storage_data_258,
            ping_storage_data_257,
            ping_storage_data_256,
            ping_storage_data_255,
            ping_storage_data_254,
            ping_storage_data_253,
            ping_storage_data_252,
            ping_storage_data_251,
            ping_storage_data_250,
            ping_storage_data_249,
            ping_storage_data_248,
            ping_storage_data_247,
            ping_storage_data_246,
            ping_storage_data_245,
            ping_storage_data_244,
            ping_storage_data_243,
            ping_storage_data_242,
            ping_storage_data_241,
            ping_storage_data_240,
            ping_storage_data_239,
            ping_storage_data_238,
            ping_storage_data_237,
            ping_storage_data_236,
            ping_storage_data_235,
            ping_storage_data_234,
            ping_storage_data_233,
            ping_storage_data_232,
            ping_storage_data_231,
            ping_storage_data_230,
            ping_storage_data_229,
            ping_storage_data_228,
            ping_storage_data_227,
            ping_storage_data_226,
            ping_storage_data_225,
            ping_storage_data_224,
            ping_storage_data_223,
            ping_storage_data_222,
            ping_storage_data_221,
            ping_storage_data_220,
            ping_storage_data_219,
            ping_storage_data_218,
            ping_storage_data_217,
            ping_storage_data_216,
            ping_storage_data_215,
            ping_storage_data_214,
            ping_storage_data_213,
            ping_storage_data_212,
            ping_storage_data_211,
            ping_storage_data_210,
            ping_storage_data_209,
            ping_storage_data_208,
            ping_storage_data_207,
            ping_storage_data_206,
            ping_storage_data_205,
            ping_storage_data_204,
            ping_storage_data_203,
            ping_storage_data_202,
            ping_storage_data_201,
            ping_storage_data_200,
            ping_storage_data_199,
            ping_storage_data_198,
            ping_storage_data_197,
            ping_storage_data_196,
            ping_storage_data_195,
            ping_storage_data_194,
            ping_storage_data_193,
            ping_storage_data_192
        };
        3: o_output_data = {
            ping_storage_data_383,
            ping_storage_data_382,
            ping_storage_data_381,
            ping_storage_data_380,
            ping_storage_data_379,
            ping_storage_data_378,
            ping_storage_data_377,
            ping_storage_data_376,
            ping_storage_data_375,
            ping_storage_data_374,
            ping_storage_data_373,
            ping_storage_data_372,
            ping_storage_data_371,
            ping_storage_data_370,
            ping_storage_data_369,
            ping_storage_data_368,
            ping_storage_data_367,
            ping_storage_data_366,
            ping_storage_data_365,
            ping_storage_data_364,
            ping_storage_data_363,
            ping_storage_data_362,
            ping_storage_data_361,
            ping_storage_data_360,
            ping_storage_data_359,
            ping_storage_data_358,
            ping_storage_data_357,
            ping_storage_data_356,
            ping_storage_data_355,
            ping_storage_data_354,
            ping_storage_data_353,
            ping_storage_data_352,
            ping_storage_data_351,
            ping_storage_data_350,
            ping_storage_data_349,
            ping_storage_data_348,
            ping_storage_data_347,
            ping_storage_data_346,
            ping_storage_data_345,
            ping_storage_data_344,
            ping_storage_data_343,
            ping_storage_data_342,
            ping_storage_data_341,
            ping_storage_data_340,
            ping_storage_data_339,
            ping_storage_data_338,
            ping_storage_data_337,
            ping_storage_data_336,
            ping_storage_data_335,
            ping_storage_data_334,
            ping_storage_data_333,
            ping_storage_data_332,
            ping_storage_data_331,
            ping_storage_data_330,
            ping_storage_data_329,
            ping_storage_data_328,
            ping_storage_data_327,
            ping_storage_data_326,
            ping_storage_data_325,
            ping_storage_data_324,
            ping_storage_data_323,
            ping_storage_data_322,
            ping_storage_data_321,
            ping_storage_data_320,
            ping_storage_data_319,
            ping_storage_data_318,
            ping_storage_data_317,
            ping_storage_data_316,
            ping_storage_data_315,
            ping_storage_data_314,
            ping_storage_data_313,
            ping_storage_data_312,
            ping_storage_data_311,
            ping_storage_data_310,
            ping_storage_data_309,
            ping_storage_data_308,
            ping_storage_data_307,
            ping_storage_data_306,
            ping_storage_data_305,
            ping_storage_data_304,
            ping_storage_data_303,
            ping_storage_data_302,
            ping_storage_data_301,
            ping_storage_data_300,
            ping_storage_data_299,
            ping_storage_data_298,
            ping_storage_data_297,
            ping_storage_data_296,
            ping_storage_data_295,
            ping_storage_data_294,
            ping_storage_data_293,
            ping_storage_data_292,
            ping_storage_data_291,
            ping_storage_data_290,
            ping_storage_data_289,
            ping_storage_data_288
        };
        4: o_output_data = {
            ping_storage_data_479,
            ping_storage_data_478,
            ping_storage_data_477,
            ping_storage_data_476,
            ping_storage_data_475,
            ping_storage_data_474,
            ping_storage_data_473,
            ping_storage_data_472,
            ping_storage_data_471,
            ping_storage_data_470,
            ping_storage_data_469,
            ping_storage_data_468,
            ping_storage_data_467,
            ping_storage_data_466,
            ping_storage_data_465,
            ping_storage_data_464,
            ping_storage_data_463,
            ping_storage_data_462,
            ping_storage_data_461,
            ping_storage_data_460,
            ping_storage_data_459,
            ping_storage_data_458,
            ping_storage_data_457,
            ping_storage_data_456,
            ping_storage_data_455,
            ping_storage_data_454,
            ping_storage_data_453,
            ping_storage_data_452,
            ping_storage_data_451,
            ping_storage_data_450,
            ping_storage_data_449,
            ping_storage_data_448,
            ping_storage_data_447,
            ping_storage_data_446,
            ping_storage_data_445,
            ping_storage_data_444,
            ping_storage_data_443,
            ping_storage_data_442,
            ping_storage_data_441,
            ping_storage_data_440,
            ping_storage_data_439,
            ping_storage_data_438,
            ping_storage_data_437,
            ping_storage_data_436,
            ping_storage_data_435,
            ping_storage_data_434,
            ping_storage_data_433,
            ping_storage_data_432,
            ping_storage_data_431,
            ping_storage_data_430,
            ping_storage_data_429,
            ping_storage_data_428,
            ping_storage_data_427,
            ping_storage_data_426,
            ping_storage_data_425,
            ping_storage_data_424,
            ping_storage_data_423,
            ping_storage_data_422,
            ping_storage_data_421,
            ping_storage_data_420,
            ping_storage_data_419,
            ping_storage_data_418,
            ping_storage_data_417,
            ping_storage_data_416,
            ping_storage_data_415,
            ping_storage_data_414,
            ping_storage_data_413,
            ping_storage_data_412,
            ping_storage_data_411,
            ping_storage_data_410,
            ping_storage_data_409,
            ping_storage_data_408,
            ping_storage_data_407,
            ping_storage_data_406,
            ping_storage_data_405,
            ping_storage_data_404,
            ping_storage_data_403,
            ping_storage_data_402,
            ping_storage_data_401,
            ping_storage_data_400,
            ping_storage_data_399,
            ping_storage_data_398,
            ping_storage_data_397,
            ping_storage_data_396,
            ping_storage_data_395,
            ping_storage_data_394,
            ping_storage_data_393,
            ping_storage_data_392,
            ping_storage_data_391,
            ping_storage_data_390,
            ping_storage_data_389,
            ping_storage_data_388,
            ping_storage_data_387,
            ping_storage_data_386,
            ping_storage_data_385,
            ping_storage_data_384
        };
        5: o_output_data = {
            ping_storage_data_575,
            ping_storage_data_574,
            ping_storage_data_573,
            ping_storage_data_572,
            ping_storage_data_571,
            ping_storage_data_570,
            ping_storage_data_569,
            ping_storage_data_568,
            ping_storage_data_567,
            ping_storage_data_566,
            ping_storage_data_565,
            ping_storage_data_564,
            ping_storage_data_563,
            ping_storage_data_562,
            ping_storage_data_561,
            ping_storage_data_560,
            ping_storage_data_559,
            ping_storage_data_558,
            ping_storage_data_557,
            ping_storage_data_556,
            ping_storage_data_555,
            ping_storage_data_554,
            ping_storage_data_553,
            ping_storage_data_552,
            ping_storage_data_551,
            ping_storage_data_550,
            ping_storage_data_549,
            ping_storage_data_548,
            ping_storage_data_547,
            ping_storage_data_546,
            ping_storage_data_545,
            ping_storage_data_544,
            ping_storage_data_543,
            ping_storage_data_542,
            ping_storage_data_541,
            ping_storage_data_540,
            ping_storage_data_539,
            ping_storage_data_538,
            ping_storage_data_537,
            ping_storage_data_536,
            ping_storage_data_535,
            ping_storage_data_534,
            ping_storage_data_533,
            ping_storage_data_532,
            ping_storage_data_531,
            ping_storage_data_530,
            ping_storage_data_529,
            ping_storage_data_528,
            ping_storage_data_527,
            ping_storage_data_526,
            ping_storage_data_525,
            ping_storage_data_524,
            ping_storage_data_523,
            ping_storage_data_522,
            ping_storage_data_521,
            ping_storage_data_520,
            ping_storage_data_519,
            ping_storage_data_518,
            ping_storage_data_517,
            ping_storage_data_516,
            ping_storage_data_515,
            ping_storage_data_514,
            ping_storage_data_513,
            ping_storage_data_512,
            ping_storage_data_511,
            ping_storage_data_510,
            ping_storage_data_509,
            ping_storage_data_508,
            ping_storage_data_507,
            ping_storage_data_506,
            ping_storage_data_505,
            ping_storage_data_504,
            ping_storage_data_503,
            ping_storage_data_502,
            ping_storage_data_501,
            ping_storage_data_500,
            ping_storage_data_499,
            ping_storage_data_498,
            ping_storage_data_497,
            ping_storage_data_496,
            ping_storage_data_495,
            ping_storage_data_494,
            ping_storage_data_493,
            ping_storage_data_492,
            ping_storage_data_491,
            ping_storage_data_490,
            ping_storage_data_489,
            ping_storage_data_488,
            ping_storage_data_487,
            ping_storage_data_486,
            ping_storage_data_485,
            ping_storage_data_484,
            ping_storage_data_483,
            ping_storage_data_482,
            ping_storage_data_481,
            ping_storage_data_480
        };
        6: o_output_data = {
            ping_storage_data_671,
            ping_storage_data_670,
            ping_storage_data_669,
            ping_storage_data_668,
            ping_storage_data_667,
            ping_storage_data_666,
            ping_storage_data_665,
            ping_storage_data_664,
            ping_storage_data_663,
            ping_storage_data_662,
            ping_storage_data_661,
            ping_storage_data_660,
            ping_storage_data_659,
            ping_storage_data_658,
            ping_storage_data_657,
            ping_storage_data_656,
            ping_storage_data_655,
            ping_storage_data_654,
            ping_storage_data_653,
            ping_storage_data_652,
            ping_storage_data_651,
            ping_storage_data_650,
            ping_storage_data_649,
            ping_storage_data_648,
            ping_storage_data_647,
            ping_storage_data_646,
            ping_storage_data_645,
            ping_storage_data_644,
            ping_storage_data_643,
            ping_storage_data_642,
            ping_storage_data_641,
            ping_storage_data_640,
            ping_storage_data_639,
            ping_storage_data_638,
            ping_storage_data_637,
            ping_storage_data_636,
            ping_storage_data_635,
            ping_storage_data_634,
            ping_storage_data_633,
            ping_storage_data_632,
            ping_storage_data_631,
            ping_storage_data_630,
            ping_storage_data_629,
            ping_storage_data_628,
            ping_storage_data_627,
            ping_storage_data_626,
            ping_storage_data_625,
            ping_storage_data_624,
            ping_storage_data_623,
            ping_storage_data_622,
            ping_storage_data_621,
            ping_storage_data_620,
            ping_storage_data_619,
            ping_storage_data_618,
            ping_storage_data_617,
            ping_storage_data_616,
            ping_storage_data_615,
            ping_storage_data_614,
            ping_storage_data_613,
            ping_storage_data_612,
            ping_storage_data_611,
            ping_storage_data_610,
            ping_storage_data_609,
            ping_storage_data_608,
            ping_storage_data_607,
            ping_storage_data_606,
            ping_storage_data_605,
            ping_storage_data_604,
            ping_storage_data_603,
            ping_storage_data_602,
            ping_storage_data_601,
            ping_storage_data_600,
            ping_storage_data_599,
            ping_storage_data_598,
            ping_storage_data_597,
            ping_storage_data_596,
            ping_storage_data_595,
            ping_storage_data_594,
            ping_storage_data_593,
            ping_storage_data_592,
            ping_storage_data_591,
            ping_storage_data_590,
            ping_storage_data_589,
            ping_storage_data_588,
            ping_storage_data_587,
            ping_storage_data_586,
            ping_storage_data_585,
            ping_storage_data_584,
            ping_storage_data_583,
            ping_storage_data_582,
            ping_storage_data_581,
            ping_storage_data_580,
            ping_storage_data_579,
            ping_storage_data_578,
            ping_storage_data_577,
            ping_storage_data_576
        };
        7: o_output_data = {
            ping_storage_data_767,
            ping_storage_data_766,
            ping_storage_data_765,
            ping_storage_data_764,
            ping_storage_data_763,
            ping_storage_data_762,
            ping_storage_data_761,
            ping_storage_data_760,
            ping_storage_data_759,
            ping_storage_data_758,
            ping_storage_data_757,
            ping_storage_data_756,
            ping_storage_data_755,
            ping_storage_data_754,
            ping_storage_data_753,
            ping_storage_data_752,
            ping_storage_data_751,
            ping_storage_data_750,
            ping_storage_data_749,
            ping_storage_data_748,
            ping_storage_data_747,
            ping_storage_data_746,
            ping_storage_data_745,
            ping_storage_data_744,
            ping_storage_data_743,
            ping_storage_data_742,
            ping_storage_data_741,
            ping_storage_data_740,
            ping_storage_data_739,
            ping_storage_data_738,
            ping_storage_data_737,
            ping_storage_data_736,
            ping_storage_data_735,
            ping_storage_data_734,
            ping_storage_data_733,
            ping_storage_data_732,
            ping_storage_data_731,
            ping_storage_data_730,
            ping_storage_data_729,
            ping_storage_data_728,
            ping_storage_data_727,
            ping_storage_data_726,
            ping_storage_data_725,
            ping_storage_data_724,
            ping_storage_data_723,
            ping_storage_data_722,
            ping_storage_data_721,
            ping_storage_data_720,
            ping_storage_data_719,
            ping_storage_data_718,
            ping_storage_data_717,
            ping_storage_data_716,
            ping_storage_data_715,
            ping_storage_data_714,
            ping_storage_data_713,
            ping_storage_data_712,
            ping_storage_data_711,
            ping_storage_data_710,
            ping_storage_data_709,
            ping_storage_data_708,
            ping_storage_data_707,
            ping_storage_data_706,
            ping_storage_data_705,
            ping_storage_data_704,
            ping_storage_data_703,
            ping_storage_data_702,
            ping_storage_data_701,
            ping_storage_data_700,
            ping_storage_data_699,
            ping_storage_data_698,
            ping_storage_data_697,
            ping_storage_data_696,
            ping_storage_data_695,
            ping_storage_data_694,
            ping_storage_data_693,
            ping_storage_data_692,
            ping_storage_data_691,
            ping_storage_data_690,
            ping_storage_data_689,
            ping_storage_data_688,
            ping_storage_data_687,
            ping_storage_data_686,
            ping_storage_data_685,
            ping_storage_data_684,
            ping_storage_data_683,
            ping_storage_data_682,
            ping_storage_data_681,
            ping_storage_data_680,
            ping_storage_data_679,
            ping_storage_data_678,
            ping_storage_data_677,
            ping_storage_data_676,
            ping_storage_data_675,
            ping_storage_data_674,
            ping_storage_data_673,
            ping_storage_data_672
        };
        8: o_output_data = {
            ping_storage_data_863,
            ping_storage_data_862,
            ping_storage_data_861,
            ping_storage_data_860,
            ping_storage_data_859,
            ping_storage_data_858,
            ping_storage_data_857,
            ping_storage_data_856,
            ping_storage_data_855,
            ping_storage_data_854,
            ping_storage_data_853,
            ping_storage_data_852,
            ping_storage_data_851,
            ping_storage_data_850,
            ping_storage_data_849,
            ping_storage_data_848,
            ping_storage_data_847,
            ping_storage_data_846,
            ping_storage_data_845,
            ping_storage_data_844,
            ping_storage_data_843,
            ping_storage_data_842,
            ping_storage_data_841,
            ping_storage_data_840,
            ping_storage_data_839,
            ping_storage_data_838,
            ping_storage_data_837,
            ping_storage_data_836,
            ping_storage_data_835,
            ping_storage_data_834,
            ping_storage_data_833,
            ping_storage_data_832,
            ping_storage_data_831,
            ping_storage_data_830,
            ping_storage_data_829,
            ping_storage_data_828,
            ping_storage_data_827,
            ping_storage_data_826,
            ping_storage_data_825,
            ping_storage_data_824,
            ping_storage_data_823,
            ping_storage_data_822,
            ping_storage_data_821,
            ping_storage_data_820,
            ping_storage_data_819,
            ping_storage_data_818,
            ping_storage_data_817,
            ping_storage_data_816,
            ping_storage_data_815,
            ping_storage_data_814,
            ping_storage_data_813,
            ping_storage_data_812,
            ping_storage_data_811,
            ping_storage_data_810,
            ping_storage_data_809,
            ping_storage_data_808,
            ping_storage_data_807,
            ping_storage_data_806,
            ping_storage_data_805,
            ping_storage_data_804,
            ping_storage_data_803,
            ping_storage_data_802,
            ping_storage_data_801,
            ping_storage_data_800,
            ping_storage_data_799,
            ping_storage_data_798,
            ping_storage_data_797,
            ping_storage_data_796,
            ping_storage_data_795,
            ping_storage_data_794,
            ping_storage_data_793,
            ping_storage_data_792,
            ping_storage_data_791,
            ping_storage_data_790,
            ping_storage_data_789,
            ping_storage_data_788,
            ping_storage_data_787,
            ping_storage_data_786,
            ping_storage_data_785,
            ping_storage_data_784,
            ping_storage_data_783,
            ping_storage_data_782,
            ping_storage_data_781,
            ping_storage_data_780,
            ping_storage_data_779,
            ping_storage_data_778,
            ping_storage_data_777,
            ping_storage_data_776,
            ping_storage_data_775,
            ping_storage_data_774,
            ping_storage_data_773,
            ping_storage_data_772,
            ping_storage_data_771,
            ping_storage_data_770,
            ping_storage_data_769,
            ping_storage_data_768
        };
        9: o_output_data = {
            ping_storage_data_959,
            ping_storage_data_958,
            ping_storage_data_957,
            ping_storage_data_956,
            ping_storage_data_955,
            ping_storage_data_954,
            ping_storage_data_953,
            ping_storage_data_952,
            ping_storage_data_951,
            ping_storage_data_950,
            ping_storage_data_949,
            ping_storage_data_948,
            ping_storage_data_947,
            ping_storage_data_946,
            ping_storage_data_945,
            ping_storage_data_944,
            ping_storage_data_943,
            ping_storage_data_942,
            ping_storage_data_941,
            ping_storage_data_940,
            ping_storage_data_939,
            ping_storage_data_938,
            ping_storage_data_937,
            ping_storage_data_936,
            ping_storage_data_935,
            ping_storage_data_934,
            ping_storage_data_933,
            ping_storage_data_932,
            ping_storage_data_931,
            ping_storage_data_930,
            ping_storage_data_929,
            ping_storage_data_928,
            ping_storage_data_927,
            ping_storage_data_926,
            ping_storage_data_925,
            ping_storage_data_924,
            ping_storage_data_923,
            ping_storage_data_922,
            ping_storage_data_921,
            ping_storage_data_920,
            ping_storage_data_919,
            ping_storage_data_918,
            ping_storage_data_917,
            ping_storage_data_916,
            ping_storage_data_915,
            ping_storage_data_914,
            ping_storage_data_913,
            ping_storage_data_912,
            ping_storage_data_911,
            ping_storage_data_910,
            ping_storage_data_909,
            ping_storage_data_908,
            ping_storage_data_907,
            ping_storage_data_906,
            ping_storage_data_905,
            ping_storage_data_904,
            ping_storage_data_903,
            ping_storage_data_902,
            ping_storage_data_901,
            ping_storage_data_900,
            ping_storage_data_899,
            ping_storage_data_898,
            ping_storage_data_897,
            ping_storage_data_896,
            ping_storage_data_895,
            ping_storage_data_894,
            ping_storage_data_893,
            ping_storage_data_892,
            ping_storage_data_891,
            ping_storage_data_890,
            ping_storage_data_889,
            ping_storage_data_888,
            ping_storage_data_887,
            ping_storage_data_886,
            ping_storage_data_885,
            ping_storage_data_884,
            ping_storage_data_883,
            ping_storage_data_882,
            ping_storage_data_881,
            ping_storage_data_880,
            ping_storage_data_879,
            ping_storage_data_878,
            ping_storage_data_877,
            ping_storage_data_876,
            ping_storage_data_875,
            ping_storage_data_874,
            ping_storage_data_873,
            ping_storage_data_872,
            ping_storage_data_871,
            ping_storage_data_870,
            ping_storage_data_869,
            ping_storage_data_868,
            ping_storage_data_867,
            ping_storage_data_866,
            ping_storage_data_865,
            ping_storage_data_864
        };
        default: o_output_data = {
            ping_storage_data_1055,
            ping_storage_data_1054,
            ping_storage_data_1053,
            ping_storage_data_1052,
            ping_storage_data_1051,
            ping_storage_data_1050,
            ping_storage_data_1049,
            ping_storage_data_1048,
            ping_storage_data_1047,
            ping_storage_data_1046,
            ping_storage_data_1045,
            ping_storage_data_1044,
            ping_storage_data_1043,
            ping_storage_data_1042,
            ping_storage_data_1041,
            ping_storage_data_1040,
            ping_storage_data_1039,
            ping_storage_data_1038,
            ping_storage_data_1037,
            ping_storage_data_1036,
            ping_storage_data_1035,
            ping_storage_data_1034,
            ping_storage_data_1033,
            ping_storage_data_1032,
            ping_storage_data_1031,
            ping_storage_data_1030,
            ping_storage_data_1029,
            ping_storage_data_1028,
            ping_storage_data_1027,
            ping_storage_data_1026,
            ping_storage_data_1025,
            ping_storage_data_1024,
            ping_storage_data_1023,
            ping_storage_data_1022,
            ping_storage_data_1021,
            ping_storage_data_1020,
            ping_storage_data_1019,
            ping_storage_data_1018,
            ping_storage_data_1017,
            ping_storage_data_1016,
            ping_storage_data_1015,
            ping_storage_data_1014,
            ping_storage_data_1013,
            ping_storage_data_1012,
            ping_storage_data_1011,
            ping_storage_data_1010,
            ping_storage_data_1009,
            ping_storage_data_1008,
            ping_storage_data_1007,
            ping_storage_data_1006,
            ping_storage_data_1005,
            ping_storage_data_1004,
            ping_storage_data_1003,
            ping_storage_data_1002,
            ping_storage_data_1001,
            ping_storage_data_1000,
            ping_storage_data_999,
            ping_storage_data_998,
            ping_storage_data_997,
            ping_storage_data_996,
            ping_storage_data_995,
            ping_storage_data_994,
            ping_storage_data_993,
            ping_storage_data_992,
            ping_storage_data_991,
            ping_storage_data_990,
            ping_storage_data_989,
            ping_storage_data_988,
            ping_storage_data_987,
            ping_storage_data_986,
            ping_storage_data_985,
            ping_storage_data_984,
            ping_storage_data_983,
            ping_storage_data_982,
            ping_storage_data_981,
            ping_storage_data_980,
            ping_storage_data_979,
            ping_storage_data_978,
            ping_storage_data_977,
            ping_storage_data_976,
            ping_storage_data_975,
            ping_storage_data_974,
            ping_storage_data_973,
            ping_storage_data_972,
            ping_storage_data_971,
            ping_storage_data_970,
            ping_storage_data_969,
            ping_storage_data_968,
            ping_storage_data_967,
            ping_storage_data_966,
            ping_storage_data_965,
            ping_storage_data_964,
            ping_storage_data_963,
            ping_storage_data_962,
            ping_storage_data_961,
            ping_storage_data_960
        };
        endcase
        o_output_valid = 1'b1;
    end
    ST_PONG: begin
        if ((output_count == OUTPUT_LENGTH - 1)
                && (i_output_ready == 1'b1)) begin
            next_readout_state = ping_is_full ? ST_PING : ST_WAIT_FOR_PING;
        end else begin
            next_readout_state = ST_PONG;
        end
        case (output_count)
        0: o_output_data = {
            pong_storage_data_95,
            pong_storage_data_94,
            pong_storage_data_93,
            pong_storage_data_92,
            pong_storage_data_91,
            pong_storage_data_90,
            pong_storage_data_89,
            pong_storage_data_88,
            pong_storage_data_87,
            pong_storage_data_86,
            pong_storage_data_85,
            pong_storage_data_84,
            pong_storage_data_83,
            pong_storage_data_82,
            pong_storage_data_81,
            pong_storage_data_80,
            pong_storage_data_79,
            pong_storage_data_78,
            pong_storage_data_77,
            pong_storage_data_76,
            pong_storage_data_75,
            pong_storage_data_74,
            pong_storage_data_73,
            pong_storage_data_72,
            pong_storage_data_71,
            pong_storage_data_70,
            pong_storage_data_69,
            pong_storage_data_68,
            pong_storage_data_67,
            pong_storage_data_66,
            pong_storage_data_65,
            pong_storage_data_64,
            pong_storage_data_63,
            pong_storage_data_62,
            pong_storage_data_61,
            pong_storage_data_60,
            pong_storage_data_59,
            pong_storage_data_58,
            pong_storage_data_57,
            pong_storage_data_56,
            pong_storage_data_55,
            pong_storage_data_54,
            pong_storage_data_53,
            pong_storage_data_52,
            pong_storage_data_51,
            pong_storage_data_50,
            pong_storage_data_49,
            pong_storage_data_48,
            pong_storage_data_47,
            pong_storage_data_46,
            pong_storage_data_45,
            pong_storage_data_44,
            pong_storage_data_43,
            pong_storage_data_42,
            pong_storage_data_41,
            pong_storage_data_40,
            pong_storage_data_39,
            pong_storage_data_38,
            pong_storage_data_37,
            pong_storage_data_36,
            pong_storage_data_35,
            pong_storage_data_34,
            pong_storage_data_33,
            pong_storage_data_32,
            pong_storage_data_31,
            pong_storage_data_30,
            pong_storage_data_29,
            pong_storage_data_28,
            pong_storage_data_27,
            pong_storage_data_26,
            pong_storage_data_25,
            pong_storage_data_24,
            pong_storage_data_23,
            pong_storage_data_22,
            pong_storage_data_21,
            pong_storage_data_20,
            pong_storage_data_19,
            pong_storage_data_18,
            pong_storage_data_17,
            pong_storage_data_16,
            pong_storage_data_15,
            pong_storage_data_14,
            pong_storage_data_13,
            pong_storage_data_12,
            pong_storage_data_11,
            pong_storage_data_10,
            pong_storage_data_9,
            pong_storage_data_8,
            pong_storage_data_7,
            pong_storage_data_6,
            pong_storage_data_5,
            pong_storage_data_4,
            pong_storage_data_3,
            pong_storage_data_2,
            pong_storage_data_1,
            pong_storage_data_0
        };
        1: o_output_data = {
            pong_storage_data_191,
            pong_storage_data_190,
            pong_storage_data_189,
            pong_storage_data_188,
            pong_storage_data_187,
            pong_storage_data_186,
            pong_storage_data_185,
            pong_storage_data_184,
            pong_storage_data_183,
            pong_storage_data_182,
            pong_storage_data_181,
            pong_storage_data_180,
            pong_storage_data_179,
            pong_storage_data_178,
            pong_storage_data_177,
            pong_storage_data_176,
            pong_storage_data_175,
            pong_storage_data_174,
            pong_storage_data_173,
            pong_storage_data_172,
            pong_storage_data_171,
            pong_storage_data_170,
            pong_storage_data_169,
            pong_storage_data_168,
            pong_storage_data_167,
            pong_storage_data_166,
            pong_storage_data_165,
            pong_storage_data_164,
            pong_storage_data_163,
            pong_storage_data_162,
            pong_storage_data_161,
            pong_storage_data_160,
            pong_storage_data_159,
            pong_storage_data_158,
            pong_storage_data_157,
            pong_storage_data_156,
            pong_storage_data_155,
            pong_storage_data_154,
            pong_storage_data_153,
            pong_storage_data_152,
            pong_storage_data_151,
            pong_storage_data_150,
            pong_storage_data_149,
            pong_storage_data_148,
            pong_storage_data_147,
            pong_storage_data_146,
            pong_storage_data_145,
            pong_storage_data_144,
            pong_storage_data_143,
            pong_storage_data_142,
            pong_storage_data_141,
            pong_storage_data_140,
            pong_storage_data_139,
            pong_storage_data_138,
            pong_storage_data_137,
            pong_storage_data_136,
            pong_storage_data_135,
            pong_storage_data_134,
            pong_storage_data_133,
            pong_storage_data_132,
            pong_storage_data_131,
            pong_storage_data_130,
            pong_storage_data_129,
            pong_storage_data_128,
            pong_storage_data_127,
            pong_storage_data_126,
            pong_storage_data_125,
            pong_storage_data_124,
            pong_storage_data_123,
            pong_storage_data_122,
            pong_storage_data_121,
            pong_storage_data_120,
            pong_storage_data_119,
            pong_storage_data_118,
            pong_storage_data_117,
            pong_storage_data_116,
            pong_storage_data_115,
            pong_storage_data_114,
            pong_storage_data_113,
            pong_storage_data_112,
            pong_storage_data_111,
            pong_storage_data_110,
            pong_storage_data_109,
            pong_storage_data_108,
            pong_storage_data_107,
            pong_storage_data_106,
            pong_storage_data_105,
            pong_storage_data_104,
            pong_storage_data_103,
            pong_storage_data_102,
            pong_storage_data_101,
            pong_storage_data_100,
            pong_storage_data_99,
            pong_storage_data_98,
            pong_storage_data_97,
            pong_storage_data_96
        };
        2: o_output_data = {
            pong_storage_data_287,
            pong_storage_data_286,
            pong_storage_data_285,
            pong_storage_data_284,
            pong_storage_data_283,
            pong_storage_data_282,
            pong_storage_data_281,
            pong_storage_data_280,
            pong_storage_data_279,
            pong_storage_data_278,
            pong_storage_data_277,
            pong_storage_data_276,
            pong_storage_data_275,
            pong_storage_data_274,
            pong_storage_data_273,
            pong_storage_data_272,
            pong_storage_data_271,
            pong_storage_data_270,
            pong_storage_data_269,
            pong_storage_data_268,
            pong_storage_data_267,
            pong_storage_data_266,
            pong_storage_data_265,
            pong_storage_data_264,
            pong_storage_data_263,
            pong_storage_data_262,
            pong_storage_data_261,
            pong_storage_data_260,
            pong_storage_data_259,
            pong_storage_data_258,
            pong_storage_data_257,
            pong_storage_data_256,
            pong_storage_data_255,
            pong_storage_data_254,
            pong_storage_data_253,
            pong_storage_data_252,
            pong_storage_data_251,
            pong_storage_data_250,
            pong_storage_data_249,
            pong_storage_data_248,
            pong_storage_data_247,
            pong_storage_data_246,
            pong_storage_data_245,
            pong_storage_data_244,
            pong_storage_data_243,
            pong_storage_data_242,
            pong_storage_data_241,
            pong_storage_data_240,
            pong_storage_data_239,
            pong_storage_data_238,
            pong_storage_data_237,
            pong_storage_data_236,
            pong_storage_data_235,
            pong_storage_data_234,
            pong_storage_data_233,
            pong_storage_data_232,
            pong_storage_data_231,
            pong_storage_data_230,
            pong_storage_data_229,
            pong_storage_data_228,
            pong_storage_data_227,
            pong_storage_data_226,
            pong_storage_data_225,
            pong_storage_data_224,
            pong_storage_data_223,
            pong_storage_data_222,
            pong_storage_data_221,
            pong_storage_data_220,
            pong_storage_data_219,
            pong_storage_data_218,
            pong_storage_data_217,
            pong_storage_data_216,
            pong_storage_data_215,
            pong_storage_data_214,
            pong_storage_data_213,
            pong_storage_data_212,
            pong_storage_data_211,
            pong_storage_data_210,
            pong_storage_data_209,
            pong_storage_data_208,
            pong_storage_data_207,
            pong_storage_data_206,
            pong_storage_data_205,
            pong_storage_data_204,
            pong_storage_data_203,
            pong_storage_data_202,
            pong_storage_data_201,
            pong_storage_data_200,
            pong_storage_data_199,
            pong_storage_data_198,
            pong_storage_data_197,
            pong_storage_data_196,
            pong_storage_data_195,
            pong_storage_data_194,
            pong_storage_data_193,
            pong_storage_data_192
        };
        3: o_output_data = {
            pong_storage_data_383,
            pong_storage_data_382,
            pong_storage_data_381,
            pong_storage_data_380,
            pong_storage_data_379,
            pong_storage_data_378,
            pong_storage_data_377,
            pong_storage_data_376,
            pong_storage_data_375,
            pong_storage_data_374,
            pong_storage_data_373,
            pong_storage_data_372,
            pong_storage_data_371,
            pong_storage_data_370,
            pong_storage_data_369,
            pong_storage_data_368,
            pong_storage_data_367,
            pong_storage_data_366,
            pong_storage_data_365,
            pong_storage_data_364,
            pong_storage_data_363,
            pong_storage_data_362,
            pong_storage_data_361,
            pong_storage_data_360,
            pong_storage_data_359,
            pong_storage_data_358,
            pong_storage_data_357,
            pong_storage_data_356,
            pong_storage_data_355,
            pong_storage_data_354,
            pong_storage_data_353,
            pong_storage_data_352,
            pong_storage_data_351,
            pong_storage_data_350,
            pong_storage_data_349,
            pong_storage_data_348,
            pong_storage_data_347,
            pong_storage_data_346,
            pong_storage_data_345,
            pong_storage_data_344,
            pong_storage_data_343,
            pong_storage_data_342,
            pong_storage_data_341,
            pong_storage_data_340,
            pong_storage_data_339,
            pong_storage_data_338,
            pong_storage_data_337,
            pong_storage_data_336,
            pong_storage_data_335,
            pong_storage_data_334,
            pong_storage_data_333,
            pong_storage_data_332,
            pong_storage_data_331,
            pong_storage_data_330,
            pong_storage_data_329,
            pong_storage_data_328,
            pong_storage_data_327,
            pong_storage_data_326,
            pong_storage_data_325,
            pong_storage_data_324,
            pong_storage_data_323,
            pong_storage_data_322,
            pong_storage_data_321,
            pong_storage_data_320,
            pong_storage_data_319,
            pong_storage_data_318,
            pong_storage_data_317,
            pong_storage_data_316,
            pong_storage_data_315,
            pong_storage_data_314,
            pong_storage_data_313,
            pong_storage_data_312,
            pong_storage_data_311,
            pong_storage_data_310,
            pong_storage_data_309,
            pong_storage_data_308,
            pong_storage_data_307,
            pong_storage_data_306,
            pong_storage_data_305,
            pong_storage_data_304,
            pong_storage_data_303,
            pong_storage_data_302,
            pong_storage_data_301,
            pong_storage_data_300,
            pong_storage_data_299,
            pong_storage_data_298,
            pong_storage_data_297,
            pong_storage_data_296,
            pong_storage_data_295,
            pong_storage_data_294,
            pong_storage_data_293,
            pong_storage_data_292,
            pong_storage_data_291,
            pong_storage_data_290,
            pong_storage_data_289,
            pong_storage_data_288
        };
        4: o_output_data = {
            pong_storage_data_479,
            pong_storage_data_478,
            pong_storage_data_477,
            pong_storage_data_476,
            pong_storage_data_475,
            pong_storage_data_474,
            pong_storage_data_473,
            pong_storage_data_472,
            pong_storage_data_471,
            pong_storage_data_470,
            pong_storage_data_469,
            pong_storage_data_468,
            pong_storage_data_467,
            pong_storage_data_466,
            pong_storage_data_465,
            pong_storage_data_464,
            pong_storage_data_463,
            pong_storage_data_462,
            pong_storage_data_461,
            pong_storage_data_460,
            pong_storage_data_459,
            pong_storage_data_458,
            pong_storage_data_457,
            pong_storage_data_456,
            pong_storage_data_455,
            pong_storage_data_454,
            pong_storage_data_453,
            pong_storage_data_452,
            pong_storage_data_451,
            pong_storage_data_450,
            pong_storage_data_449,
            pong_storage_data_448,
            pong_storage_data_447,
            pong_storage_data_446,
            pong_storage_data_445,
            pong_storage_data_444,
            pong_storage_data_443,
            pong_storage_data_442,
            pong_storage_data_441,
            pong_storage_data_440,
            pong_storage_data_439,
            pong_storage_data_438,
            pong_storage_data_437,
            pong_storage_data_436,
            pong_storage_data_435,
            pong_storage_data_434,
            pong_storage_data_433,
            pong_storage_data_432,
            pong_storage_data_431,
            pong_storage_data_430,
            pong_storage_data_429,
            pong_storage_data_428,
            pong_storage_data_427,
            pong_storage_data_426,
            pong_storage_data_425,
            pong_storage_data_424,
            pong_storage_data_423,
            pong_storage_data_422,
            pong_storage_data_421,
            pong_storage_data_420,
            pong_storage_data_419,
            pong_storage_data_418,
            pong_storage_data_417,
            pong_storage_data_416,
            pong_storage_data_415,
            pong_storage_data_414,
            pong_storage_data_413,
            pong_storage_data_412,
            pong_storage_data_411,
            pong_storage_data_410,
            pong_storage_data_409,
            pong_storage_data_408,
            pong_storage_data_407,
            pong_storage_data_406,
            pong_storage_data_405,
            pong_storage_data_404,
            pong_storage_data_403,
            pong_storage_data_402,
            pong_storage_data_401,
            pong_storage_data_400,
            pong_storage_data_399,
            pong_storage_data_398,
            pong_storage_data_397,
            pong_storage_data_396,
            pong_storage_data_395,
            pong_storage_data_394,
            pong_storage_data_393,
            pong_storage_data_392,
            pong_storage_data_391,
            pong_storage_data_390,
            pong_storage_data_389,
            pong_storage_data_388,
            pong_storage_data_387,
            pong_storage_data_386,
            pong_storage_data_385,
            pong_storage_data_384
        };
        5: o_output_data = {
            pong_storage_data_575,
            pong_storage_data_574,
            pong_storage_data_573,
            pong_storage_data_572,
            pong_storage_data_571,
            pong_storage_data_570,
            pong_storage_data_569,
            pong_storage_data_568,
            pong_storage_data_567,
            pong_storage_data_566,
            pong_storage_data_565,
            pong_storage_data_564,
            pong_storage_data_563,
            pong_storage_data_562,
            pong_storage_data_561,
            pong_storage_data_560,
            pong_storage_data_559,
            pong_storage_data_558,
            pong_storage_data_557,
            pong_storage_data_556,
            pong_storage_data_555,
            pong_storage_data_554,
            pong_storage_data_553,
            pong_storage_data_552,
            pong_storage_data_551,
            pong_storage_data_550,
            pong_storage_data_549,
            pong_storage_data_548,
            pong_storage_data_547,
            pong_storage_data_546,
            pong_storage_data_545,
            pong_storage_data_544,
            pong_storage_data_543,
            pong_storage_data_542,
            pong_storage_data_541,
            pong_storage_data_540,
            pong_storage_data_539,
            pong_storage_data_538,
            pong_storage_data_537,
            pong_storage_data_536,
            pong_storage_data_535,
            pong_storage_data_534,
            pong_storage_data_533,
            pong_storage_data_532,
            pong_storage_data_531,
            pong_storage_data_530,
            pong_storage_data_529,
            pong_storage_data_528,
            pong_storage_data_527,
            pong_storage_data_526,
            pong_storage_data_525,
            pong_storage_data_524,
            pong_storage_data_523,
            pong_storage_data_522,
            pong_storage_data_521,
            pong_storage_data_520,
            pong_storage_data_519,
            pong_storage_data_518,
            pong_storage_data_517,
            pong_storage_data_516,
            pong_storage_data_515,
            pong_storage_data_514,
            pong_storage_data_513,
            pong_storage_data_512,
            pong_storage_data_511,
            pong_storage_data_510,
            pong_storage_data_509,
            pong_storage_data_508,
            pong_storage_data_507,
            pong_storage_data_506,
            pong_storage_data_505,
            pong_storage_data_504,
            pong_storage_data_503,
            pong_storage_data_502,
            pong_storage_data_501,
            pong_storage_data_500,
            pong_storage_data_499,
            pong_storage_data_498,
            pong_storage_data_497,
            pong_storage_data_496,
            pong_storage_data_495,
            pong_storage_data_494,
            pong_storage_data_493,
            pong_storage_data_492,
            pong_storage_data_491,
            pong_storage_data_490,
            pong_storage_data_489,
            pong_storage_data_488,
            pong_storage_data_487,
            pong_storage_data_486,
            pong_storage_data_485,
            pong_storage_data_484,
            pong_storage_data_483,
            pong_storage_data_482,
            pong_storage_data_481,
            pong_storage_data_480
        };
        6: o_output_data = {
            pong_storage_data_671,
            pong_storage_data_670,
            pong_storage_data_669,
            pong_storage_data_668,
            pong_storage_data_667,
            pong_storage_data_666,
            pong_storage_data_665,
            pong_storage_data_664,
            pong_storage_data_663,
            pong_storage_data_662,
            pong_storage_data_661,
            pong_storage_data_660,
            pong_storage_data_659,
            pong_storage_data_658,
            pong_storage_data_657,
            pong_storage_data_656,
            pong_storage_data_655,
            pong_storage_data_654,
            pong_storage_data_653,
            pong_storage_data_652,
            pong_storage_data_651,
            pong_storage_data_650,
            pong_storage_data_649,
            pong_storage_data_648,
            pong_storage_data_647,
            pong_storage_data_646,
            pong_storage_data_645,
            pong_storage_data_644,
            pong_storage_data_643,
            pong_storage_data_642,
            pong_storage_data_641,
            pong_storage_data_640,
            pong_storage_data_639,
            pong_storage_data_638,
            pong_storage_data_637,
            pong_storage_data_636,
            pong_storage_data_635,
            pong_storage_data_634,
            pong_storage_data_633,
            pong_storage_data_632,
            pong_storage_data_631,
            pong_storage_data_630,
            pong_storage_data_629,
            pong_storage_data_628,
            pong_storage_data_627,
            pong_storage_data_626,
            pong_storage_data_625,
            pong_storage_data_624,
            pong_storage_data_623,
            pong_storage_data_622,
            pong_storage_data_621,
            pong_storage_data_620,
            pong_storage_data_619,
            pong_storage_data_618,
            pong_storage_data_617,
            pong_storage_data_616,
            pong_storage_data_615,
            pong_storage_data_614,
            pong_storage_data_613,
            pong_storage_data_612,
            pong_storage_data_611,
            pong_storage_data_610,
            pong_storage_data_609,
            pong_storage_data_608,
            pong_storage_data_607,
            pong_storage_data_606,
            pong_storage_data_605,
            pong_storage_data_604,
            pong_storage_data_603,
            pong_storage_data_602,
            pong_storage_data_601,
            pong_storage_data_600,
            pong_storage_data_599,
            pong_storage_data_598,
            pong_storage_data_597,
            pong_storage_data_596,
            pong_storage_data_595,
            pong_storage_data_594,
            pong_storage_data_593,
            pong_storage_data_592,
            pong_storage_data_591,
            pong_storage_data_590,
            pong_storage_data_589,
            pong_storage_data_588,
            pong_storage_data_587,
            pong_storage_data_586,
            pong_storage_data_585,
            pong_storage_data_584,
            pong_storage_data_583,
            pong_storage_data_582,
            pong_storage_data_581,
            pong_storage_data_580,
            pong_storage_data_579,
            pong_storage_data_578,
            pong_storage_data_577,
            pong_storage_data_576
        };
        7: o_output_data = {
            pong_storage_data_767,
            pong_storage_data_766,
            pong_storage_data_765,
            pong_storage_data_764,
            pong_storage_data_763,
            pong_storage_data_762,
            pong_storage_data_761,
            pong_storage_data_760,
            pong_storage_data_759,
            pong_storage_data_758,
            pong_storage_data_757,
            pong_storage_data_756,
            pong_storage_data_755,
            pong_storage_data_754,
            pong_storage_data_753,
            pong_storage_data_752,
            pong_storage_data_751,
            pong_storage_data_750,
            pong_storage_data_749,
            pong_storage_data_748,
            pong_storage_data_747,
            pong_storage_data_746,
            pong_storage_data_745,
            pong_storage_data_744,
            pong_storage_data_743,
            pong_storage_data_742,
            pong_storage_data_741,
            pong_storage_data_740,
            pong_storage_data_739,
            pong_storage_data_738,
            pong_storage_data_737,
            pong_storage_data_736,
            pong_storage_data_735,
            pong_storage_data_734,
            pong_storage_data_733,
            pong_storage_data_732,
            pong_storage_data_731,
            pong_storage_data_730,
            pong_storage_data_729,
            pong_storage_data_728,
            pong_storage_data_727,
            pong_storage_data_726,
            pong_storage_data_725,
            pong_storage_data_724,
            pong_storage_data_723,
            pong_storage_data_722,
            pong_storage_data_721,
            pong_storage_data_720,
            pong_storage_data_719,
            pong_storage_data_718,
            pong_storage_data_717,
            pong_storage_data_716,
            pong_storage_data_715,
            pong_storage_data_714,
            pong_storage_data_713,
            pong_storage_data_712,
            pong_storage_data_711,
            pong_storage_data_710,
            pong_storage_data_709,
            pong_storage_data_708,
            pong_storage_data_707,
            pong_storage_data_706,
            pong_storage_data_705,
            pong_storage_data_704,
            pong_storage_data_703,
            pong_storage_data_702,
            pong_storage_data_701,
            pong_storage_data_700,
            pong_storage_data_699,
            pong_storage_data_698,
            pong_storage_data_697,
            pong_storage_data_696,
            pong_storage_data_695,
            pong_storage_data_694,
            pong_storage_data_693,
            pong_storage_data_692,
            pong_storage_data_691,
            pong_storage_data_690,
            pong_storage_data_689,
            pong_storage_data_688,
            pong_storage_data_687,
            pong_storage_data_686,
            pong_storage_data_685,
            pong_storage_data_684,
            pong_storage_data_683,
            pong_storage_data_682,
            pong_storage_data_681,
            pong_storage_data_680,
            pong_storage_data_679,
            pong_storage_data_678,
            pong_storage_data_677,
            pong_storage_data_676,
            pong_storage_data_675,
            pong_storage_data_674,
            pong_storage_data_673,
            pong_storage_data_672
        };
        8: o_output_data = {
            pong_storage_data_863,
            pong_storage_data_862,
            pong_storage_data_861,
            pong_storage_data_860,
            pong_storage_data_859,
            pong_storage_data_858,
            pong_storage_data_857,
            pong_storage_data_856,
            pong_storage_data_855,
            pong_storage_data_854,
            pong_storage_data_853,
            pong_storage_data_852,
            pong_storage_data_851,
            pong_storage_data_850,
            pong_storage_data_849,
            pong_storage_data_848,
            pong_storage_data_847,
            pong_storage_data_846,
            pong_storage_data_845,
            pong_storage_data_844,
            pong_storage_data_843,
            pong_storage_data_842,
            pong_storage_data_841,
            pong_storage_data_840,
            pong_storage_data_839,
            pong_storage_data_838,
            pong_storage_data_837,
            pong_storage_data_836,
            pong_storage_data_835,
            pong_storage_data_834,
            pong_storage_data_833,
            pong_storage_data_832,
            pong_storage_data_831,
            pong_storage_data_830,
            pong_storage_data_829,
            pong_storage_data_828,
            pong_storage_data_827,
            pong_storage_data_826,
            pong_storage_data_825,
            pong_storage_data_824,
            pong_storage_data_823,
            pong_storage_data_822,
            pong_storage_data_821,
            pong_storage_data_820,
            pong_storage_data_819,
            pong_storage_data_818,
            pong_storage_data_817,
            pong_storage_data_816,
            pong_storage_data_815,
            pong_storage_data_814,
            pong_storage_data_813,
            pong_storage_data_812,
            pong_storage_data_811,
            pong_storage_data_810,
            pong_storage_data_809,
            pong_storage_data_808,
            pong_storage_data_807,
            pong_storage_data_806,
            pong_storage_data_805,
            pong_storage_data_804,
            pong_storage_data_803,
            pong_storage_data_802,
            pong_storage_data_801,
            pong_storage_data_800,
            pong_storage_data_799,
            pong_storage_data_798,
            pong_storage_data_797,
            pong_storage_data_796,
            pong_storage_data_795,
            pong_storage_data_794,
            pong_storage_data_793,
            pong_storage_data_792,
            pong_storage_data_791,
            pong_storage_data_790,
            pong_storage_data_789,
            pong_storage_data_788,
            pong_storage_data_787,
            pong_storage_data_786,
            pong_storage_data_785,
            pong_storage_data_784,
            pong_storage_data_783,
            pong_storage_data_782,
            pong_storage_data_781,
            pong_storage_data_780,
            pong_storage_data_779,
            pong_storage_data_778,
            pong_storage_data_777,
            pong_storage_data_776,
            pong_storage_data_775,
            pong_storage_data_774,
            pong_storage_data_773,
            pong_storage_data_772,
            pong_storage_data_771,
            pong_storage_data_770,
            pong_storage_data_769,
            pong_storage_data_768
        };
        9: o_output_data = {
            pong_storage_data_959,
            pong_storage_data_958,
            pong_storage_data_957,
            pong_storage_data_956,
            pong_storage_data_955,
            pong_storage_data_954,
            pong_storage_data_953,
            pong_storage_data_952,
            pong_storage_data_951,
            pong_storage_data_950,
            pong_storage_data_949,
            pong_storage_data_948,
            pong_storage_data_947,
            pong_storage_data_946,
            pong_storage_data_945,
            pong_storage_data_944,
            pong_storage_data_943,
            pong_storage_data_942,
            pong_storage_data_941,
            pong_storage_data_940,
            pong_storage_data_939,
            pong_storage_data_938,
            pong_storage_data_937,
            pong_storage_data_936,
            pong_storage_data_935,
            pong_storage_data_934,
            pong_storage_data_933,
            pong_storage_data_932,
            pong_storage_data_931,
            pong_storage_data_930,
            pong_storage_data_929,
            pong_storage_data_928,
            pong_storage_data_927,
            pong_storage_data_926,
            pong_storage_data_925,
            pong_storage_data_924,
            pong_storage_data_923,
            pong_storage_data_922,
            pong_storage_data_921,
            pong_storage_data_920,
            pong_storage_data_919,
            pong_storage_data_918,
            pong_storage_data_917,
            pong_storage_data_916,
            pong_storage_data_915,
            pong_storage_data_914,
            pong_storage_data_913,
            pong_storage_data_912,
            pong_storage_data_911,
            pong_storage_data_910,
            pong_storage_data_909,
            pong_storage_data_908,
            pong_storage_data_907,
            pong_storage_data_906,
            pong_storage_data_905,
            pong_storage_data_904,
            pong_storage_data_903,
            pong_storage_data_902,
            pong_storage_data_901,
            pong_storage_data_900,
            pong_storage_data_899,
            pong_storage_data_898,
            pong_storage_data_897,
            pong_storage_data_896,
            pong_storage_data_895,
            pong_storage_data_894,
            pong_storage_data_893,
            pong_storage_data_892,
            pong_storage_data_891,
            pong_storage_data_890,
            pong_storage_data_889,
            pong_storage_data_888,
            pong_storage_data_887,
            pong_storage_data_886,
            pong_storage_data_885,
            pong_storage_data_884,
            pong_storage_data_883,
            pong_storage_data_882,
            pong_storage_data_881,
            pong_storage_data_880,
            pong_storage_data_879,
            pong_storage_data_878,
            pong_storage_data_877,
            pong_storage_data_876,
            pong_storage_data_875,
            pong_storage_data_874,
            pong_storage_data_873,
            pong_storage_data_872,
            pong_storage_data_871,
            pong_storage_data_870,
            pong_storage_data_869,
            pong_storage_data_868,
            pong_storage_data_867,
            pong_storage_data_866,
            pong_storage_data_865,
            pong_storage_data_864
        };
        default: o_output_data = {
            pong_storage_data_1055,
            pong_storage_data_1054,
            pong_storage_data_1053,
            pong_storage_data_1052,
            pong_storage_data_1051,
            pong_storage_data_1050,
            pong_storage_data_1049,
            pong_storage_data_1048,
            pong_storage_data_1047,
            pong_storage_data_1046,
            pong_storage_data_1045,
            pong_storage_data_1044,
            pong_storage_data_1043,
            pong_storage_data_1042,
            pong_storage_data_1041,
            pong_storage_data_1040,
            pong_storage_data_1039,
            pong_storage_data_1038,
            pong_storage_data_1037,
            pong_storage_data_1036,
            pong_storage_data_1035,
            pong_storage_data_1034,
            pong_storage_data_1033,
            pong_storage_data_1032,
            pong_storage_data_1031,
            pong_storage_data_1030,
            pong_storage_data_1029,
            pong_storage_data_1028,
            pong_storage_data_1027,
            pong_storage_data_1026,
            pong_storage_data_1025,
            pong_storage_data_1024,
            pong_storage_data_1023,
            pong_storage_data_1022,
            pong_storage_data_1021,
            pong_storage_data_1020,
            pong_storage_data_1019,
            pong_storage_data_1018,
            pong_storage_data_1017,
            pong_storage_data_1016,
            pong_storage_data_1015,
            pong_storage_data_1014,
            pong_storage_data_1013,
            pong_storage_data_1012,
            pong_storage_data_1011,
            pong_storage_data_1010,
            pong_storage_data_1009,
            pong_storage_data_1008,
            pong_storage_data_1007,
            pong_storage_data_1006,
            pong_storage_data_1005,
            pong_storage_data_1004,
            pong_storage_data_1003,
            pong_storage_data_1002,
            pong_storage_data_1001,
            pong_storage_data_1000,
            pong_storage_data_999,
            pong_storage_data_998,
            pong_storage_data_997,
            pong_storage_data_996,
            pong_storage_data_995,
            pong_storage_data_994,
            pong_storage_data_993,
            pong_storage_data_992,
            pong_storage_data_991,
            pong_storage_data_990,
            pong_storage_data_989,
            pong_storage_data_988,
            pong_storage_data_987,
            pong_storage_data_986,
            pong_storage_data_985,
            pong_storage_data_984,
            pong_storage_data_983,
            pong_storage_data_982,
            pong_storage_data_981,
            pong_storage_data_980,
            pong_storage_data_979,
            pong_storage_data_978,
            pong_storage_data_977,
            pong_storage_data_976,
            pong_storage_data_975,
            pong_storage_data_974,
            pong_storage_data_973,
            pong_storage_data_972,
            pong_storage_data_971,
            pong_storage_data_970,
            pong_storage_data_969,
            pong_storage_data_968,
            pong_storage_data_967,
            pong_storage_data_966,
            pong_storage_data_965,
            pong_storage_data_964,
            pong_storage_data_963,
            pong_storage_data_962,
            pong_storage_data_961,
            pong_storage_data_960
        };
        endcase
        o_output_valid = 1'b1;
    end
    ST_WAIT_FOR_PING: begin
        if (ping_is_full == 1'b1) begin
            next_readout_state = ST_PING;
        end else begin
            next_readout_state = ST_WAIT_FOR_PING;
        end
        o_output_data = 0;
        o_output_valid = 1'b0;
    end
    ST_WAIT_FOR_PONG: begin
        if (pong_is_full == 1'b1) begin
            next_readout_state = ST_PONG;
        end else begin
            next_readout_state = ST_WAIT_FOR_PONG;
        end
        o_output_data = 0;
        o_output_valid = 1'b0;
    end
    default: begin // ST_INIT
        next_readout_state = ST_WAIT_FOR_PING;
        o_output_data = 0;
        o_output_valid = 1'b0;
    end
    endcase
end

logic ping_storage_data_0;
logic pong_storage_data_0;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_0 <= 1'b0;
        pong_storage_data_0 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                98 / IN_WIDTH: ping_storage_data_0 <= (fillup_transition == 1'b1) ? i_input_data[98 % IN_WIDTH] : ping_storage_data_0 ^ i_input_data[98 % IN_WIDTH];
                215 / IN_WIDTH: ping_storage_data_0 <= (fillup_transition == 1'b1) ? i_input_data[215 % IN_WIDTH] : ping_storage_data_0 ^ i_input_data[215 % IN_WIDTH];
                809 / IN_WIDTH: ping_storage_data_0 <= (fillup_transition == 1'b1) ? i_input_data[809 % IN_WIDTH] : ping_storage_data_0 ^ i_input_data[809 % IN_WIDTH];
                877 / IN_WIDTH: ping_storage_data_0 <= (fillup_transition == 1'b1) ? i_input_data[877 % IN_WIDTH] : ping_storage_data_0 ^ i_input_data[877 % IN_WIDTH];
                default: ping_storage_data_0 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_0;
                endcase
            end else begin
                case (input_count)
                98 / IN_WIDTH: pong_storage_data_0 <= (fillup_transition == 1'b1) ? i_input_data[98 % IN_WIDTH] : pong_storage_data_0 ^ i_input_data[98 % IN_WIDTH];
                215 / IN_WIDTH: pong_storage_data_0 <= (fillup_transition == 1'b1) ? i_input_data[215 % IN_WIDTH] : pong_storage_data_0 ^ i_input_data[215 % IN_WIDTH];
                809 / IN_WIDTH: pong_storage_data_0 <= (fillup_transition == 1'b1) ? i_input_data[809 % IN_WIDTH] : pong_storage_data_0 ^ i_input_data[809 % IN_WIDTH];
                877 / IN_WIDTH: pong_storage_data_0 <= (fillup_transition == 1'b1) ? i_input_data[877 % IN_WIDTH] : pong_storage_data_0 ^ i_input_data[877 % IN_WIDTH];
                default: pong_storage_data_0 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_0;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_0 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_0;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_0 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_0;
            end
        end
    end
end

logic ping_storage_data_1;
logic pong_storage_data_1;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1 <= 1'b0;
        pong_storage_data_1 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                99 / IN_WIDTH: ping_storage_data_1 <= (fillup_transition == 1'b1) ? i_input_data[99 % IN_WIDTH] : ping_storage_data_1 ^ i_input_data[99 % IN_WIDTH];
                216 / IN_WIDTH: ping_storage_data_1 <= (fillup_transition == 1'b1) ? i_input_data[216 % IN_WIDTH] : ping_storage_data_1 ^ i_input_data[216 % IN_WIDTH];
                810 / IN_WIDTH: ping_storage_data_1 <= (fillup_transition == 1'b1) ? i_input_data[810 % IN_WIDTH] : ping_storage_data_1 ^ i_input_data[810 % IN_WIDTH];
                878 / IN_WIDTH: ping_storage_data_1 <= (fillup_transition == 1'b1) ? i_input_data[878 % IN_WIDTH] : ping_storage_data_1 ^ i_input_data[878 % IN_WIDTH];
                default: ping_storage_data_1 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1;
                endcase
            end else begin
                case (input_count)
                99 / IN_WIDTH: pong_storage_data_1 <= (fillup_transition == 1'b1) ? i_input_data[99 % IN_WIDTH] : pong_storage_data_1 ^ i_input_data[99 % IN_WIDTH];
                216 / IN_WIDTH: pong_storage_data_1 <= (fillup_transition == 1'b1) ? i_input_data[216 % IN_WIDTH] : pong_storage_data_1 ^ i_input_data[216 % IN_WIDTH];
                810 / IN_WIDTH: pong_storage_data_1 <= (fillup_transition == 1'b1) ? i_input_data[810 % IN_WIDTH] : pong_storage_data_1 ^ i_input_data[810 % IN_WIDTH];
                878 / IN_WIDTH: pong_storage_data_1 <= (fillup_transition == 1'b1) ? i_input_data[878 % IN_WIDTH] : pong_storage_data_1 ^ i_input_data[878 % IN_WIDTH];
                default: pong_storage_data_1 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1;
            end
        end
    end
end

logic ping_storage_data_2;
logic pong_storage_data_2;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_2 <= 1'b0;
        pong_storage_data_2 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                100 / IN_WIDTH: ping_storage_data_2 <= (fillup_transition == 1'b1) ? i_input_data[100 % IN_WIDTH] : ping_storage_data_2 ^ i_input_data[100 % IN_WIDTH];
                217 / IN_WIDTH: ping_storage_data_2 <= (fillup_transition == 1'b1) ? i_input_data[217 % IN_WIDTH] : ping_storage_data_2 ^ i_input_data[217 % IN_WIDTH];
                811 / IN_WIDTH: ping_storage_data_2 <= (fillup_transition == 1'b1) ? i_input_data[811 % IN_WIDTH] : ping_storage_data_2 ^ i_input_data[811 % IN_WIDTH];
                879 / IN_WIDTH: ping_storage_data_2 <= (fillup_transition == 1'b1) ? i_input_data[879 % IN_WIDTH] : ping_storage_data_2 ^ i_input_data[879 % IN_WIDTH];
                default: ping_storage_data_2 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_2;
                endcase
            end else begin
                case (input_count)
                100 / IN_WIDTH: pong_storage_data_2 <= (fillup_transition == 1'b1) ? i_input_data[100 % IN_WIDTH] : pong_storage_data_2 ^ i_input_data[100 % IN_WIDTH];
                217 / IN_WIDTH: pong_storage_data_2 <= (fillup_transition == 1'b1) ? i_input_data[217 % IN_WIDTH] : pong_storage_data_2 ^ i_input_data[217 % IN_WIDTH];
                811 / IN_WIDTH: pong_storage_data_2 <= (fillup_transition == 1'b1) ? i_input_data[811 % IN_WIDTH] : pong_storage_data_2 ^ i_input_data[811 % IN_WIDTH];
                879 / IN_WIDTH: pong_storage_data_2 <= (fillup_transition == 1'b1) ? i_input_data[879 % IN_WIDTH] : pong_storage_data_2 ^ i_input_data[879 % IN_WIDTH];
                default: pong_storage_data_2 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_2;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_2 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_2;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_2 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_2;
            end
        end
    end
end

logic ping_storage_data_3;
logic pong_storage_data_3;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_3 <= 1'b0;
        pong_storage_data_3 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                101 / IN_WIDTH: ping_storage_data_3 <= (fillup_transition == 1'b1) ? i_input_data[101 % IN_WIDTH] : ping_storage_data_3 ^ i_input_data[101 % IN_WIDTH];
                218 / IN_WIDTH: ping_storage_data_3 <= (fillup_transition == 1'b1) ? i_input_data[218 % IN_WIDTH] : ping_storage_data_3 ^ i_input_data[218 % IN_WIDTH];
                812 / IN_WIDTH: ping_storage_data_3 <= (fillup_transition == 1'b1) ? i_input_data[812 % IN_WIDTH] : ping_storage_data_3 ^ i_input_data[812 % IN_WIDTH];
                880 / IN_WIDTH: ping_storage_data_3 <= (fillup_transition == 1'b1) ? i_input_data[880 % IN_WIDTH] : ping_storage_data_3 ^ i_input_data[880 % IN_WIDTH];
                default: ping_storage_data_3 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_3;
                endcase
            end else begin
                case (input_count)
                101 / IN_WIDTH: pong_storage_data_3 <= (fillup_transition == 1'b1) ? i_input_data[101 % IN_WIDTH] : pong_storage_data_3 ^ i_input_data[101 % IN_WIDTH];
                218 / IN_WIDTH: pong_storage_data_3 <= (fillup_transition == 1'b1) ? i_input_data[218 % IN_WIDTH] : pong_storage_data_3 ^ i_input_data[218 % IN_WIDTH];
                812 / IN_WIDTH: pong_storage_data_3 <= (fillup_transition == 1'b1) ? i_input_data[812 % IN_WIDTH] : pong_storage_data_3 ^ i_input_data[812 % IN_WIDTH];
                880 / IN_WIDTH: pong_storage_data_3 <= (fillup_transition == 1'b1) ? i_input_data[880 % IN_WIDTH] : pong_storage_data_3 ^ i_input_data[880 % IN_WIDTH];
                default: pong_storage_data_3 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_3;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_3 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_3;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_3 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_3;
            end
        end
    end
end

logic ping_storage_data_4;
logic pong_storage_data_4;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_4 <= 1'b0;
        pong_storage_data_4 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                102 / IN_WIDTH: ping_storage_data_4 <= (fillup_transition == 1'b1) ? i_input_data[102 % IN_WIDTH] : ping_storage_data_4 ^ i_input_data[102 % IN_WIDTH];
                219 / IN_WIDTH: ping_storage_data_4 <= (fillup_transition == 1'b1) ? i_input_data[219 % IN_WIDTH] : ping_storage_data_4 ^ i_input_data[219 % IN_WIDTH];
                813 / IN_WIDTH: ping_storage_data_4 <= (fillup_transition == 1'b1) ? i_input_data[813 % IN_WIDTH] : ping_storage_data_4 ^ i_input_data[813 % IN_WIDTH];
                881 / IN_WIDTH: ping_storage_data_4 <= (fillup_transition == 1'b1) ? i_input_data[881 % IN_WIDTH] : ping_storage_data_4 ^ i_input_data[881 % IN_WIDTH];
                default: ping_storage_data_4 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_4;
                endcase
            end else begin
                case (input_count)
                102 / IN_WIDTH: pong_storage_data_4 <= (fillup_transition == 1'b1) ? i_input_data[102 % IN_WIDTH] : pong_storage_data_4 ^ i_input_data[102 % IN_WIDTH];
                219 / IN_WIDTH: pong_storage_data_4 <= (fillup_transition == 1'b1) ? i_input_data[219 % IN_WIDTH] : pong_storage_data_4 ^ i_input_data[219 % IN_WIDTH];
                813 / IN_WIDTH: pong_storage_data_4 <= (fillup_transition == 1'b1) ? i_input_data[813 % IN_WIDTH] : pong_storage_data_4 ^ i_input_data[813 % IN_WIDTH];
                881 / IN_WIDTH: pong_storage_data_4 <= (fillup_transition == 1'b1) ? i_input_data[881 % IN_WIDTH] : pong_storage_data_4 ^ i_input_data[881 % IN_WIDTH];
                default: pong_storage_data_4 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_4;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_4 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_4;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_4 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_4;
            end
        end
    end
end

logic ping_storage_data_5;
logic pong_storage_data_5;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_5 <= 1'b0;
        pong_storage_data_5 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                103 / IN_WIDTH: ping_storage_data_5 <= (fillup_transition == 1'b1) ? i_input_data[103 % IN_WIDTH] : ping_storage_data_5 ^ i_input_data[103 % IN_WIDTH];
                220 / IN_WIDTH: ping_storage_data_5 <= (fillup_transition == 1'b1) ? i_input_data[220 % IN_WIDTH] : ping_storage_data_5 ^ i_input_data[220 % IN_WIDTH];
                814 / IN_WIDTH: ping_storage_data_5 <= (fillup_transition == 1'b1) ? i_input_data[814 % IN_WIDTH] : ping_storage_data_5 ^ i_input_data[814 % IN_WIDTH];
                882 / IN_WIDTH: ping_storage_data_5 <= (fillup_transition == 1'b1) ? i_input_data[882 % IN_WIDTH] : ping_storage_data_5 ^ i_input_data[882 % IN_WIDTH];
                default: ping_storage_data_5 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_5;
                endcase
            end else begin
                case (input_count)
                103 / IN_WIDTH: pong_storage_data_5 <= (fillup_transition == 1'b1) ? i_input_data[103 % IN_WIDTH] : pong_storage_data_5 ^ i_input_data[103 % IN_WIDTH];
                220 / IN_WIDTH: pong_storage_data_5 <= (fillup_transition == 1'b1) ? i_input_data[220 % IN_WIDTH] : pong_storage_data_5 ^ i_input_data[220 % IN_WIDTH];
                814 / IN_WIDTH: pong_storage_data_5 <= (fillup_transition == 1'b1) ? i_input_data[814 % IN_WIDTH] : pong_storage_data_5 ^ i_input_data[814 % IN_WIDTH];
                882 / IN_WIDTH: pong_storage_data_5 <= (fillup_transition == 1'b1) ? i_input_data[882 % IN_WIDTH] : pong_storage_data_5 ^ i_input_data[882 % IN_WIDTH];
                default: pong_storage_data_5 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_5;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_5 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_5;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_5 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_5;
            end
        end
    end
end

logic ping_storage_data_6;
logic pong_storage_data_6;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_6 <= 1'b0;
        pong_storage_data_6 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                104 / IN_WIDTH: ping_storage_data_6 <= (fillup_transition == 1'b1) ? i_input_data[104 % IN_WIDTH] : ping_storage_data_6 ^ i_input_data[104 % IN_WIDTH];
                221 / IN_WIDTH: ping_storage_data_6 <= (fillup_transition == 1'b1) ? i_input_data[221 % IN_WIDTH] : ping_storage_data_6 ^ i_input_data[221 % IN_WIDTH];
                815 / IN_WIDTH: ping_storage_data_6 <= (fillup_transition == 1'b1) ? i_input_data[815 % IN_WIDTH] : ping_storage_data_6 ^ i_input_data[815 % IN_WIDTH];
                883 / IN_WIDTH: ping_storage_data_6 <= (fillup_transition == 1'b1) ? i_input_data[883 % IN_WIDTH] : ping_storage_data_6 ^ i_input_data[883 % IN_WIDTH];
                default: ping_storage_data_6 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_6;
                endcase
            end else begin
                case (input_count)
                104 / IN_WIDTH: pong_storage_data_6 <= (fillup_transition == 1'b1) ? i_input_data[104 % IN_WIDTH] : pong_storage_data_6 ^ i_input_data[104 % IN_WIDTH];
                221 / IN_WIDTH: pong_storage_data_6 <= (fillup_transition == 1'b1) ? i_input_data[221 % IN_WIDTH] : pong_storage_data_6 ^ i_input_data[221 % IN_WIDTH];
                815 / IN_WIDTH: pong_storage_data_6 <= (fillup_transition == 1'b1) ? i_input_data[815 % IN_WIDTH] : pong_storage_data_6 ^ i_input_data[815 % IN_WIDTH];
                883 / IN_WIDTH: pong_storage_data_6 <= (fillup_transition == 1'b1) ? i_input_data[883 % IN_WIDTH] : pong_storage_data_6 ^ i_input_data[883 % IN_WIDTH];
                default: pong_storage_data_6 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_6;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_6 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_6;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_6 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_6;
            end
        end
    end
end

logic ping_storage_data_7;
logic pong_storage_data_7;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_7 <= 1'b0;
        pong_storage_data_7 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                105 / IN_WIDTH: ping_storage_data_7 <= (fillup_transition == 1'b1) ? i_input_data[105 % IN_WIDTH] : ping_storage_data_7 ^ i_input_data[105 % IN_WIDTH];
                222 / IN_WIDTH: ping_storage_data_7 <= (fillup_transition == 1'b1) ? i_input_data[222 % IN_WIDTH] : ping_storage_data_7 ^ i_input_data[222 % IN_WIDTH];
                816 / IN_WIDTH: ping_storage_data_7 <= (fillup_transition == 1'b1) ? i_input_data[816 % IN_WIDTH] : ping_storage_data_7 ^ i_input_data[816 % IN_WIDTH];
                884 / IN_WIDTH: ping_storage_data_7 <= (fillup_transition == 1'b1) ? i_input_data[884 % IN_WIDTH] : ping_storage_data_7 ^ i_input_data[884 % IN_WIDTH];
                default: ping_storage_data_7 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_7;
                endcase
            end else begin
                case (input_count)
                105 / IN_WIDTH: pong_storage_data_7 <= (fillup_transition == 1'b1) ? i_input_data[105 % IN_WIDTH] : pong_storage_data_7 ^ i_input_data[105 % IN_WIDTH];
                222 / IN_WIDTH: pong_storage_data_7 <= (fillup_transition == 1'b1) ? i_input_data[222 % IN_WIDTH] : pong_storage_data_7 ^ i_input_data[222 % IN_WIDTH];
                816 / IN_WIDTH: pong_storage_data_7 <= (fillup_transition == 1'b1) ? i_input_data[816 % IN_WIDTH] : pong_storage_data_7 ^ i_input_data[816 % IN_WIDTH];
                884 / IN_WIDTH: pong_storage_data_7 <= (fillup_transition == 1'b1) ? i_input_data[884 % IN_WIDTH] : pong_storage_data_7 ^ i_input_data[884 % IN_WIDTH];
                default: pong_storage_data_7 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_7;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_7 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_7;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_7 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_7;
            end
        end
    end
end

logic ping_storage_data_8;
logic pong_storage_data_8;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_8 <= 1'b0;
        pong_storage_data_8 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                106 / IN_WIDTH: ping_storage_data_8 <= (fillup_transition == 1'b1) ? i_input_data[106 % IN_WIDTH] : ping_storage_data_8 ^ i_input_data[106 % IN_WIDTH];
                223 / IN_WIDTH: ping_storage_data_8 <= (fillup_transition == 1'b1) ? i_input_data[223 % IN_WIDTH] : ping_storage_data_8 ^ i_input_data[223 % IN_WIDTH];
                817 / IN_WIDTH: ping_storage_data_8 <= (fillup_transition == 1'b1) ? i_input_data[817 % IN_WIDTH] : ping_storage_data_8 ^ i_input_data[817 % IN_WIDTH];
                885 / IN_WIDTH: ping_storage_data_8 <= (fillup_transition == 1'b1) ? i_input_data[885 % IN_WIDTH] : ping_storage_data_8 ^ i_input_data[885 % IN_WIDTH];
                default: ping_storage_data_8 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_8;
                endcase
            end else begin
                case (input_count)
                106 / IN_WIDTH: pong_storage_data_8 <= (fillup_transition == 1'b1) ? i_input_data[106 % IN_WIDTH] : pong_storage_data_8 ^ i_input_data[106 % IN_WIDTH];
                223 / IN_WIDTH: pong_storage_data_8 <= (fillup_transition == 1'b1) ? i_input_data[223 % IN_WIDTH] : pong_storage_data_8 ^ i_input_data[223 % IN_WIDTH];
                817 / IN_WIDTH: pong_storage_data_8 <= (fillup_transition == 1'b1) ? i_input_data[817 % IN_WIDTH] : pong_storage_data_8 ^ i_input_data[817 % IN_WIDTH];
                885 / IN_WIDTH: pong_storage_data_8 <= (fillup_transition == 1'b1) ? i_input_data[885 % IN_WIDTH] : pong_storage_data_8 ^ i_input_data[885 % IN_WIDTH];
                default: pong_storage_data_8 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_8;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_8 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_8;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_8 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_8;
            end
        end
    end
end

logic ping_storage_data_9;
logic pong_storage_data_9;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_9 <= 1'b0;
        pong_storage_data_9 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                107 / IN_WIDTH: ping_storage_data_9 <= (fillup_transition == 1'b1) ? i_input_data[107 % IN_WIDTH] : ping_storage_data_9 ^ i_input_data[107 % IN_WIDTH];
                224 / IN_WIDTH: ping_storage_data_9 <= (fillup_transition == 1'b1) ? i_input_data[224 % IN_WIDTH] : ping_storage_data_9 ^ i_input_data[224 % IN_WIDTH];
                818 / IN_WIDTH: ping_storage_data_9 <= (fillup_transition == 1'b1) ? i_input_data[818 % IN_WIDTH] : ping_storage_data_9 ^ i_input_data[818 % IN_WIDTH];
                886 / IN_WIDTH: ping_storage_data_9 <= (fillup_transition == 1'b1) ? i_input_data[886 % IN_WIDTH] : ping_storage_data_9 ^ i_input_data[886 % IN_WIDTH];
                default: ping_storage_data_9 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_9;
                endcase
            end else begin
                case (input_count)
                107 / IN_WIDTH: pong_storage_data_9 <= (fillup_transition == 1'b1) ? i_input_data[107 % IN_WIDTH] : pong_storage_data_9 ^ i_input_data[107 % IN_WIDTH];
                224 / IN_WIDTH: pong_storage_data_9 <= (fillup_transition == 1'b1) ? i_input_data[224 % IN_WIDTH] : pong_storage_data_9 ^ i_input_data[224 % IN_WIDTH];
                818 / IN_WIDTH: pong_storage_data_9 <= (fillup_transition == 1'b1) ? i_input_data[818 % IN_WIDTH] : pong_storage_data_9 ^ i_input_data[818 % IN_WIDTH];
                886 / IN_WIDTH: pong_storage_data_9 <= (fillup_transition == 1'b1) ? i_input_data[886 % IN_WIDTH] : pong_storage_data_9 ^ i_input_data[886 % IN_WIDTH];
                default: pong_storage_data_9 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_9;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_9 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_9;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_9 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_9;
            end
        end
    end
end

logic ping_storage_data_10;
logic pong_storage_data_10;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_10 <= 1'b0;
        pong_storage_data_10 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                108 / IN_WIDTH: ping_storage_data_10 <= (fillup_transition == 1'b1) ? i_input_data[108 % IN_WIDTH] : ping_storage_data_10 ^ i_input_data[108 % IN_WIDTH];
                225 / IN_WIDTH: ping_storage_data_10 <= (fillup_transition == 1'b1) ? i_input_data[225 % IN_WIDTH] : ping_storage_data_10 ^ i_input_data[225 % IN_WIDTH];
                819 / IN_WIDTH: ping_storage_data_10 <= (fillup_transition == 1'b1) ? i_input_data[819 % IN_WIDTH] : ping_storage_data_10 ^ i_input_data[819 % IN_WIDTH];
                887 / IN_WIDTH: ping_storage_data_10 <= (fillup_transition == 1'b1) ? i_input_data[887 % IN_WIDTH] : ping_storage_data_10 ^ i_input_data[887 % IN_WIDTH];
                default: ping_storage_data_10 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_10;
                endcase
            end else begin
                case (input_count)
                108 / IN_WIDTH: pong_storage_data_10 <= (fillup_transition == 1'b1) ? i_input_data[108 % IN_WIDTH] : pong_storage_data_10 ^ i_input_data[108 % IN_WIDTH];
                225 / IN_WIDTH: pong_storage_data_10 <= (fillup_transition == 1'b1) ? i_input_data[225 % IN_WIDTH] : pong_storage_data_10 ^ i_input_data[225 % IN_WIDTH];
                819 / IN_WIDTH: pong_storage_data_10 <= (fillup_transition == 1'b1) ? i_input_data[819 % IN_WIDTH] : pong_storage_data_10 ^ i_input_data[819 % IN_WIDTH];
                887 / IN_WIDTH: pong_storage_data_10 <= (fillup_transition == 1'b1) ? i_input_data[887 % IN_WIDTH] : pong_storage_data_10 ^ i_input_data[887 % IN_WIDTH];
                default: pong_storage_data_10 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_10;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_10 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_10;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_10 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_10;
            end
        end
    end
end

logic ping_storage_data_11;
logic pong_storage_data_11;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_11 <= 1'b0;
        pong_storage_data_11 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                109 / IN_WIDTH: ping_storage_data_11 <= (fillup_transition == 1'b1) ? i_input_data[109 % IN_WIDTH] : ping_storage_data_11 ^ i_input_data[109 % IN_WIDTH];
                226 / IN_WIDTH: ping_storage_data_11 <= (fillup_transition == 1'b1) ? i_input_data[226 % IN_WIDTH] : ping_storage_data_11 ^ i_input_data[226 % IN_WIDTH];
                820 / IN_WIDTH: ping_storage_data_11 <= (fillup_transition == 1'b1) ? i_input_data[820 % IN_WIDTH] : ping_storage_data_11 ^ i_input_data[820 % IN_WIDTH];
                888 / IN_WIDTH: ping_storage_data_11 <= (fillup_transition == 1'b1) ? i_input_data[888 % IN_WIDTH] : ping_storage_data_11 ^ i_input_data[888 % IN_WIDTH];
                default: ping_storage_data_11 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_11;
                endcase
            end else begin
                case (input_count)
                109 / IN_WIDTH: pong_storage_data_11 <= (fillup_transition == 1'b1) ? i_input_data[109 % IN_WIDTH] : pong_storage_data_11 ^ i_input_data[109 % IN_WIDTH];
                226 / IN_WIDTH: pong_storage_data_11 <= (fillup_transition == 1'b1) ? i_input_data[226 % IN_WIDTH] : pong_storage_data_11 ^ i_input_data[226 % IN_WIDTH];
                820 / IN_WIDTH: pong_storage_data_11 <= (fillup_transition == 1'b1) ? i_input_data[820 % IN_WIDTH] : pong_storage_data_11 ^ i_input_data[820 % IN_WIDTH];
                888 / IN_WIDTH: pong_storage_data_11 <= (fillup_transition == 1'b1) ? i_input_data[888 % IN_WIDTH] : pong_storage_data_11 ^ i_input_data[888 % IN_WIDTH];
                default: pong_storage_data_11 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_11;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_11 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_11;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_11 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_11;
            end
        end
    end
end

logic ping_storage_data_12;
logic pong_storage_data_12;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_12 <= 1'b0;
        pong_storage_data_12 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                110 / IN_WIDTH: ping_storage_data_12 <= (fillup_transition == 1'b1) ? i_input_data[110 % IN_WIDTH] : ping_storage_data_12 ^ i_input_data[110 % IN_WIDTH];
                227 / IN_WIDTH: ping_storage_data_12 <= (fillup_transition == 1'b1) ? i_input_data[227 % IN_WIDTH] : ping_storage_data_12 ^ i_input_data[227 % IN_WIDTH];
                821 / IN_WIDTH: ping_storage_data_12 <= (fillup_transition == 1'b1) ? i_input_data[821 % IN_WIDTH] : ping_storage_data_12 ^ i_input_data[821 % IN_WIDTH];
                889 / IN_WIDTH: ping_storage_data_12 <= (fillup_transition == 1'b1) ? i_input_data[889 % IN_WIDTH] : ping_storage_data_12 ^ i_input_data[889 % IN_WIDTH];
                default: ping_storage_data_12 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_12;
                endcase
            end else begin
                case (input_count)
                110 / IN_WIDTH: pong_storage_data_12 <= (fillup_transition == 1'b1) ? i_input_data[110 % IN_WIDTH] : pong_storage_data_12 ^ i_input_data[110 % IN_WIDTH];
                227 / IN_WIDTH: pong_storage_data_12 <= (fillup_transition == 1'b1) ? i_input_data[227 % IN_WIDTH] : pong_storage_data_12 ^ i_input_data[227 % IN_WIDTH];
                821 / IN_WIDTH: pong_storage_data_12 <= (fillup_transition == 1'b1) ? i_input_data[821 % IN_WIDTH] : pong_storage_data_12 ^ i_input_data[821 % IN_WIDTH];
                889 / IN_WIDTH: pong_storage_data_12 <= (fillup_transition == 1'b1) ? i_input_data[889 % IN_WIDTH] : pong_storage_data_12 ^ i_input_data[889 % IN_WIDTH];
                default: pong_storage_data_12 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_12;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_12 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_12;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_12 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_12;
            end
        end
    end
end

logic ping_storage_data_13;
logic pong_storage_data_13;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_13 <= 1'b0;
        pong_storage_data_13 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                111 / IN_WIDTH: ping_storage_data_13 <= (fillup_transition == 1'b1) ? i_input_data[111 % IN_WIDTH] : ping_storage_data_13 ^ i_input_data[111 % IN_WIDTH];
                228 / IN_WIDTH: ping_storage_data_13 <= (fillup_transition == 1'b1) ? i_input_data[228 % IN_WIDTH] : ping_storage_data_13 ^ i_input_data[228 % IN_WIDTH];
                822 / IN_WIDTH: ping_storage_data_13 <= (fillup_transition == 1'b1) ? i_input_data[822 % IN_WIDTH] : ping_storage_data_13 ^ i_input_data[822 % IN_WIDTH];
                890 / IN_WIDTH: ping_storage_data_13 <= (fillup_transition == 1'b1) ? i_input_data[890 % IN_WIDTH] : ping_storage_data_13 ^ i_input_data[890 % IN_WIDTH];
                default: ping_storage_data_13 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_13;
                endcase
            end else begin
                case (input_count)
                111 / IN_WIDTH: pong_storage_data_13 <= (fillup_transition == 1'b1) ? i_input_data[111 % IN_WIDTH] : pong_storage_data_13 ^ i_input_data[111 % IN_WIDTH];
                228 / IN_WIDTH: pong_storage_data_13 <= (fillup_transition == 1'b1) ? i_input_data[228 % IN_WIDTH] : pong_storage_data_13 ^ i_input_data[228 % IN_WIDTH];
                822 / IN_WIDTH: pong_storage_data_13 <= (fillup_transition == 1'b1) ? i_input_data[822 % IN_WIDTH] : pong_storage_data_13 ^ i_input_data[822 % IN_WIDTH];
                890 / IN_WIDTH: pong_storage_data_13 <= (fillup_transition == 1'b1) ? i_input_data[890 % IN_WIDTH] : pong_storage_data_13 ^ i_input_data[890 % IN_WIDTH];
                default: pong_storage_data_13 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_13;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_13 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_13;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_13 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_13;
            end
        end
    end
end

logic ping_storage_data_14;
logic pong_storage_data_14;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_14 <= 1'b0;
        pong_storage_data_14 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                112 / IN_WIDTH: ping_storage_data_14 <= (fillup_transition == 1'b1) ? i_input_data[112 % IN_WIDTH] : ping_storage_data_14 ^ i_input_data[112 % IN_WIDTH];
                229 / IN_WIDTH: ping_storage_data_14 <= (fillup_transition == 1'b1) ? i_input_data[229 % IN_WIDTH] : ping_storage_data_14 ^ i_input_data[229 % IN_WIDTH];
                823 / IN_WIDTH: ping_storage_data_14 <= (fillup_transition == 1'b1) ? i_input_data[823 % IN_WIDTH] : ping_storage_data_14 ^ i_input_data[823 % IN_WIDTH];
                891 / IN_WIDTH: ping_storage_data_14 <= (fillup_transition == 1'b1) ? i_input_data[891 % IN_WIDTH] : ping_storage_data_14 ^ i_input_data[891 % IN_WIDTH];
                default: ping_storage_data_14 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_14;
                endcase
            end else begin
                case (input_count)
                112 / IN_WIDTH: pong_storage_data_14 <= (fillup_transition == 1'b1) ? i_input_data[112 % IN_WIDTH] : pong_storage_data_14 ^ i_input_data[112 % IN_WIDTH];
                229 / IN_WIDTH: pong_storage_data_14 <= (fillup_transition == 1'b1) ? i_input_data[229 % IN_WIDTH] : pong_storage_data_14 ^ i_input_data[229 % IN_WIDTH];
                823 / IN_WIDTH: pong_storage_data_14 <= (fillup_transition == 1'b1) ? i_input_data[823 % IN_WIDTH] : pong_storage_data_14 ^ i_input_data[823 % IN_WIDTH];
                891 / IN_WIDTH: pong_storage_data_14 <= (fillup_transition == 1'b1) ? i_input_data[891 % IN_WIDTH] : pong_storage_data_14 ^ i_input_data[891 % IN_WIDTH];
                default: pong_storage_data_14 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_14;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_14 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_14;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_14 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_14;
            end
        end
    end
end

logic ping_storage_data_15;
logic pong_storage_data_15;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_15 <= 1'b0;
        pong_storage_data_15 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                113 / IN_WIDTH: ping_storage_data_15 <= (fillup_transition == 1'b1) ? i_input_data[113 % IN_WIDTH] : ping_storage_data_15 ^ i_input_data[113 % IN_WIDTH];
                230 / IN_WIDTH: ping_storage_data_15 <= (fillup_transition == 1'b1) ? i_input_data[230 % IN_WIDTH] : ping_storage_data_15 ^ i_input_data[230 % IN_WIDTH];
                824 / IN_WIDTH: ping_storage_data_15 <= (fillup_transition == 1'b1) ? i_input_data[824 % IN_WIDTH] : ping_storage_data_15 ^ i_input_data[824 % IN_WIDTH];
                892 / IN_WIDTH: ping_storage_data_15 <= (fillup_transition == 1'b1) ? i_input_data[892 % IN_WIDTH] : ping_storage_data_15 ^ i_input_data[892 % IN_WIDTH];
                default: ping_storage_data_15 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_15;
                endcase
            end else begin
                case (input_count)
                113 / IN_WIDTH: pong_storage_data_15 <= (fillup_transition == 1'b1) ? i_input_data[113 % IN_WIDTH] : pong_storage_data_15 ^ i_input_data[113 % IN_WIDTH];
                230 / IN_WIDTH: pong_storage_data_15 <= (fillup_transition == 1'b1) ? i_input_data[230 % IN_WIDTH] : pong_storage_data_15 ^ i_input_data[230 % IN_WIDTH];
                824 / IN_WIDTH: pong_storage_data_15 <= (fillup_transition == 1'b1) ? i_input_data[824 % IN_WIDTH] : pong_storage_data_15 ^ i_input_data[824 % IN_WIDTH];
                892 / IN_WIDTH: pong_storage_data_15 <= (fillup_transition == 1'b1) ? i_input_data[892 % IN_WIDTH] : pong_storage_data_15 ^ i_input_data[892 % IN_WIDTH];
                default: pong_storage_data_15 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_15;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_15 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_15;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_15 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_15;
            end
        end
    end
end

logic ping_storage_data_16;
logic pong_storage_data_16;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_16 <= 1'b0;
        pong_storage_data_16 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                114 / IN_WIDTH: ping_storage_data_16 <= (fillup_transition == 1'b1) ? i_input_data[114 % IN_WIDTH] : ping_storage_data_16 ^ i_input_data[114 % IN_WIDTH];
                231 / IN_WIDTH: ping_storage_data_16 <= (fillup_transition == 1'b1) ? i_input_data[231 % IN_WIDTH] : ping_storage_data_16 ^ i_input_data[231 % IN_WIDTH];
                825 / IN_WIDTH: ping_storage_data_16 <= (fillup_transition == 1'b1) ? i_input_data[825 % IN_WIDTH] : ping_storage_data_16 ^ i_input_data[825 % IN_WIDTH];
                893 / IN_WIDTH: ping_storage_data_16 <= (fillup_transition == 1'b1) ? i_input_data[893 % IN_WIDTH] : ping_storage_data_16 ^ i_input_data[893 % IN_WIDTH];
                default: ping_storage_data_16 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_16;
                endcase
            end else begin
                case (input_count)
                114 / IN_WIDTH: pong_storage_data_16 <= (fillup_transition == 1'b1) ? i_input_data[114 % IN_WIDTH] : pong_storage_data_16 ^ i_input_data[114 % IN_WIDTH];
                231 / IN_WIDTH: pong_storage_data_16 <= (fillup_transition == 1'b1) ? i_input_data[231 % IN_WIDTH] : pong_storage_data_16 ^ i_input_data[231 % IN_WIDTH];
                825 / IN_WIDTH: pong_storage_data_16 <= (fillup_transition == 1'b1) ? i_input_data[825 % IN_WIDTH] : pong_storage_data_16 ^ i_input_data[825 % IN_WIDTH];
                893 / IN_WIDTH: pong_storage_data_16 <= (fillup_transition == 1'b1) ? i_input_data[893 % IN_WIDTH] : pong_storage_data_16 ^ i_input_data[893 % IN_WIDTH];
                default: pong_storage_data_16 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_16;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_16 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_16;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_16 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_16;
            end
        end
    end
end

logic ping_storage_data_17;
logic pong_storage_data_17;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_17 <= 1'b0;
        pong_storage_data_17 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                115 / IN_WIDTH: ping_storage_data_17 <= (fillup_transition == 1'b1) ? i_input_data[115 % IN_WIDTH] : ping_storage_data_17 ^ i_input_data[115 % IN_WIDTH];
                232 / IN_WIDTH: ping_storage_data_17 <= (fillup_transition == 1'b1) ? i_input_data[232 % IN_WIDTH] : ping_storage_data_17 ^ i_input_data[232 % IN_WIDTH];
                826 / IN_WIDTH: ping_storage_data_17 <= (fillup_transition == 1'b1) ? i_input_data[826 % IN_WIDTH] : ping_storage_data_17 ^ i_input_data[826 % IN_WIDTH];
                894 / IN_WIDTH: ping_storage_data_17 <= (fillup_transition == 1'b1) ? i_input_data[894 % IN_WIDTH] : ping_storage_data_17 ^ i_input_data[894 % IN_WIDTH];
                default: ping_storage_data_17 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_17;
                endcase
            end else begin
                case (input_count)
                115 / IN_WIDTH: pong_storage_data_17 <= (fillup_transition == 1'b1) ? i_input_data[115 % IN_WIDTH] : pong_storage_data_17 ^ i_input_data[115 % IN_WIDTH];
                232 / IN_WIDTH: pong_storage_data_17 <= (fillup_transition == 1'b1) ? i_input_data[232 % IN_WIDTH] : pong_storage_data_17 ^ i_input_data[232 % IN_WIDTH];
                826 / IN_WIDTH: pong_storage_data_17 <= (fillup_transition == 1'b1) ? i_input_data[826 % IN_WIDTH] : pong_storage_data_17 ^ i_input_data[826 % IN_WIDTH];
                894 / IN_WIDTH: pong_storage_data_17 <= (fillup_transition == 1'b1) ? i_input_data[894 % IN_WIDTH] : pong_storage_data_17 ^ i_input_data[894 % IN_WIDTH];
                default: pong_storage_data_17 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_17;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_17 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_17;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_17 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_17;
            end
        end
    end
end

logic ping_storage_data_18;
logic pong_storage_data_18;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_18 <= 1'b0;
        pong_storage_data_18 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                116 / IN_WIDTH: ping_storage_data_18 <= (fillup_transition == 1'b1) ? i_input_data[116 % IN_WIDTH] : ping_storage_data_18 ^ i_input_data[116 % IN_WIDTH];
                233 / IN_WIDTH: ping_storage_data_18 <= (fillup_transition == 1'b1) ? i_input_data[233 % IN_WIDTH] : ping_storage_data_18 ^ i_input_data[233 % IN_WIDTH];
                827 / IN_WIDTH: ping_storage_data_18 <= (fillup_transition == 1'b1) ? i_input_data[827 % IN_WIDTH] : ping_storage_data_18 ^ i_input_data[827 % IN_WIDTH];
                895 / IN_WIDTH: ping_storage_data_18 <= (fillup_transition == 1'b1) ? i_input_data[895 % IN_WIDTH] : ping_storage_data_18 ^ i_input_data[895 % IN_WIDTH];
                default: ping_storage_data_18 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_18;
                endcase
            end else begin
                case (input_count)
                116 / IN_WIDTH: pong_storage_data_18 <= (fillup_transition == 1'b1) ? i_input_data[116 % IN_WIDTH] : pong_storage_data_18 ^ i_input_data[116 % IN_WIDTH];
                233 / IN_WIDTH: pong_storage_data_18 <= (fillup_transition == 1'b1) ? i_input_data[233 % IN_WIDTH] : pong_storage_data_18 ^ i_input_data[233 % IN_WIDTH];
                827 / IN_WIDTH: pong_storage_data_18 <= (fillup_transition == 1'b1) ? i_input_data[827 % IN_WIDTH] : pong_storage_data_18 ^ i_input_data[827 % IN_WIDTH];
                895 / IN_WIDTH: pong_storage_data_18 <= (fillup_transition == 1'b1) ? i_input_data[895 % IN_WIDTH] : pong_storage_data_18 ^ i_input_data[895 % IN_WIDTH];
                default: pong_storage_data_18 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_18;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_18 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_18;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_18 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_18;
            end
        end
    end
end

logic ping_storage_data_19;
logic pong_storage_data_19;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_19 <= 1'b0;
        pong_storage_data_19 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                117 / IN_WIDTH: ping_storage_data_19 <= (fillup_transition == 1'b1) ? i_input_data[117 % IN_WIDTH] : ping_storage_data_19 ^ i_input_data[117 % IN_WIDTH];
                234 / IN_WIDTH: ping_storage_data_19 <= (fillup_transition == 1'b1) ? i_input_data[234 % IN_WIDTH] : ping_storage_data_19 ^ i_input_data[234 % IN_WIDTH];
                828 / IN_WIDTH: ping_storage_data_19 <= (fillup_transition == 1'b1) ? i_input_data[828 % IN_WIDTH] : ping_storage_data_19 ^ i_input_data[828 % IN_WIDTH];
                896 / IN_WIDTH: ping_storage_data_19 <= (fillup_transition == 1'b1) ? i_input_data[896 % IN_WIDTH] : ping_storage_data_19 ^ i_input_data[896 % IN_WIDTH];
                default: ping_storage_data_19 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_19;
                endcase
            end else begin
                case (input_count)
                117 / IN_WIDTH: pong_storage_data_19 <= (fillup_transition == 1'b1) ? i_input_data[117 % IN_WIDTH] : pong_storage_data_19 ^ i_input_data[117 % IN_WIDTH];
                234 / IN_WIDTH: pong_storage_data_19 <= (fillup_transition == 1'b1) ? i_input_data[234 % IN_WIDTH] : pong_storage_data_19 ^ i_input_data[234 % IN_WIDTH];
                828 / IN_WIDTH: pong_storage_data_19 <= (fillup_transition == 1'b1) ? i_input_data[828 % IN_WIDTH] : pong_storage_data_19 ^ i_input_data[828 % IN_WIDTH];
                896 / IN_WIDTH: pong_storage_data_19 <= (fillup_transition == 1'b1) ? i_input_data[896 % IN_WIDTH] : pong_storage_data_19 ^ i_input_data[896 % IN_WIDTH];
                default: pong_storage_data_19 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_19;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_19 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_19;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_19 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_19;
            end
        end
    end
end

logic ping_storage_data_20;
logic pong_storage_data_20;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_20 <= 1'b0;
        pong_storage_data_20 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                118 / IN_WIDTH: ping_storage_data_20 <= (fillup_transition == 1'b1) ? i_input_data[118 % IN_WIDTH] : ping_storage_data_20 ^ i_input_data[118 % IN_WIDTH];
                235 / IN_WIDTH: ping_storage_data_20 <= (fillup_transition == 1'b1) ? i_input_data[235 % IN_WIDTH] : ping_storage_data_20 ^ i_input_data[235 % IN_WIDTH];
                829 / IN_WIDTH: ping_storage_data_20 <= (fillup_transition == 1'b1) ? i_input_data[829 % IN_WIDTH] : ping_storage_data_20 ^ i_input_data[829 % IN_WIDTH];
                897 / IN_WIDTH: ping_storage_data_20 <= (fillup_transition == 1'b1) ? i_input_data[897 % IN_WIDTH] : ping_storage_data_20 ^ i_input_data[897 % IN_WIDTH];
                default: ping_storage_data_20 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_20;
                endcase
            end else begin
                case (input_count)
                118 / IN_WIDTH: pong_storage_data_20 <= (fillup_transition == 1'b1) ? i_input_data[118 % IN_WIDTH] : pong_storage_data_20 ^ i_input_data[118 % IN_WIDTH];
                235 / IN_WIDTH: pong_storage_data_20 <= (fillup_transition == 1'b1) ? i_input_data[235 % IN_WIDTH] : pong_storage_data_20 ^ i_input_data[235 % IN_WIDTH];
                829 / IN_WIDTH: pong_storage_data_20 <= (fillup_transition == 1'b1) ? i_input_data[829 % IN_WIDTH] : pong_storage_data_20 ^ i_input_data[829 % IN_WIDTH];
                897 / IN_WIDTH: pong_storage_data_20 <= (fillup_transition == 1'b1) ? i_input_data[897 % IN_WIDTH] : pong_storage_data_20 ^ i_input_data[897 % IN_WIDTH];
                default: pong_storage_data_20 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_20;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_20 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_20;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_20 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_20;
            end
        end
    end
end

logic ping_storage_data_21;
logic pong_storage_data_21;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_21 <= 1'b0;
        pong_storage_data_21 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                119 / IN_WIDTH: ping_storage_data_21 <= (fillup_transition == 1'b1) ? i_input_data[119 % IN_WIDTH] : ping_storage_data_21 ^ i_input_data[119 % IN_WIDTH];
                236 / IN_WIDTH: ping_storage_data_21 <= (fillup_transition == 1'b1) ? i_input_data[236 % IN_WIDTH] : ping_storage_data_21 ^ i_input_data[236 % IN_WIDTH];
                830 / IN_WIDTH: ping_storage_data_21 <= (fillup_transition == 1'b1) ? i_input_data[830 % IN_WIDTH] : ping_storage_data_21 ^ i_input_data[830 % IN_WIDTH];
                898 / IN_WIDTH: ping_storage_data_21 <= (fillup_transition == 1'b1) ? i_input_data[898 % IN_WIDTH] : ping_storage_data_21 ^ i_input_data[898 % IN_WIDTH];
                default: ping_storage_data_21 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_21;
                endcase
            end else begin
                case (input_count)
                119 / IN_WIDTH: pong_storage_data_21 <= (fillup_transition == 1'b1) ? i_input_data[119 % IN_WIDTH] : pong_storage_data_21 ^ i_input_data[119 % IN_WIDTH];
                236 / IN_WIDTH: pong_storage_data_21 <= (fillup_transition == 1'b1) ? i_input_data[236 % IN_WIDTH] : pong_storage_data_21 ^ i_input_data[236 % IN_WIDTH];
                830 / IN_WIDTH: pong_storage_data_21 <= (fillup_transition == 1'b1) ? i_input_data[830 % IN_WIDTH] : pong_storage_data_21 ^ i_input_data[830 % IN_WIDTH];
                898 / IN_WIDTH: pong_storage_data_21 <= (fillup_transition == 1'b1) ? i_input_data[898 % IN_WIDTH] : pong_storage_data_21 ^ i_input_data[898 % IN_WIDTH];
                default: pong_storage_data_21 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_21;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_21 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_21;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_21 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_21;
            end
        end
    end
end

logic ping_storage_data_22;
logic pong_storage_data_22;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_22 <= 1'b0;
        pong_storage_data_22 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                120 / IN_WIDTH: ping_storage_data_22 <= (fillup_transition == 1'b1) ? i_input_data[120 % IN_WIDTH] : ping_storage_data_22 ^ i_input_data[120 % IN_WIDTH];
                237 / IN_WIDTH: ping_storage_data_22 <= (fillup_transition == 1'b1) ? i_input_data[237 % IN_WIDTH] : ping_storage_data_22 ^ i_input_data[237 % IN_WIDTH];
                831 / IN_WIDTH: ping_storage_data_22 <= (fillup_transition == 1'b1) ? i_input_data[831 % IN_WIDTH] : ping_storage_data_22 ^ i_input_data[831 % IN_WIDTH];
                899 / IN_WIDTH: ping_storage_data_22 <= (fillup_transition == 1'b1) ? i_input_data[899 % IN_WIDTH] : ping_storage_data_22 ^ i_input_data[899 % IN_WIDTH];
                default: ping_storage_data_22 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_22;
                endcase
            end else begin
                case (input_count)
                120 / IN_WIDTH: pong_storage_data_22 <= (fillup_transition == 1'b1) ? i_input_data[120 % IN_WIDTH] : pong_storage_data_22 ^ i_input_data[120 % IN_WIDTH];
                237 / IN_WIDTH: pong_storage_data_22 <= (fillup_transition == 1'b1) ? i_input_data[237 % IN_WIDTH] : pong_storage_data_22 ^ i_input_data[237 % IN_WIDTH];
                831 / IN_WIDTH: pong_storage_data_22 <= (fillup_transition == 1'b1) ? i_input_data[831 % IN_WIDTH] : pong_storage_data_22 ^ i_input_data[831 % IN_WIDTH];
                899 / IN_WIDTH: pong_storage_data_22 <= (fillup_transition == 1'b1) ? i_input_data[899 % IN_WIDTH] : pong_storage_data_22 ^ i_input_data[899 % IN_WIDTH];
                default: pong_storage_data_22 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_22;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_22 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_22;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_22 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_22;
            end
        end
    end
end

logic ping_storage_data_23;
logic pong_storage_data_23;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_23 <= 1'b0;
        pong_storage_data_23 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                121 / IN_WIDTH: ping_storage_data_23 <= (fillup_transition == 1'b1) ? i_input_data[121 % IN_WIDTH] : ping_storage_data_23 ^ i_input_data[121 % IN_WIDTH];
                238 / IN_WIDTH: ping_storage_data_23 <= (fillup_transition == 1'b1) ? i_input_data[238 % IN_WIDTH] : ping_storage_data_23 ^ i_input_data[238 % IN_WIDTH];
                832 / IN_WIDTH: ping_storage_data_23 <= (fillup_transition == 1'b1) ? i_input_data[832 % IN_WIDTH] : ping_storage_data_23 ^ i_input_data[832 % IN_WIDTH];
                900 / IN_WIDTH: ping_storage_data_23 <= (fillup_transition == 1'b1) ? i_input_data[900 % IN_WIDTH] : ping_storage_data_23 ^ i_input_data[900 % IN_WIDTH];
                default: ping_storage_data_23 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_23;
                endcase
            end else begin
                case (input_count)
                121 / IN_WIDTH: pong_storage_data_23 <= (fillup_transition == 1'b1) ? i_input_data[121 % IN_WIDTH] : pong_storage_data_23 ^ i_input_data[121 % IN_WIDTH];
                238 / IN_WIDTH: pong_storage_data_23 <= (fillup_transition == 1'b1) ? i_input_data[238 % IN_WIDTH] : pong_storage_data_23 ^ i_input_data[238 % IN_WIDTH];
                832 / IN_WIDTH: pong_storage_data_23 <= (fillup_transition == 1'b1) ? i_input_data[832 % IN_WIDTH] : pong_storage_data_23 ^ i_input_data[832 % IN_WIDTH];
                900 / IN_WIDTH: pong_storage_data_23 <= (fillup_transition == 1'b1) ? i_input_data[900 % IN_WIDTH] : pong_storage_data_23 ^ i_input_data[900 % IN_WIDTH];
                default: pong_storage_data_23 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_23;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_23 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_23;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_23 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_23;
            end
        end
    end
end

logic ping_storage_data_24;
logic pong_storage_data_24;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_24 <= 1'b0;
        pong_storage_data_24 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                122 / IN_WIDTH: ping_storage_data_24 <= (fillup_transition == 1'b1) ? i_input_data[122 % IN_WIDTH] : ping_storage_data_24 ^ i_input_data[122 % IN_WIDTH];
                239 / IN_WIDTH: ping_storage_data_24 <= (fillup_transition == 1'b1) ? i_input_data[239 % IN_WIDTH] : ping_storage_data_24 ^ i_input_data[239 % IN_WIDTH];
                833 / IN_WIDTH: ping_storage_data_24 <= (fillup_transition == 1'b1) ? i_input_data[833 % IN_WIDTH] : ping_storage_data_24 ^ i_input_data[833 % IN_WIDTH];
                901 / IN_WIDTH: ping_storage_data_24 <= (fillup_transition == 1'b1) ? i_input_data[901 % IN_WIDTH] : ping_storage_data_24 ^ i_input_data[901 % IN_WIDTH];
                default: ping_storage_data_24 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_24;
                endcase
            end else begin
                case (input_count)
                122 / IN_WIDTH: pong_storage_data_24 <= (fillup_transition == 1'b1) ? i_input_data[122 % IN_WIDTH] : pong_storage_data_24 ^ i_input_data[122 % IN_WIDTH];
                239 / IN_WIDTH: pong_storage_data_24 <= (fillup_transition == 1'b1) ? i_input_data[239 % IN_WIDTH] : pong_storage_data_24 ^ i_input_data[239 % IN_WIDTH];
                833 / IN_WIDTH: pong_storage_data_24 <= (fillup_transition == 1'b1) ? i_input_data[833 % IN_WIDTH] : pong_storage_data_24 ^ i_input_data[833 % IN_WIDTH];
                901 / IN_WIDTH: pong_storage_data_24 <= (fillup_transition == 1'b1) ? i_input_data[901 % IN_WIDTH] : pong_storage_data_24 ^ i_input_data[901 % IN_WIDTH];
                default: pong_storage_data_24 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_24;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_24 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_24;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_24 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_24;
            end
        end
    end
end

logic ping_storage_data_25;
logic pong_storage_data_25;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_25 <= 1'b0;
        pong_storage_data_25 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                123 / IN_WIDTH: ping_storage_data_25 <= (fillup_transition == 1'b1) ? i_input_data[123 % IN_WIDTH] : ping_storage_data_25 ^ i_input_data[123 % IN_WIDTH];
                240 / IN_WIDTH: ping_storage_data_25 <= (fillup_transition == 1'b1) ? i_input_data[240 % IN_WIDTH] : ping_storage_data_25 ^ i_input_data[240 % IN_WIDTH];
                834 / IN_WIDTH: ping_storage_data_25 <= (fillup_transition == 1'b1) ? i_input_data[834 % IN_WIDTH] : ping_storage_data_25 ^ i_input_data[834 % IN_WIDTH];
                902 / IN_WIDTH: ping_storage_data_25 <= (fillup_transition == 1'b1) ? i_input_data[902 % IN_WIDTH] : ping_storage_data_25 ^ i_input_data[902 % IN_WIDTH];
                default: ping_storage_data_25 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_25;
                endcase
            end else begin
                case (input_count)
                123 / IN_WIDTH: pong_storage_data_25 <= (fillup_transition == 1'b1) ? i_input_data[123 % IN_WIDTH] : pong_storage_data_25 ^ i_input_data[123 % IN_WIDTH];
                240 / IN_WIDTH: pong_storage_data_25 <= (fillup_transition == 1'b1) ? i_input_data[240 % IN_WIDTH] : pong_storage_data_25 ^ i_input_data[240 % IN_WIDTH];
                834 / IN_WIDTH: pong_storage_data_25 <= (fillup_transition == 1'b1) ? i_input_data[834 % IN_WIDTH] : pong_storage_data_25 ^ i_input_data[834 % IN_WIDTH];
                902 / IN_WIDTH: pong_storage_data_25 <= (fillup_transition == 1'b1) ? i_input_data[902 % IN_WIDTH] : pong_storage_data_25 ^ i_input_data[902 % IN_WIDTH];
                default: pong_storage_data_25 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_25;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_25 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_25;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_25 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_25;
            end
        end
    end
end

logic ping_storage_data_26;
logic pong_storage_data_26;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_26 <= 1'b0;
        pong_storage_data_26 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                124 / IN_WIDTH: ping_storage_data_26 <= (fillup_transition == 1'b1) ? i_input_data[124 % IN_WIDTH] : ping_storage_data_26 ^ i_input_data[124 % IN_WIDTH];
                241 / IN_WIDTH: ping_storage_data_26 <= (fillup_transition == 1'b1) ? i_input_data[241 % IN_WIDTH] : ping_storage_data_26 ^ i_input_data[241 % IN_WIDTH];
                835 / IN_WIDTH: ping_storage_data_26 <= (fillup_transition == 1'b1) ? i_input_data[835 % IN_WIDTH] : ping_storage_data_26 ^ i_input_data[835 % IN_WIDTH];
                903 / IN_WIDTH: ping_storage_data_26 <= (fillup_transition == 1'b1) ? i_input_data[903 % IN_WIDTH] : ping_storage_data_26 ^ i_input_data[903 % IN_WIDTH];
                default: ping_storage_data_26 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_26;
                endcase
            end else begin
                case (input_count)
                124 / IN_WIDTH: pong_storage_data_26 <= (fillup_transition == 1'b1) ? i_input_data[124 % IN_WIDTH] : pong_storage_data_26 ^ i_input_data[124 % IN_WIDTH];
                241 / IN_WIDTH: pong_storage_data_26 <= (fillup_transition == 1'b1) ? i_input_data[241 % IN_WIDTH] : pong_storage_data_26 ^ i_input_data[241 % IN_WIDTH];
                835 / IN_WIDTH: pong_storage_data_26 <= (fillup_transition == 1'b1) ? i_input_data[835 % IN_WIDTH] : pong_storage_data_26 ^ i_input_data[835 % IN_WIDTH];
                903 / IN_WIDTH: pong_storage_data_26 <= (fillup_transition == 1'b1) ? i_input_data[903 % IN_WIDTH] : pong_storage_data_26 ^ i_input_data[903 % IN_WIDTH];
                default: pong_storage_data_26 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_26;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_26 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_26;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_26 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_26;
            end
        end
    end
end

logic ping_storage_data_27;
logic pong_storage_data_27;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_27 <= 1'b0;
        pong_storage_data_27 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                125 / IN_WIDTH: ping_storage_data_27 <= (fillup_transition == 1'b1) ? i_input_data[125 % IN_WIDTH] : ping_storage_data_27 ^ i_input_data[125 % IN_WIDTH];
                242 / IN_WIDTH: ping_storage_data_27 <= (fillup_transition == 1'b1) ? i_input_data[242 % IN_WIDTH] : ping_storage_data_27 ^ i_input_data[242 % IN_WIDTH];
                836 / IN_WIDTH: ping_storage_data_27 <= (fillup_transition == 1'b1) ? i_input_data[836 % IN_WIDTH] : ping_storage_data_27 ^ i_input_data[836 % IN_WIDTH];
                904 / IN_WIDTH: ping_storage_data_27 <= (fillup_transition == 1'b1) ? i_input_data[904 % IN_WIDTH] : ping_storage_data_27 ^ i_input_data[904 % IN_WIDTH];
                default: ping_storage_data_27 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_27;
                endcase
            end else begin
                case (input_count)
                125 / IN_WIDTH: pong_storage_data_27 <= (fillup_transition == 1'b1) ? i_input_data[125 % IN_WIDTH] : pong_storage_data_27 ^ i_input_data[125 % IN_WIDTH];
                242 / IN_WIDTH: pong_storage_data_27 <= (fillup_transition == 1'b1) ? i_input_data[242 % IN_WIDTH] : pong_storage_data_27 ^ i_input_data[242 % IN_WIDTH];
                836 / IN_WIDTH: pong_storage_data_27 <= (fillup_transition == 1'b1) ? i_input_data[836 % IN_WIDTH] : pong_storage_data_27 ^ i_input_data[836 % IN_WIDTH];
                904 / IN_WIDTH: pong_storage_data_27 <= (fillup_transition == 1'b1) ? i_input_data[904 % IN_WIDTH] : pong_storage_data_27 ^ i_input_data[904 % IN_WIDTH];
                default: pong_storage_data_27 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_27;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_27 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_27;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_27 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_27;
            end
        end
    end
end

logic ping_storage_data_28;
logic pong_storage_data_28;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_28 <= 1'b0;
        pong_storage_data_28 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                126 / IN_WIDTH: ping_storage_data_28 <= (fillup_transition == 1'b1) ? i_input_data[126 % IN_WIDTH] : ping_storage_data_28 ^ i_input_data[126 % IN_WIDTH];
                243 / IN_WIDTH: ping_storage_data_28 <= (fillup_transition == 1'b1) ? i_input_data[243 % IN_WIDTH] : ping_storage_data_28 ^ i_input_data[243 % IN_WIDTH];
                837 / IN_WIDTH: ping_storage_data_28 <= (fillup_transition == 1'b1) ? i_input_data[837 % IN_WIDTH] : ping_storage_data_28 ^ i_input_data[837 % IN_WIDTH];
                905 / IN_WIDTH: ping_storage_data_28 <= (fillup_transition == 1'b1) ? i_input_data[905 % IN_WIDTH] : ping_storage_data_28 ^ i_input_data[905 % IN_WIDTH];
                default: ping_storage_data_28 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_28;
                endcase
            end else begin
                case (input_count)
                126 / IN_WIDTH: pong_storage_data_28 <= (fillup_transition == 1'b1) ? i_input_data[126 % IN_WIDTH] : pong_storage_data_28 ^ i_input_data[126 % IN_WIDTH];
                243 / IN_WIDTH: pong_storage_data_28 <= (fillup_transition == 1'b1) ? i_input_data[243 % IN_WIDTH] : pong_storage_data_28 ^ i_input_data[243 % IN_WIDTH];
                837 / IN_WIDTH: pong_storage_data_28 <= (fillup_transition == 1'b1) ? i_input_data[837 % IN_WIDTH] : pong_storage_data_28 ^ i_input_data[837 % IN_WIDTH];
                905 / IN_WIDTH: pong_storage_data_28 <= (fillup_transition == 1'b1) ? i_input_data[905 % IN_WIDTH] : pong_storage_data_28 ^ i_input_data[905 % IN_WIDTH];
                default: pong_storage_data_28 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_28;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_28 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_28;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_28 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_28;
            end
        end
    end
end

logic ping_storage_data_29;
logic pong_storage_data_29;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_29 <= 1'b0;
        pong_storage_data_29 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                127 / IN_WIDTH: ping_storage_data_29 <= (fillup_transition == 1'b1) ? i_input_data[127 % IN_WIDTH] : ping_storage_data_29 ^ i_input_data[127 % IN_WIDTH];
                244 / IN_WIDTH: ping_storage_data_29 <= (fillup_transition == 1'b1) ? i_input_data[244 % IN_WIDTH] : ping_storage_data_29 ^ i_input_data[244 % IN_WIDTH];
                838 / IN_WIDTH: ping_storage_data_29 <= (fillup_transition == 1'b1) ? i_input_data[838 % IN_WIDTH] : ping_storage_data_29 ^ i_input_data[838 % IN_WIDTH];
                906 / IN_WIDTH: ping_storage_data_29 <= (fillup_transition == 1'b1) ? i_input_data[906 % IN_WIDTH] : ping_storage_data_29 ^ i_input_data[906 % IN_WIDTH];
                default: ping_storage_data_29 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_29;
                endcase
            end else begin
                case (input_count)
                127 / IN_WIDTH: pong_storage_data_29 <= (fillup_transition == 1'b1) ? i_input_data[127 % IN_WIDTH] : pong_storage_data_29 ^ i_input_data[127 % IN_WIDTH];
                244 / IN_WIDTH: pong_storage_data_29 <= (fillup_transition == 1'b1) ? i_input_data[244 % IN_WIDTH] : pong_storage_data_29 ^ i_input_data[244 % IN_WIDTH];
                838 / IN_WIDTH: pong_storage_data_29 <= (fillup_transition == 1'b1) ? i_input_data[838 % IN_WIDTH] : pong_storage_data_29 ^ i_input_data[838 % IN_WIDTH];
                906 / IN_WIDTH: pong_storage_data_29 <= (fillup_transition == 1'b1) ? i_input_data[906 % IN_WIDTH] : pong_storage_data_29 ^ i_input_data[906 % IN_WIDTH];
                default: pong_storage_data_29 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_29;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_29 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_29;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_29 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_29;
            end
        end
    end
end

logic ping_storage_data_30;
logic pong_storage_data_30;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_30 <= 1'b0;
        pong_storage_data_30 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                128 / IN_WIDTH: ping_storage_data_30 <= (fillup_transition == 1'b1) ? i_input_data[128 % IN_WIDTH] : ping_storage_data_30 ^ i_input_data[128 % IN_WIDTH];
                245 / IN_WIDTH: ping_storage_data_30 <= (fillup_transition == 1'b1) ? i_input_data[245 % IN_WIDTH] : ping_storage_data_30 ^ i_input_data[245 % IN_WIDTH];
                839 / IN_WIDTH: ping_storage_data_30 <= (fillup_transition == 1'b1) ? i_input_data[839 % IN_WIDTH] : ping_storage_data_30 ^ i_input_data[839 % IN_WIDTH];
                907 / IN_WIDTH: ping_storage_data_30 <= (fillup_transition == 1'b1) ? i_input_data[907 % IN_WIDTH] : ping_storage_data_30 ^ i_input_data[907 % IN_WIDTH];
                default: ping_storage_data_30 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_30;
                endcase
            end else begin
                case (input_count)
                128 / IN_WIDTH: pong_storage_data_30 <= (fillup_transition == 1'b1) ? i_input_data[128 % IN_WIDTH] : pong_storage_data_30 ^ i_input_data[128 % IN_WIDTH];
                245 / IN_WIDTH: pong_storage_data_30 <= (fillup_transition == 1'b1) ? i_input_data[245 % IN_WIDTH] : pong_storage_data_30 ^ i_input_data[245 % IN_WIDTH];
                839 / IN_WIDTH: pong_storage_data_30 <= (fillup_transition == 1'b1) ? i_input_data[839 % IN_WIDTH] : pong_storage_data_30 ^ i_input_data[839 % IN_WIDTH];
                907 / IN_WIDTH: pong_storage_data_30 <= (fillup_transition == 1'b1) ? i_input_data[907 % IN_WIDTH] : pong_storage_data_30 ^ i_input_data[907 % IN_WIDTH];
                default: pong_storage_data_30 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_30;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_30 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_30;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_30 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_30;
            end
        end
    end
end

logic ping_storage_data_31;
logic pong_storage_data_31;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_31 <= 1'b0;
        pong_storage_data_31 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                129 / IN_WIDTH: ping_storage_data_31 <= (fillup_transition == 1'b1) ? i_input_data[129 % IN_WIDTH] : ping_storage_data_31 ^ i_input_data[129 % IN_WIDTH];
                246 / IN_WIDTH: ping_storage_data_31 <= (fillup_transition == 1'b1) ? i_input_data[246 % IN_WIDTH] : ping_storage_data_31 ^ i_input_data[246 % IN_WIDTH];
                840 / IN_WIDTH: ping_storage_data_31 <= (fillup_transition == 1'b1) ? i_input_data[840 % IN_WIDTH] : ping_storage_data_31 ^ i_input_data[840 % IN_WIDTH];
                908 / IN_WIDTH: ping_storage_data_31 <= (fillup_transition == 1'b1) ? i_input_data[908 % IN_WIDTH] : ping_storage_data_31 ^ i_input_data[908 % IN_WIDTH];
                default: ping_storage_data_31 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_31;
                endcase
            end else begin
                case (input_count)
                129 / IN_WIDTH: pong_storage_data_31 <= (fillup_transition == 1'b1) ? i_input_data[129 % IN_WIDTH] : pong_storage_data_31 ^ i_input_data[129 % IN_WIDTH];
                246 / IN_WIDTH: pong_storage_data_31 <= (fillup_transition == 1'b1) ? i_input_data[246 % IN_WIDTH] : pong_storage_data_31 ^ i_input_data[246 % IN_WIDTH];
                840 / IN_WIDTH: pong_storage_data_31 <= (fillup_transition == 1'b1) ? i_input_data[840 % IN_WIDTH] : pong_storage_data_31 ^ i_input_data[840 % IN_WIDTH];
                908 / IN_WIDTH: pong_storage_data_31 <= (fillup_transition == 1'b1) ? i_input_data[908 % IN_WIDTH] : pong_storage_data_31 ^ i_input_data[908 % IN_WIDTH];
                default: pong_storage_data_31 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_31;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_31 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_31;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_31 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_31;
            end
        end
    end
end

logic ping_storage_data_32;
logic pong_storage_data_32;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_32 <= 1'b0;
        pong_storage_data_32 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                130 / IN_WIDTH: ping_storage_data_32 <= (fillup_transition == 1'b1) ? i_input_data[130 % IN_WIDTH] : ping_storage_data_32 ^ i_input_data[130 % IN_WIDTH];
                247 / IN_WIDTH: ping_storage_data_32 <= (fillup_transition == 1'b1) ? i_input_data[247 % IN_WIDTH] : ping_storage_data_32 ^ i_input_data[247 % IN_WIDTH];
                841 / IN_WIDTH: ping_storage_data_32 <= (fillup_transition == 1'b1) ? i_input_data[841 % IN_WIDTH] : ping_storage_data_32 ^ i_input_data[841 % IN_WIDTH];
                909 / IN_WIDTH: ping_storage_data_32 <= (fillup_transition == 1'b1) ? i_input_data[909 % IN_WIDTH] : ping_storage_data_32 ^ i_input_data[909 % IN_WIDTH];
                default: ping_storage_data_32 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_32;
                endcase
            end else begin
                case (input_count)
                130 / IN_WIDTH: pong_storage_data_32 <= (fillup_transition == 1'b1) ? i_input_data[130 % IN_WIDTH] : pong_storage_data_32 ^ i_input_data[130 % IN_WIDTH];
                247 / IN_WIDTH: pong_storage_data_32 <= (fillup_transition == 1'b1) ? i_input_data[247 % IN_WIDTH] : pong_storage_data_32 ^ i_input_data[247 % IN_WIDTH];
                841 / IN_WIDTH: pong_storage_data_32 <= (fillup_transition == 1'b1) ? i_input_data[841 % IN_WIDTH] : pong_storage_data_32 ^ i_input_data[841 % IN_WIDTH];
                909 / IN_WIDTH: pong_storage_data_32 <= (fillup_transition == 1'b1) ? i_input_data[909 % IN_WIDTH] : pong_storage_data_32 ^ i_input_data[909 % IN_WIDTH];
                default: pong_storage_data_32 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_32;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_32 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_32;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_32 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_32;
            end
        end
    end
end

logic ping_storage_data_33;
logic pong_storage_data_33;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_33 <= 1'b0;
        pong_storage_data_33 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                131 / IN_WIDTH: ping_storage_data_33 <= (fillup_transition == 1'b1) ? i_input_data[131 % IN_WIDTH] : ping_storage_data_33 ^ i_input_data[131 % IN_WIDTH];
                248 / IN_WIDTH: ping_storage_data_33 <= (fillup_transition == 1'b1) ? i_input_data[248 % IN_WIDTH] : ping_storage_data_33 ^ i_input_data[248 % IN_WIDTH];
                842 / IN_WIDTH: ping_storage_data_33 <= (fillup_transition == 1'b1) ? i_input_data[842 % IN_WIDTH] : ping_storage_data_33 ^ i_input_data[842 % IN_WIDTH];
                910 / IN_WIDTH: ping_storage_data_33 <= (fillup_transition == 1'b1) ? i_input_data[910 % IN_WIDTH] : ping_storage_data_33 ^ i_input_data[910 % IN_WIDTH];
                default: ping_storage_data_33 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_33;
                endcase
            end else begin
                case (input_count)
                131 / IN_WIDTH: pong_storage_data_33 <= (fillup_transition == 1'b1) ? i_input_data[131 % IN_WIDTH] : pong_storage_data_33 ^ i_input_data[131 % IN_WIDTH];
                248 / IN_WIDTH: pong_storage_data_33 <= (fillup_transition == 1'b1) ? i_input_data[248 % IN_WIDTH] : pong_storage_data_33 ^ i_input_data[248 % IN_WIDTH];
                842 / IN_WIDTH: pong_storage_data_33 <= (fillup_transition == 1'b1) ? i_input_data[842 % IN_WIDTH] : pong_storage_data_33 ^ i_input_data[842 % IN_WIDTH];
                910 / IN_WIDTH: pong_storage_data_33 <= (fillup_transition == 1'b1) ? i_input_data[910 % IN_WIDTH] : pong_storage_data_33 ^ i_input_data[910 % IN_WIDTH];
                default: pong_storage_data_33 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_33;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_33 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_33;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_33 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_33;
            end
        end
    end
end

logic ping_storage_data_34;
logic pong_storage_data_34;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_34 <= 1'b0;
        pong_storage_data_34 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                132 / IN_WIDTH: ping_storage_data_34 <= (fillup_transition == 1'b1) ? i_input_data[132 % IN_WIDTH] : ping_storage_data_34 ^ i_input_data[132 % IN_WIDTH];
                249 / IN_WIDTH: ping_storage_data_34 <= (fillup_transition == 1'b1) ? i_input_data[249 % IN_WIDTH] : ping_storage_data_34 ^ i_input_data[249 % IN_WIDTH];
                843 / IN_WIDTH: ping_storage_data_34 <= (fillup_transition == 1'b1) ? i_input_data[843 % IN_WIDTH] : ping_storage_data_34 ^ i_input_data[843 % IN_WIDTH];
                911 / IN_WIDTH: ping_storage_data_34 <= (fillup_transition == 1'b1) ? i_input_data[911 % IN_WIDTH] : ping_storage_data_34 ^ i_input_data[911 % IN_WIDTH];
                default: ping_storage_data_34 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_34;
                endcase
            end else begin
                case (input_count)
                132 / IN_WIDTH: pong_storage_data_34 <= (fillup_transition == 1'b1) ? i_input_data[132 % IN_WIDTH] : pong_storage_data_34 ^ i_input_data[132 % IN_WIDTH];
                249 / IN_WIDTH: pong_storage_data_34 <= (fillup_transition == 1'b1) ? i_input_data[249 % IN_WIDTH] : pong_storage_data_34 ^ i_input_data[249 % IN_WIDTH];
                843 / IN_WIDTH: pong_storage_data_34 <= (fillup_transition == 1'b1) ? i_input_data[843 % IN_WIDTH] : pong_storage_data_34 ^ i_input_data[843 % IN_WIDTH];
                911 / IN_WIDTH: pong_storage_data_34 <= (fillup_transition == 1'b1) ? i_input_data[911 % IN_WIDTH] : pong_storage_data_34 ^ i_input_data[911 % IN_WIDTH];
                default: pong_storage_data_34 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_34;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_34 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_34;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_34 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_34;
            end
        end
    end
end

logic ping_storage_data_35;
logic pong_storage_data_35;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_35 <= 1'b0;
        pong_storage_data_35 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                133 / IN_WIDTH: ping_storage_data_35 <= (fillup_transition == 1'b1) ? i_input_data[133 % IN_WIDTH] : ping_storage_data_35 ^ i_input_data[133 % IN_WIDTH];
                250 / IN_WIDTH: ping_storage_data_35 <= (fillup_transition == 1'b1) ? i_input_data[250 % IN_WIDTH] : ping_storage_data_35 ^ i_input_data[250 % IN_WIDTH];
                844 / IN_WIDTH: ping_storage_data_35 <= (fillup_transition == 1'b1) ? i_input_data[844 % IN_WIDTH] : ping_storage_data_35 ^ i_input_data[844 % IN_WIDTH];
                912 / IN_WIDTH: ping_storage_data_35 <= (fillup_transition == 1'b1) ? i_input_data[912 % IN_WIDTH] : ping_storage_data_35 ^ i_input_data[912 % IN_WIDTH];
                default: ping_storage_data_35 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_35;
                endcase
            end else begin
                case (input_count)
                133 / IN_WIDTH: pong_storage_data_35 <= (fillup_transition == 1'b1) ? i_input_data[133 % IN_WIDTH] : pong_storage_data_35 ^ i_input_data[133 % IN_WIDTH];
                250 / IN_WIDTH: pong_storage_data_35 <= (fillup_transition == 1'b1) ? i_input_data[250 % IN_WIDTH] : pong_storage_data_35 ^ i_input_data[250 % IN_WIDTH];
                844 / IN_WIDTH: pong_storage_data_35 <= (fillup_transition == 1'b1) ? i_input_data[844 % IN_WIDTH] : pong_storage_data_35 ^ i_input_data[844 % IN_WIDTH];
                912 / IN_WIDTH: pong_storage_data_35 <= (fillup_transition == 1'b1) ? i_input_data[912 % IN_WIDTH] : pong_storage_data_35 ^ i_input_data[912 % IN_WIDTH];
                default: pong_storage_data_35 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_35;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_35 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_35;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_35 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_35;
            end
        end
    end
end

logic ping_storage_data_36;
logic pong_storage_data_36;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_36 <= 1'b0;
        pong_storage_data_36 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                134 / IN_WIDTH: ping_storage_data_36 <= (fillup_transition == 1'b1) ? i_input_data[134 % IN_WIDTH] : ping_storage_data_36 ^ i_input_data[134 % IN_WIDTH];
                251 / IN_WIDTH: ping_storage_data_36 <= (fillup_transition == 1'b1) ? i_input_data[251 % IN_WIDTH] : ping_storage_data_36 ^ i_input_data[251 % IN_WIDTH];
                845 / IN_WIDTH: ping_storage_data_36 <= (fillup_transition == 1'b1) ? i_input_data[845 % IN_WIDTH] : ping_storage_data_36 ^ i_input_data[845 % IN_WIDTH];
                913 / IN_WIDTH: ping_storage_data_36 <= (fillup_transition == 1'b1) ? i_input_data[913 % IN_WIDTH] : ping_storage_data_36 ^ i_input_data[913 % IN_WIDTH];
                default: ping_storage_data_36 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_36;
                endcase
            end else begin
                case (input_count)
                134 / IN_WIDTH: pong_storage_data_36 <= (fillup_transition == 1'b1) ? i_input_data[134 % IN_WIDTH] : pong_storage_data_36 ^ i_input_data[134 % IN_WIDTH];
                251 / IN_WIDTH: pong_storage_data_36 <= (fillup_transition == 1'b1) ? i_input_data[251 % IN_WIDTH] : pong_storage_data_36 ^ i_input_data[251 % IN_WIDTH];
                845 / IN_WIDTH: pong_storage_data_36 <= (fillup_transition == 1'b1) ? i_input_data[845 % IN_WIDTH] : pong_storage_data_36 ^ i_input_data[845 % IN_WIDTH];
                913 / IN_WIDTH: pong_storage_data_36 <= (fillup_transition == 1'b1) ? i_input_data[913 % IN_WIDTH] : pong_storage_data_36 ^ i_input_data[913 % IN_WIDTH];
                default: pong_storage_data_36 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_36;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_36 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_36;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_36 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_36;
            end
        end
    end
end

logic ping_storage_data_37;
logic pong_storage_data_37;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_37 <= 1'b0;
        pong_storage_data_37 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                135 / IN_WIDTH: ping_storage_data_37 <= (fillup_transition == 1'b1) ? i_input_data[135 % IN_WIDTH] : ping_storage_data_37 ^ i_input_data[135 % IN_WIDTH];
                252 / IN_WIDTH: ping_storage_data_37 <= (fillup_transition == 1'b1) ? i_input_data[252 % IN_WIDTH] : ping_storage_data_37 ^ i_input_data[252 % IN_WIDTH];
                846 / IN_WIDTH: ping_storage_data_37 <= (fillup_transition == 1'b1) ? i_input_data[846 % IN_WIDTH] : ping_storage_data_37 ^ i_input_data[846 % IN_WIDTH];
                914 / IN_WIDTH: ping_storage_data_37 <= (fillup_transition == 1'b1) ? i_input_data[914 % IN_WIDTH] : ping_storage_data_37 ^ i_input_data[914 % IN_WIDTH];
                default: ping_storage_data_37 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_37;
                endcase
            end else begin
                case (input_count)
                135 / IN_WIDTH: pong_storage_data_37 <= (fillup_transition == 1'b1) ? i_input_data[135 % IN_WIDTH] : pong_storage_data_37 ^ i_input_data[135 % IN_WIDTH];
                252 / IN_WIDTH: pong_storage_data_37 <= (fillup_transition == 1'b1) ? i_input_data[252 % IN_WIDTH] : pong_storage_data_37 ^ i_input_data[252 % IN_WIDTH];
                846 / IN_WIDTH: pong_storage_data_37 <= (fillup_transition == 1'b1) ? i_input_data[846 % IN_WIDTH] : pong_storage_data_37 ^ i_input_data[846 % IN_WIDTH];
                914 / IN_WIDTH: pong_storage_data_37 <= (fillup_transition == 1'b1) ? i_input_data[914 % IN_WIDTH] : pong_storage_data_37 ^ i_input_data[914 % IN_WIDTH];
                default: pong_storage_data_37 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_37;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_37 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_37;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_37 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_37;
            end
        end
    end
end

logic ping_storage_data_38;
logic pong_storage_data_38;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_38 <= 1'b0;
        pong_storage_data_38 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                136 / IN_WIDTH: ping_storage_data_38 <= (fillup_transition == 1'b1) ? i_input_data[136 % IN_WIDTH] : ping_storage_data_38 ^ i_input_data[136 % IN_WIDTH];
                253 / IN_WIDTH: ping_storage_data_38 <= (fillup_transition == 1'b1) ? i_input_data[253 % IN_WIDTH] : ping_storage_data_38 ^ i_input_data[253 % IN_WIDTH];
                847 / IN_WIDTH: ping_storage_data_38 <= (fillup_transition == 1'b1) ? i_input_data[847 % IN_WIDTH] : ping_storage_data_38 ^ i_input_data[847 % IN_WIDTH];
                915 / IN_WIDTH: ping_storage_data_38 <= (fillup_transition == 1'b1) ? i_input_data[915 % IN_WIDTH] : ping_storage_data_38 ^ i_input_data[915 % IN_WIDTH];
                default: ping_storage_data_38 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_38;
                endcase
            end else begin
                case (input_count)
                136 / IN_WIDTH: pong_storage_data_38 <= (fillup_transition == 1'b1) ? i_input_data[136 % IN_WIDTH] : pong_storage_data_38 ^ i_input_data[136 % IN_WIDTH];
                253 / IN_WIDTH: pong_storage_data_38 <= (fillup_transition == 1'b1) ? i_input_data[253 % IN_WIDTH] : pong_storage_data_38 ^ i_input_data[253 % IN_WIDTH];
                847 / IN_WIDTH: pong_storage_data_38 <= (fillup_transition == 1'b1) ? i_input_data[847 % IN_WIDTH] : pong_storage_data_38 ^ i_input_data[847 % IN_WIDTH];
                915 / IN_WIDTH: pong_storage_data_38 <= (fillup_transition == 1'b1) ? i_input_data[915 % IN_WIDTH] : pong_storage_data_38 ^ i_input_data[915 % IN_WIDTH];
                default: pong_storage_data_38 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_38;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_38 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_38;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_38 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_38;
            end
        end
    end
end

logic ping_storage_data_39;
logic pong_storage_data_39;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_39 <= 1'b0;
        pong_storage_data_39 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                137 / IN_WIDTH: ping_storage_data_39 <= (fillup_transition == 1'b1) ? i_input_data[137 % IN_WIDTH] : ping_storage_data_39 ^ i_input_data[137 % IN_WIDTH];
                254 / IN_WIDTH: ping_storage_data_39 <= (fillup_transition == 1'b1) ? i_input_data[254 % IN_WIDTH] : ping_storage_data_39 ^ i_input_data[254 % IN_WIDTH];
                848 / IN_WIDTH: ping_storage_data_39 <= (fillup_transition == 1'b1) ? i_input_data[848 % IN_WIDTH] : ping_storage_data_39 ^ i_input_data[848 % IN_WIDTH];
                916 / IN_WIDTH: ping_storage_data_39 <= (fillup_transition == 1'b1) ? i_input_data[916 % IN_WIDTH] : ping_storage_data_39 ^ i_input_data[916 % IN_WIDTH];
                default: ping_storage_data_39 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_39;
                endcase
            end else begin
                case (input_count)
                137 / IN_WIDTH: pong_storage_data_39 <= (fillup_transition == 1'b1) ? i_input_data[137 % IN_WIDTH] : pong_storage_data_39 ^ i_input_data[137 % IN_WIDTH];
                254 / IN_WIDTH: pong_storage_data_39 <= (fillup_transition == 1'b1) ? i_input_data[254 % IN_WIDTH] : pong_storage_data_39 ^ i_input_data[254 % IN_WIDTH];
                848 / IN_WIDTH: pong_storage_data_39 <= (fillup_transition == 1'b1) ? i_input_data[848 % IN_WIDTH] : pong_storage_data_39 ^ i_input_data[848 % IN_WIDTH];
                916 / IN_WIDTH: pong_storage_data_39 <= (fillup_transition == 1'b1) ? i_input_data[916 % IN_WIDTH] : pong_storage_data_39 ^ i_input_data[916 % IN_WIDTH];
                default: pong_storage_data_39 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_39;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_39 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_39;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_39 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_39;
            end
        end
    end
end

logic ping_storage_data_40;
logic pong_storage_data_40;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_40 <= 1'b0;
        pong_storage_data_40 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                138 / IN_WIDTH: ping_storage_data_40 <= (fillup_transition == 1'b1) ? i_input_data[138 % IN_WIDTH] : ping_storage_data_40 ^ i_input_data[138 % IN_WIDTH];
                255 / IN_WIDTH: ping_storage_data_40 <= (fillup_transition == 1'b1) ? i_input_data[255 % IN_WIDTH] : ping_storage_data_40 ^ i_input_data[255 % IN_WIDTH];
                849 / IN_WIDTH: ping_storage_data_40 <= (fillup_transition == 1'b1) ? i_input_data[849 % IN_WIDTH] : ping_storage_data_40 ^ i_input_data[849 % IN_WIDTH];
                917 / IN_WIDTH: ping_storage_data_40 <= (fillup_transition == 1'b1) ? i_input_data[917 % IN_WIDTH] : ping_storage_data_40 ^ i_input_data[917 % IN_WIDTH];
                default: ping_storage_data_40 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_40;
                endcase
            end else begin
                case (input_count)
                138 / IN_WIDTH: pong_storage_data_40 <= (fillup_transition == 1'b1) ? i_input_data[138 % IN_WIDTH] : pong_storage_data_40 ^ i_input_data[138 % IN_WIDTH];
                255 / IN_WIDTH: pong_storage_data_40 <= (fillup_transition == 1'b1) ? i_input_data[255 % IN_WIDTH] : pong_storage_data_40 ^ i_input_data[255 % IN_WIDTH];
                849 / IN_WIDTH: pong_storage_data_40 <= (fillup_transition == 1'b1) ? i_input_data[849 % IN_WIDTH] : pong_storage_data_40 ^ i_input_data[849 % IN_WIDTH];
                917 / IN_WIDTH: pong_storage_data_40 <= (fillup_transition == 1'b1) ? i_input_data[917 % IN_WIDTH] : pong_storage_data_40 ^ i_input_data[917 % IN_WIDTH];
                default: pong_storage_data_40 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_40;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_40 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_40;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_40 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_40;
            end
        end
    end
end

logic ping_storage_data_41;
logic pong_storage_data_41;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_41 <= 1'b0;
        pong_storage_data_41 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                139 / IN_WIDTH: ping_storage_data_41 <= (fillup_transition == 1'b1) ? i_input_data[139 % IN_WIDTH] : ping_storage_data_41 ^ i_input_data[139 % IN_WIDTH];
                256 / IN_WIDTH: ping_storage_data_41 <= (fillup_transition == 1'b1) ? i_input_data[256 % IN_WIDTH] : ping_storage_data_41 ^ i_input_data[256 % IN_WIDTH];
                850 / IN_WIDTH: ping_storage_data_41 <= (fillup_transition == 1'b1) ? i_input_data[850 % IN_WIDTH] : ping_storage_data_41 ^ i_input_data[850 % IN_WIDTH];
                918 / IN_WIDTH: ping_storage_data_41 <= (fillup_transition == 1'b1) ? i_input_data[918 % IN_WIDTH] : ping_storage_data_41 ^ i_input_data[918 % IN_WIDTH];
                default: ping_storage_data_41 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_41;
                endcase
            end else begin
                case (input_count)
                139 / IN_WIDTH: pong_storage_data_41 <= (fillup_transition == 1'b1) ? i_input_data[139 % IN_WIDTH] : pong_storage_data_41 ^ i_input_data[139 % IN_WIDTH];
                256 / IN_WIDTH: pong_storage_data_41 <= (fillup_transition == 1'b1) ? i_input_data[256 % IN_WIDTH] : pong_storage_data_41 ^ i_input_data[256 % IN_WIDTH];
                850 / IN_WIDTH: pong_storage_data_41 <= (fillup_transition == 1'b1) ? i_input_data[850 % IN_WIDTH] : pong_storage_data_41 ^ i_input_data[850 % IN_WIDTH];
                918 / IN_WIDTH: pong_storage_data_41 <= (fillup_transition == 1'b1) ? i_input_data[918 % IN_WIDTH] : pong_storage_data_41 ^ i_input_data[918 % IN_WIDTH];
                default: pong_storage_data_41 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_41;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_41 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_41;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_41 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_41;
            end
        end
    end
end

logic ping_storage_data_42;
logic pong_storage_data_42;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_42 <= 1'b0;
        pong_storage_data_42 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                140 / IN_WIDTH: ping_storage_data_42 <= (fillup_transition == 1'b1) ? i_input_data[140 % IN_WIDTH] : ping_storage_data_42 ^ i_input_data[140 % IN_WIDTH];
                257 / IN_WIDTH: ping_storage_data_42 <= (fillup_transition == 1'b1) ? i_input_data[257 % IN_WIDTH] : ping_storage_data_42 ^ i_input_data[257 % IN_WIDTH];
                851 / IN_WIDTH: ping_storage_data_42 <= (fillup_transition == 1'b1) ? i_input_data[851 % IN_WIDTH] : ping_storage_data_42 ^ i_input_data[851 % IN_WIDTH];
                919 / IN_WIDTH: ping_storage_data_42 <= (fillup_transition == 1'b1) ? i_input_data[919 % IN_WIDTH] : ping_storage_data_42 ^ i_input_data[919 % IN_WIDTH];
                default: ping_storage_data_42 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_42;
                endcase
            end else begin
                case (input_count)
                140 / IN_WIDTH: pong_storage_data_42 <= (fillup_transition == 1'b1) ? i_input_data[140 % IN_WIDTH] : pong_storage_data_42 ^ i_input_data[140 % IN_WIDTH];
                257 / IN_WIDTH: pong_storage_data_42 <= (fillup_transition == 1'b1) ? i_input_data[257 % IN_WIDTH] : pong_storage_data_42 ^ i_input_data[257 % IN_WIDTH];
                851 / IN_WIDTH: pong_storage_data_42 <= (fillup_transition == 1'b1) ? i_input_data[851 % IN_WIDTH] : pong_storage_data_42 ^ i_input_data[851 % IN_WIDTH];
                919 / IN_WIDTH: pong_storage_data_42 <= (fillup_transition == 1'b1) ? i_input_data[919 % IN_WIDTH] : pong_storage_data_42 ^ i_input_data[919 % IN_WIDTH];
                default: pong_storage_data_42 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_42;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_42 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_42;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_42 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_42;
            end
        end
    end
end

logic ping_storage_data_43;
logic pong_storage_data_43;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_43 <= 1'b0;
        pong_storage_data_43 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                141 / IN_WIDTH: ping_storage_data_43 <= (fillup_transition == 1'b1) ? i_input_data[141 % IN_WIDTH] : ping_storage_data_43 ^ i_input_data[141 % IN_WIDTH];
                258 / IN_WIDTH: ping_storage_data_43 <= (fillup_transition == 1'b1) ? i_input_data[258 % IN_WIDTH] : ping_storage_data_43 ^ i_input_data[258 % IN_WIDTH];
                852 / IN_WIDTH: ping_storage_data_43 <= (fillup_transition == 1'b1) ? i_input_data[852 % IN_WIDTH] : ping_storage_data_43 ^ i_input_data[852 % IN_WIDTH];
                920 / IN_WIDTH: ping_storage_data_43 <= (fillup_transition == 1'b1) ? i_input_data[920 % IN_WIDTH] : ping_storage_data_43 ^ i_input_data[920 % IN_WIDTH];
                default: ping_storage_data_43 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_43;
                endcase
            end else begin
                case (input_count)
                141 / IN_WIDTH: pong_storage_data_43 <= (fillup_transition == 1'b1) ? i_input_data[141 % IN_WIDTH] : pong_storage_data_43 ^ i_input_data[141 % IN_WIDTH];
                258 / IN_WIDTH: pong_storage_data_43 <= (fillup_transition == 1'b1) ? i_input_data[258 % IN_WIDTH] : pong_storage_data_43 ^ i_input_data[258 % IN_WIDTH];
                852 / IN_WIDTH: pong_storage_data_43 <= (fillup_transition == 1'b1) ? i_input_data[852 % IN_WIDTH] : pong_storage_data_43 ^ i_input_data[852 % IN_WIDTH];
                920 / IN_WIDTH: pong_storage_data_43 <= (fillup_transition == 1'b1) ? i_input_data[920 % IN_WIDTH] : pong_storage_data_43 ^ i_input_data[920 % IN_WIDTH];
                default: pong_storage_data_43 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_43;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_43 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_43;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_43 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_43;
            end
        end
    end
end

logic ping_storage_data_44;
logic pong_storage_data_44;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_44 <= 1'b0;
        pong_storage_data_44 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                142 / IN_WIDTH: ping_storage_data_44 <= (fillup_transition == 1'b1) ? i_input_data[142 % IN_WIDTH] : ping_storage_data_44 ^ i_input_data[142 % IN_WIDTH];
                259 / IN_WIDTH: ping_storage_data_44 <= (fillup_transition == 1'b1) ? i_input_data[259 % IN_WIDTH] : ping_storage_data_44 ^ i_input_data[259 % IN_WIDTH];
                853 / IN_WIDTH: ping_storage_data_44 <= (fillup_transition == 1'b1) ? i_input_data[853 % IN_WIDTH] : ping_storage_data_44 ^ i_input_data[853 % IN_WIDTH];
                921 / IN_WIDTH: ping_storage_data_44 <= (fillup_transition == 1'b1) ? i_input_data[921 % IN_WIDTH] : ping_storage_data_44 ^ i_input_data[921 % IN_WIDTH];
                default: ping_storage_data_44 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_44;
                endcase
            end else begin
                case (input_count)
                142 / IN_WIDTH: pong_storage_data_44 <= (fillup_transition == 1'b1) ? i_input_data[142 % IN_WIDTH] : pong_storage_data_44 ^ i_input_data[142 % IN_WIDTH];
                259 / IN_WIDTH: pong_storage_data_44 <= (fillup_transition == 1'b1) ? i_input_data[259 % IN_WIDTH] : pong_storage_data_44 ^ i_input_data[259 % IN_WIDTH];
                853 / IN_WIDTH: pong_storage_data_44 <= (fillup_transition == 1'b1) ? i_input_data[853 % IN_WIDTH] : pong_storage_data_44 ^ i_input_data[853 % IN_WIDTH];
                921 / IN_WIDTH: pong_storage_data_44 <= (fillup_transition == 1'b1) ? i_input_data[921 % IN_WIDTH] : pong_storage_data_44 ^ i_input_data[921 % IN_WIDTH];
                default: pong_storage_data_44 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_44;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_44 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_44;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_44 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_44;
            end
        end
    end
end

logic ping_storage_data_45;
logic pong_storage_data_45;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_45 <= 1'b0;
        pong_storage_data_45 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                143 / IN_WIDTH: ping_storage_data_45 <= (fillup_transition == 1'b1) ? i_input_data[143 % IN_WIDTH] : ping_storage_data_45 ^ i_input_data[143 % IN_WIDTH];
                260 / IN_WIDTH: ping_storage_data_45 <= (fillup_transition == 1'b1) ? i_input_data[260 % IN_WIDTH] : ping_storage_data_45 ^ i_input_data[260 % IN_WIDTH];
                854 / IN_WIDTH: ping_storage_data_45 <= (fillup_transition == 1'b1) ? i_input_data[854 % IN_WIDTH] : ping_storage_data_45 ^ i_input_data[854 % IN_WIDTH];
                922 / IN_WIDTH: ping_storage_data_45 <= (fillup_transition == 1'b1) ? i_input_data[922 % IN_WIDTH] : ping_storage_data_45 ^ i_input_data[922 % IN_WIDTH];
                default: ping_storage_data_45 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_45;
                endcase
            end else begin
                case (input_count)
                143 / IN_WIDTH: pong_storage_data_45 <= (fillup_transition == 1'b1) ? i_input_data[143 % IN_WIDTH] : pong_storage_data_45 ^ i_input_data[143 % IN_WIDTH];
                260 / IN_WIDTH: pong_storage_data_45 <= (fillup_transition == 1'b1) ? i_input_data[260 % IN_WIDTH] : pong_storage_data_45 ^ i_input_data[260 % IN_WIDTH];
                854 / IN_WIDTH: pong_storage_data_45 <= (fillup_transition == 1'b1) ? i_input_data[854 % IN_WIDTH] : pong_storage_data_45 ^ i_input_data[854 % IN_WIDTH];
                922 / IN_WIDTH: pong_storage_data_45 <= (fillup_transition == 1'b1) ? i_input_data[922 % IN_WIDTH] : pong_storage_data_45 ^ i_input_data[922 % IN_WIDTH];
                default: pong_storage_data_45 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_45;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_45 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_45;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_45 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_45;
            end
        end
    end
end

logic ping_storage_data_46;
logic pong_storage_data_46;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_46 <= 1'b0;
        pong_storage_data_46 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                144 / IN_WIDTH: ping_storage_data_46 <= (fillup_transition == 1'b1) ? i_input_data[144 % IN_WIDTH] : ping_storage_data_46 ^ i_input_data[144 % IN_WIDTH];
                261 / IN_WIDTH: ping_storage_data_46 <= (fillup_transition == 1'b1) ? i_input_data[261 % IN_WIDTH] : ping_storage_data_46 ^ i_input_data[261 % IN_WIDTH];
                855 / IN_WIDTH: ping_storage_data_46 <= (fillup_transition == 1'b1) ? i_input_data[855 % IN_WIDTH] : ping_storage_data_46 ^ i_input_data[855 % IN_WIDTH];
                923 / IN_WIDTH: ping_storage_data_46 <= (fillup_transition == 1'b1) ? i_input_data[923 % IN_WIDTH] : ping_storage_data_46 ^ i_input_data[923 % IN_WIDTH];
                default: ping_storage_data_46 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_46;
                endcase
            end else begin
                case (input_count)
                144 / IN_WIDTH: pong_storage_data_46 <= (fillup_transition == 1'b1) ? i_input_data[144 % IN_WIDTH] : pong_storage_data_46 ^ i_input_data[144 % IN_WIDTH];
                261 / IN_WIDTH: pong_storage_data_46 <= (fillup_transition == 1'b1) ? i_input_data[261 % IN_WIDTH] : pong_storage_data_46 ^ i_input_data[261 % IN_WIDTH];
                855 / IN_WIDTH: pong_storage_data_46 <= (fillup_transition == 1'b1) ? i_input_data[855 % IN_WIDTH] : pong_storage_data_46 ^ i_input_data[855 % IN_WIDTH];
                923 / IN_WIDTH: pong_storage_data_46 <= (fillup_transition == 1'b1) ? i_input_data[923 % IN_WIDTH] : pong_storage_data_46 ^ i_input_data[923 % IN_WIDTH];
                default: pong_storage_data_46 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_46;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_46 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_46;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_46 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_46;
            end
        end
    end
end

logic ping_storage_data_47;
logic pong_storage_data_47;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_47 <= 1'b0;
        pong_storage_data_47 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                145 / IN_WIDTH: ping_storage_data_47 <= (fillup_transition == 1'b1) ? i_input_data[145 % IN_WIDTH] : ping_storage_data_47 ^ i_input_data[145 % IN_WIDTH];
                262 / IN_WIDTH: ping_storage_data_47 <= (fillup_transition == 1'b1) ? i_input_data[262 % IN_WIDTH] : ping_storage_data_47 ^ i_input_data[262 % IN_WIDTH];
                856 / IN_WIDTH: ping_storage_data_47 <= (fillup_transition == 1'b1) ? i_input_data[856 % IN_WIDTH] : ping_storage_data_47 ^ i_input_data[856 % IN_WIDTH];
                924 / IN_WIDTH: ping_storage_data_47 <= (fillup_transition == 1'b1) ? i_input_data[924 % IN_WIDTH] : ping_storage_data_47 ^ i_input_data[924 % IN_WIDTH];
                default: ping_storage_data_47 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_47;
                endcase
            end else begin
                case (input_count)
                145 / IN_WIDTH: pong_storage_data_47 <= (fillup_transition == 1'b1) ? i_input_data[145 % IN_WIDTH] : pong_storage_data_47 ^ i_input_data[145 % IN_WIDTH];
                262 / IN_WIDTH: pong_storage_data_47 <= (fillup_transition == 1'b1) ? i_input_data[262 % IN_WIDTH] : pong_storage_data_47 ^ i_input_data[262 % IN_WIDTH];
                856 / IN_WIDTH: pong_storage_data_47 <= (fillup_transition == 1'b1) ? i_input_data[856 % IN_WIDTH] : pong_storage_data_47 ^ i_input_data[856 % IN_WIDTH];
                924 / IN_WIDTH: pong_storage_data_47 <= (fillup_transition == 1'b1) ? i_input_data[924 % IN_WIDTH] : pong_storage_data_47 ^ i_input_data[924 % IN_WIDTH];
                default: pong_storage_data_47 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_47;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_47 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_47;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_47 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_47;
            end
        end
    end
end

logic ping_storage_data_48;
logic pong_storage_data_48;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_48 <= 1'b0;
        pong_storage_data_48 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                146 / IN_WIDTH: ping_storage_data_48 <= (fillup_transition == 1'b1) ? i_input_data[146 % IN_WIDTH] : ping_storage_data_48 ^ i_input_data[146 % IN_WIDTH];
                263 / IN_WIDTH: ping_storage_data_48 <= (fillup_transition == 1'b1) ? i_input_data[263 % IN_WIDTH] : ping_storage_data_48 ^ i_input_data[263 % IN_WIDTH];
                857 / IN_WIDTH: ping_storage_data_48 <= (fillup_transition == 1'b1) ? i_input_data[857 % IN_WIDTH] : ping_storage_data_48 ^ i_input_data[857 % IN_WIDTH];
                925 / IN_WIDTH: ping_storage_data_48 <= (fillup_transition == 1'b1) ? i_input_data[925 % IN_WIDTH] : ping_storage_data_48 ^ i_input_data[925 % IN_WIDTH];
                default: ping_storage_data_48 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_48;
                endcase
            end else begin
                case (input_count)
                146 / IN_WIDTH: pong_storage_data_48 <= (fillup_transition == 1'b1) ? i_input_data[146 % IN_WIDTH] : pong_storage_data_48 ^ i_input_data[146 % IN_WIDTH];
                263 / IN_WIDTH: pong_storage_data_48 <= (fillup_transition == 1'b1) ? i_input_data[263 % IN_WIDTH] : pong_storage_data_48 ^ i_input_data[263 % IN_WIDTH];
                857 / IN_WIDTH: pong_storage_data_48 <= (fillup_transition == 1'b1) ? i_input_data[857 % IN_WIDTH] : pong_storage_data_48 ^ i_input_data[857 % IN_WIDTH];
                925 / IN_WIDTH: pong_storage_data_48 <= (fillup_transition == 1'b1) ? i_input_data[925 % IN_WIDTH] : pong_storage_data_48 ^ i_input_data[925 % IN_WIDTH];
                default: pong_storage_data_48 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_48;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_48 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_48;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_48 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_48;
            end
        end
    end
end

logic ping_storage_data_49;
logic pong_storage_data_49;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_49 <= 1'b0;
        pong_storage_data_49 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                147 / IN_WIDTH: ping_storage_data_49 <= (fillup_transition == 1'b1) ? i_input_data[147 % IN_WIDTH] : ping_storage_data_49 ^ i_input_data[147 % IN_WIDTH];
                264 / IN_WIDTH: ping_storage_data_49 <= (fillup_transition == 1'b1) ? i_input_data[264 % IN_WIDTH] : ping_storage_data_49 ^ i_input_data[264 % IN_WIDTH];
                858 / IN_WIDTH: ping_storage_data_49 <= (fillup_transition == 1'b1) ? i_input_data[858 % IN_WIDTH] : ping_storage_data_49 ^ i_input_data[858 % IN_WIDTH];
                926 / IN_WIDTH: ping_storage_data_49 <= (fillup_transition == 1'b1) ? i_input_data[926 % IN_WIDTH] : ping_storage_data_49 ^ i_input_data[926 % IN_WIDTH];
                default: ping_storage_data_49 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_49;
                endcase
            end else begin
                case (input_count)
                147 / IN_WIDTH: pong_storage_data_49 <= (fillup_transition == 1'b1) ? i_input_data[147 % IN_WIDTH] : pong_storage_data_49 ^ i_input_data[147 % IN_WIDTH];
                264 / IN_WIDTH: pong_storage_data_49 <= (fillup_transition == 1'b1) ? i_input_data[264 % IN_WIDTH] : pong_storage_data_49 ^ i_input_data[264 % IN_WIDTH];
                858 / IN_WIDTH: pong_storage_data_49 <= (fillup_transition == 1'b1) ? i_input_data[858 % IN_WIDTH] : pong_storage_data_49 ^ i_input_data[858 % IN_WIDTH];
                926 / IN_WIDTH: pong_storage_data_49 <= (fillup_transition == 1'b1) ? i_input_data[926 % IN_WIDTH] : pong_storage_data_49 ^ i_input_data[926 % IN_WIDTH];
                default: pong_storage_data_49 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_49;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_49 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_49;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_49 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_49;
            end
        end
    end
end

logic ping_storage_data_50;
logic pong_storage_data_50;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_50 <= 1'b0;
        pong_storage_data_50 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                148 / IN_WIDTH: ping_storage_data_50 <= (fillup_transition == 1'b1) ? i_input_data[148 % IN_WIDTH] : ping_storage_data_50 ^ i_input_data[148 % IN_WIDTH];
                265 / IN_WIDTH: ping_storage_data_50 <= (fillup_transition == 1'b1) ? i_input_data[265 % IN_WIDTH] : ping_storage_data_50 ^ i_input_data[265 % IN_WIDTH];
                859 / IN_WIDTH: ping_storage_data_50 <= (fillup_transition == 1'b1) ? i_input_data[859 % IN_WIDTH] : ping_storage_data_50 ^ i_input_data[859 % IN_WIDTH];
                927 / IN_WIDTH: ping_storage_data_50 <= (fillup_transition == 1'b1) ? i_input_data[927 % IN_WIDTH] : ping_storage_data_50 ^ i_input_data[927 % IN_WIDTH];
                default: ping_storage_data_50 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_50;
                endcase
            end else begin
                case (input_count)
                148 / IN_WIDTH: pong_storage_data_50 <= (fillup_transition == 1'b1) ? i_input_data[148 % IN_WIDTH] : pong_storage_data_50 ^ i_input_data[148 % IN_WIDTH];
                265 / IN_WIDTH: pong_storage_data_50 <= (fillup_transition == 1'b1) ? i_input_data[265 % IN_WIDTH] : pong_storage_data_50 ^ i_input_data[265 % IN_WIDTH];
                859 / IN_WIDTH: pong_storage_data_50 <= (fillup_transition == 1'b1) ? i_input_data[859 % IN_WIDTH] : pong_storage_data_50 ^ i_input_data[859 % IN_WIDTH];
                927 / IN_WIDTH: pong_storage_data_50 <= (fillup_transition == 1'b1) ? i_input_data[927 % IN_WIDTH] : pong_storage_data_50 ^ i_input_data[927 % IN_WIDTH];
                default: pong_storage_data_50 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_50;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_50 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_50;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_50 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_50;
            end
        end
    end
end

logic ping_storage_data_51;
logic pong_storage_data_51;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_51 <= 1'b0;
        pong_storage_data_51 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                149 / IN_WIDTH: ping_storage_data_51 <= (fillup_transition == 1'b1) ? i_input_data[149 % IN_WIDTH] : ping_storage_data_51 ^ i_input_data[149 % IN_WIDTH];
                266 / IN_WIDTH: ping_storage_data_51 <= (fillup_transition == 1'b1) ? i_input_data[266 % IN_WIDTH] : ping_storage_data_51 ^ i_input_data[266 % IN_WIDTH];
                860 / IN_WIDTH: ping_storage_data_51 <= (fillup_transition == 1'b1) ? i_input_data[860 % IN_WIDTH] : ping_storage_data_51 ^ i_input_data[860 % IN_WIDTH];
                928 / IN_WIDTH: ping_storage_data_51 <= (fillup_transition == 1'b1) ? i_input_data[928 % IN_WIDTH] : ping_storage_data_51 ^ i_input_data[928 % IN_WIDTH];
                default: ping_storage_data_51 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_51;
                endcase
            end else begin
                case (input_count)
                149 / IN_WIDTH: pong_storage_data_51 <= (fillup_transition == 1'b1) ? i_input_data[149 % IN_WIDTH] : pong_storage_data_51 ^ i_input_data[149 % IN_WIDTH];
                266 / IN_WIDTH: pong_storage_data_51 <= (fillup_transition == 1'b1) ? i_input_data[266 % IN_WIDTH] : pong_storage_data_51 ^ i_input_data[266 % IN_WIDTH];
                860 / IN_WIDTH: pong_storage_data_51 <= (fillup_transition == 1'b1) ? i_input_data[860 % IN_WIDTH] : pong_storage_data_51 ^ i_input_data[860 % IN_WIDTH];
                928 / IN_WIDTH: pong_storage_data_51 <= (fillup_transition == 1'b1) ? i_input_data[928 % IN_WIDTH] : pong_storage_data_51 ^ i_input_data[928 % IN_WIDTH];
                default: pong_storage_data_51 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_51;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_51 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_51;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_51 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_51;
            end
        end
    end
end

logic ping_storage_data_52;
logic pong_storage_data_52;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_52 <= 1'b0;
        pong_storage_data_52 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                150 / IN_WIDTH: ping_storage_data_52 <= (fillup_transition == 1'b1) ? i_input_data[150 % IN_WIDTH] : ping_storage_data_52 ^ i_input_data[150 % IN_WIDTH];
                267 / IN_WIDTH: ping_storage_data_52 <= (fillup_transition == 1'b1) ? i_input_data[267 % IN_WIDTH] : ping_storage_data_52 ^ i_input_data[267 % IN_WIDTH];
                861 / IN_WIDTH: ping_storage_data_52 <= (fillup_transition == 1'b1) ? i_input_data[861 % IN_WIDTH] : ping_storage_data_52 ^ i_input_data[861 % IN_WIDTH];
                929 / IN_WIDTH: ping_storage_data_52 <= (fillup_transition == 1'b1) ? i_input_data[929 % IN_WIDTH] : ping_storage_data_52 ^ i_input_data[929 % IN_WIDTH];
                default: ping_storage_data_52 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_52;
                endcase
            end else begin
                case (input_count)
                150 / IN_WIDTH: pong_storage_data_52 <= (fillup_transition == 1'b1) ? i_input_data[150 % IN_WIDTH] : pong_storage_data_52 ^ i_input_data[150 % IN_WIDTH];
                267 / IN_WIDTH: pong_storage_data_52 <= (fillup_transition == 1'b1) ? i_input_data[267 % IN_WIDTH] : pong_storage_data_52 ^ i_input_data[267 % IN_WIDTH];
                861 / IN_WIDTH: pong_storage_data_52 <= (fillup_transition == 1'b1) ? i_input_data[861 % IN_WIDTH] : pong_storage_data_52 ^ i_input_data[861 % IN_WIDTH];
                929 / IN_WIDTH: pong_storage_data_52 <= (fillup_transition == 1'b1) ? i_input_data[929 % IN_WIDTH] : pong_storage_data_52 ^ i_input_data[929 % IN_WIDTH];
                default: pong_storage_data_52 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_52;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_52 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_52;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_52 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_52;
            end
        end
    end
end

logic ping_storage_data_53;
logic pong_storage_data_53;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_53 <= 1'b0;
        pong_storage_data_53 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                151 / IN_WIDTH: ping_storage_data_53 <= (fillup_transition == 1'b1) ? i_input_data[151 % IN_WIDTH] : ping_storage_data_53 ^ i_input_data[151 % IN_WIDTH];
                268 / IN_WIDTH: ping_storage_data_53 <= (fillup_transition == 1'b1) ? i_input_data[268 % IN_WIDTH] : ping_storage_data_53 ^ i_input_data[268 % IN_WIDTH];
                862 / IN_WIDTH: ping_storage_data_53 <= (fillup_transition == 1'b1) ? i_input_data[862 % IN_WIDTH] : ping_storage_data_53 ^ i_input_data[862 % IN_WIDTH];
                930 / IN_WIDTH: ping_storage_data_53 <= (fillup_transition == 1'b1) ? i_input_data[930 % IN_WIDTH] : ping_storage_data_53 ^ i_input_data[930 % IN_WIDTH];
                default: ping_storage_data_53 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_53;
                endcase
            end else begin
                case (input_count)
                151 / IN_WIDTH: pong_storage_data_53 <= (fillup_transition == 1'b1) ? i_input_data[151 % IN_WIDTH] : pong_storage_data_53 ^ i_input_data[151 % IN_WIDTH];
                268 / IN_WIDTH: pong_storage_data_53 <= (fillup_transition == 1'b1) ? i_input_data[268 % IN_WIDTH] : pong_storage_data_53 ^ i_input_data[268 % IN_WIDTH];
                862 / IN_WIDTH: pong_storage_data_53 <= (fillup_transition == 1'b1) ? i_input_data[862 % IN_WIDTH] : pong_storage_data_53 ^ i_input_data[862 % IN_WIDTH];
                930 / IN_WIDTH: pong_storage_data_53 <= (fillup_transition == 1'b1) ? i_input_data[930 % IN_WIDTH] : pong_storage_data_53 ^ i_input_data[930 % IN_WIDTH];
                default: pong_storage_data_53 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_53;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_53 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_53;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_53 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_53;
            end
        end
    end
end

logic ping_storage_data_54;
logic pong_storage_data_54;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_54 <= 1'b0;
        pong_storage_data_54 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                152 / IN_WIDTH: ping_storage_data_54 <= (fillup_transition == 1'b1) ? i_input_data[152 % IN_WIDTH] : ping_storage_data_54 ^ i_input_data[152 % IN_WIDTH];
                269 / IN_WIDTH: ping_storage_data_54 <= (fillup_transition == 1'b1) ? i_input_data[269 % IN_WIDTH] : ping_storage_data_54 ^ i_input_data[269 % IN_WIDTH];
                863 / IN_WIDTH: ping_storage_data_54 <= (fillup_transition == 1'b1) ? i_input_data[863 % IN_WIDTH] : ping_storage_data_54 ^ i_input_data[863 % IN_WIDTH];
                931 / IN_WIDTH: ping_storage_data_54 <= (fillup_transition == 1'b1) ? i_input_data[931 % IN_WIDTH] : ping_storage_data_54 ^ i_input_data[931 % IN_WIDTH];
                default: ping_storage_data_54 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_54;
                endcase
            end else begin
                case (input_count)
                152 / IN_WIDTH: pong_storage_data_54 <= (fillup_transition == 1'b1) ? i_input_data[152 % IN_WIDTH] : pong_storage_data_54 ^ i_input_data[152 % IN_WIDTH];
                269 / IN_WIDTH: pong_storage_data_54 <= (fillup_transition == 1'b1) ? i_input_data[269 % IN_WIDTH] : pong_storage_data_54 ^ i_input_data[269 % IN_WIDTH];
                863 / IN_WIDTH: pong_storage_data_54 <= (fillup_transition == 1'b1) ? i_input_data[863 % IN_WIDTH] : pong_storage_data_54 ^ i_input_data[863 % IN_WIDTH];
                931 / IN_WIDTH: pong_storage_data_54 <= (fillup_transition == 1'b1) ? i_input_data[931 % IN_WIDTH] : pong_storage_data_54 ^ i_input_data[931 % IN_WIDTH];
                default: pong_storage_data_54 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_54;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_54 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_54;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_54 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_54;
            end
        end
    end
end

logic ping_storage_data_55;
logic pong_storage_data_55;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_55 <= 1'b0;
        pong_storage_data_55 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                153 / IN_WIDTH: ping_storage_data_55 <= (fillup_transition == 1'b1) ? i_input_data[153 % IN_WIDTH] : ping_storage_data_55 ^ i_input_data[153 % IN_WIDTH];
                270 / IN_WIDTH: ping_storage_data_55 <= (fillup_transition == 1'b1) ? i_input_data[270 % IN_WIDTH] : ping_storage_data_55 ^ i_input_data[270 % IN_WIDTH];
                768 / IN_WIDTH: ping_storage_data_55 <= (fillup_transition == 1'b1) ? i_input_data[768 % IN_WIDTH] : ping_storage_data_55 ^ i_input_data[768 % IN_WIDTH];
                932 / IN_WIDTH: ping_storage_data_55 <= (fillup_transition == 1'b1) ? i_input_data[932 % IN_WIDTH] : ping_storage_data_55 ^ i_input_data[932 % IN_WIDTH];
                default: ping_storage_data_55 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_55;
                endcase
            end else begin
                case (input_count)
                153 / IN_WIDTH: pong_storage_data_55 <= (fillup_transition == 1'b1) ? i_input_data[153 % IN_WIDTH] : pong_storage_data_55 ^ i_input_data[153 % IN_WIDTH];
                270 / IN_WIDTH: pong_storage_data_55 <= (fillup_transition == 1'b1) ? i_input_data[270 % IN_WIDTH] : pong_storage_data_55 ^ i_input_data[270 % IN_WIDTH];
                768 / IN_WIDTH: pong_storage_data_55 <= (fillup_transition == 1'b1) ? i_input_data[768 % IN_WIDTH] : pong_storage_data_55 ^ i_input_data[768 % IN_WIDTH];
                932 / IN_WIDTH: pong_storage_data_55 <= (fillup_transition == 1'b1) ? i_input_data[932 % IN_WIDTH] : pong_storage_data_55 ^ i_input_data[932 % IN_WIDTH];
                default: pong_storage_data_55 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_55;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_55 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_55;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_55 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_55;
            end
        end
    end
end

logic ping_storage_data_56;
logic pong_storage_data_56;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_56 <= 1'b0;
        pong_storage_data_56 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                154 / IN_WIDTH: ping_storage_data_56 <= (fillup_transition == 1'b1) ? i_input_data[154 % IN_WIDTH] : ping_storage_data_56 ^ i_input_data[154 % IN_WIDTH];
                271 / IN_WIDTH: ping_storage_data_56 <= (fillup_transition == 1'b1) ? i_input_data[271 % IN_WIDTH] : ping_storage_data_56 ^ i_input_data[271 % IN_WIDTH];
                769 / IN_WIDTH: ping_storage_data_56 <= (fillup_transition == 1'b1) ? i_input_data[769 % IN_WIDTH] : ping_storage_data_56 ^ i_input_data[769 % IN_WIDTH];
                933 / IN_WIDTH: ping_storage_data_56 <= (fillup_transition == 1'b1) ? i_input_data[933 % IN_WIDTH] : ping_storage_data_56 ^ i_input_data[933 % IN_WIDTH];
                default: ping_storage_data_56 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_56;
                endcase
            end else begin
                case (input_count)
                154 / IN_WIDTH: pong_storage_data_56 <= (fillup_transition == 1'b1) ? i_input_data[154 % IN_WIDTH] : pong_storage_data_56 ^ i_input_data[154 % IN_WIDTH];
                271 / IN_WIDTH: pong_storage_data_56 <= (fillup_transition == 1'b1) ? i_input_data[271 % IN_WIDTH] : pong_storage_data_56 ^ i_input_data[271 % IN_WIDTH];
                769 / IN_WIDTH: pong_storage_data_56 <= (fillup_transition == 1'b1) ? i_input_data[769 % IN_WIDTH] : pong_storage_data_56 ^ i_input_data[769 % IN_WIDTH];
                933 / IN_WIDTH: pong_storage_data_56 <= (fillup_transition == 1'b1) ? i_input_data[933 % IN_WIDTH] : pong_storage_data_56 ^ i_input_data[933 % IN_WIDTH];
                default: pong_storage_data_56 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_56;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_56 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_56;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_56 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_56;
            end
        end
    end
end

logic ping_storage_data_57;
logic pong_storage_data_57;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_57 <= 1'b0;
        pong_storage_data_57 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                155 / IN_WIDTH: ping_storage_data_57 <= (fillup_transition == 1'b1) ? i_input_data[155 % IN_WIDTH] : ping_storage_data_57 ^ i_input_data[155 % IN_WIDTH];
                272 / IN_WIDTH: ping_storage_data_57 <= (fillup_transition == 1'b1) ? i_input_data[272 % IN_WIDTH] : ping_storage_data_57 ^ i_input_data[272 % IN_WIDTH];
                770 / IN_WIDTH: ping_storage_data_57 <= (fillup_transition == 1'b1) ? i_input_data[770 % IN_WIDTH] : ping_storage_data_57 ^ i_input_data[770 % IN_WIDTH];
                934 / IN_WIDTH: ping_storage_data_57 <= (fillup_transition == 1'b1) ? i_input_data[934 % IN_WIDTH] : ping_storage_data_57 ^ i_input_data[934 % IN_WIDTH];
                default: ping_storage_data_57 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_57;
                endcase
            end else begin
                case (input_count)
                155 / IN_WIDTH: pong_storage_data_57 <= (fillup_transition == 1'b1) ? i_input_data[155 % IN_WIDTH] : pong_storage_data_57 ^ i_input_data[155 % IN_WIDTH];
                272 / IN_WIDTH: pong_storage_data_57 <= (fillup_transition == 1'b1) ? i_input_data[272 % IN_WIDTH] : pong_storage_data_57 ^ i_input_data[272 % IN_WIDTH];
                770 / IN_WIDTH: pong_storage_data_57 <= (fillup_transition == 1'b1) ? i_input_data[770 % IN_WIDTH] : pong_storage_data_57 ^ i_input_data[770 % IN_WIDTH];
                934 / IN_WIDTH: pong_storage_data_57 <= (fillup_transition == 1'b1) ? i_input_data[934 % IN_WIDTH] : pong_storage_data_57 ^ i_input_data[934 % IN_WIDTH];
                default: pong_storage_data_57 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_57;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_57 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_57;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_57 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_57;
            end
        end
    end
end

logic ping_storage_data_58;
logic pong_storage_data_58;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_58 <= 1'b0;
        pong_storage_data_58 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                156 / IN_WIDTH: ping_storage_data_58 <= (fillup_transition == 1'b1) ? i_input_data[156 % IN_WIDTH] : ping_storage_data_58 ^ i_input_data[156 % IN_WIDTH];
                273 / IN_WIDTH: ping_storage_data_58 <= (fillup_transition == 1'b1) ? i_input_data[273 % IN_WIDTH] : ping_storage_data_58 ^ i_input_data[273 % IN_WIDTH];
                771 / IN_WIDTH: ping_storage_data_58 <= (fillup_transition == 1'b1) ? i_input_data[771 % IN_WIDTH] : ping_storage_data_58 ^ i_input_data[771 % IN_WIDTH];
                935 / IN_WIDTH: ping_storage_data_58 <= (fillup_transition == 1'b1) ? i_input_data[935 % IN_WIDTH] : ping_storage_data_58 ^ i_input_data[935 % IN_WIDTH];
                default: ping_storage_data_58 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_58;
                endcase
            end else begin
                case (input_count)
                156 / IN_WIDTH: pong_storage_data_58 <= (fillup_transition == 1'b1) ? i_input_data[156 % IN_WIDTH] : pong_storage_data_58 ^ i_input_data[156 % IN_WIDTH];
                273 / IN_WIDTH: pong_storage_data_58 <= (fillup_transition == 1'b1) ? i_input_data[273 % IN_WIDTH] : pong_storage_data_58 ^ i_input_data[273 % IN_WIDTH];
                771 / IN_WIDTH: pong_storage_data_58 <= (fillup_transition == 1'b1) ? i_input_data[771 % IN_WIDTH] : pong_storage_data_58 ^ i_input_data[771 % IN_WIDTH];
                935 / IN_WIDTH: pong_storage_data_58 <= (fillup_transition == 1'b1) ? i_input_data[935 % IN_WIDTH] : pong_storage_data_58 ^ i_input_data[935 % IN_WIDTH];
                default: pong_storage_data_58 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_58;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_58 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_58;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_58 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_58;
            end
        end
    end
end

logic ping_storage_data_59;
logic pong_storage_data_59;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_59 <= 1'b0;
        pong_storage_data_59 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                157 / IN_WIDTH: ping_storage_data_59 <= (fillup_transition == 1'b1) ? i_input_data[157 % IN_WIDTH] : ping_storage_data_59 ^ i_input_data[157 % IN_WIDTH];
                274 / IN_WIDTH: ping_storage_data_59 <= (fillup_transition == 1'b1) ? i_input_data[274 % IN_WIDTH] : ping_storage_data_59 ^ i_input_data[274 % IN_WIDTH];
                772 / IN_WIDTH: ping_storage_data_59 <= (fillup_transition == 1'b1) ? i_input_data[772 % IN_WIDTH] : ping_storage_data_59 ^ i_input_data[772 % IN_WIDTH];
                936 / IN_WIDTH: ping_storage_data_59 <= (fillup_transition == 1'b1) ? i_input_data[936 % IN_WIDTH] : ping_storage_data_59 ^ i_input_data[936 % IN_WIDTH];
                default: ping_storage_data_59 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_59;
                endcase
            end else begin
                case (input_count)
                157 / IN_WIDTH: pong_storage_data_59 <= (fillup_transition == 1'b1) ? i_input_data[157 % IN_WIDTH] : pong_storage_data_59 ^ i_input_data[157 % IN_WIDTH];
                274 / IN_WIDTH: pong_storage_data_59 <= (fillup_transition == 1'b1) ? i_input_data[274 % IN_WIDTH] : pong_storage_data_59 ^ i_input_data[274 % IN_WIDTH];
                772 / IN_WIDTH: pong_storage_data_59 <= (fillup_transition == 1'b1) ? i_input_data[772 % IN_WIDTH] : pong_storage_data_59 ^ i_input_data[772 % IN_WIDTH];
                936 / IN_WIDTH: pong_storage_data_59 <= (fillup_transition == 1'b1) ? i_input_data[936 % IN_WIDTH] : pong_storage_data_59 ^ i_input_data[936 % IN_WIDTH];
                default: pong_storage_data_59 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_59;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_59 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_59;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_59 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_59;
            end
        end
    end
end

logic ping_storage_data_60;
logic pong_storage_data_60;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_60 <= 1'b0;
        pong_storage_data_60 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                158 / IN_WIDTH: ping_storage_data_60 <= (fillup_transition == 1'b1) ? i_input_data[158 % IN_WIDTH] : ping_storage_data_60 ^ i_input_data[158 % IN_WIDTH];
                275 / IN_WIDTH: ping_storage_data_60 <= (fillup_transition == 1'b1) ? i_input_data[275 % IN_WIDTH] : ping_storage_data_60 ^ i_input_data[275 % IN_WIDTH];
                773 / IN_WIDTH: ping_storage_data_60 <= (fillup_transition == 1'b1) ? i_input_data[773 % IN_WIDTH] : ping_storage_data_60 ^ i_input_data[773 % IN_WIDTH];
                937 / IN_WIDTH: ping_storage_data_60 <= (fillup_transition == 1'b1) ? i_input_data[937 % IN_WIDTH] : ping_storage_data_60 ^ i_input_data[937 % IN_WIDTH];
                default: ping_storage_data_60 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_60;
                endcase
            end else begin
                case (input_count)
                158 / IN_WIDTH: pong_storage_data_60 <= (fillup_transition == 1'b1) ? i_input_data[158 % IN_WIDTH] : pong_storage_data_60 ^ i_input_data[158 % IN_WIDTH];
                275 / IN_WIDTH: pong_storage_data_60 <= (fillup_transition == 1'b1) ? i_input_data[275 % IN_WIDTH] : pong_storage_data_60 ^ i_input_data[275 % IN_WIDTH];
                773 / IN_WIDTH: pong_storage_data_60 <= (fillup_transition == 1'b1) ? i_input_data[773 % IN_WIDTH] : pong_storage_data_60 ^ i_input_data[773 % IN_WIDTH];
                937 / IN_WIDTH: pong_storage_data_60 <= (fillup_transition == 1'b1) ? i_input_data[937 % IN_WIDTH] : pong_storage_data_60 ^ i_input_data[937 % IN_WIDTH];
                default: pong_storage_data_60 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_60;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_60 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_60;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_60 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_60;
            end
        end
    end
end

logic ping_storage_data_61;
logic pong_storage_data_61;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_61 <= 1'b0;
        pong_storage_data_61 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                159 / IN_WIDTH: ping_storage_data_61 <= (fillup_transition == 1'b1) ? i_input_data[159 % IN_WIDTH] : ping_storage_data_61 ^ i_input_data[159 % IN_WIDTH];
                276 / IN_WIDTH: ping_storage_data_61 <= (fillup_transition == 1'b1) ? i_input_data[276 % IN_WIDTH] : ping_storage_data_61 ^ i_input_data[276 % IN_WIDTH];
                774 / IN_WIDTH: ping_storage_data_61 <= (fillup_transition == 1'b1) ? i_input_data[774 % IN_WIDTH] : ping_storage_data_61 ^ i_input_data[774 % IN_WIDTH];
                938 / IN_WIDTH: ping_storage_data_61 <= (fillup_transition == 1'b1) ? i_input_data[938 % IN_WIDTH] : ping_storage_data_61 ^ i_input_data[938 % IN_WIDTH];
                default: ping_storage_data_61 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_61;
                endcase
            end else begin
                case (input_count)
                159 / IN_WIDTH: pong_storage_data_61 <= (fillup_transition == 1'b1) ? i_input_data[159 % IN_WIDTH] : pong_storage_data_61 ^ i_input_data[159 % IN_WIDTH];
                276 / IN_WIDTH: pong_storage_data_61 <= (fillup_transition == 1'b1) ? i_input_data[276 % IN_WIDTH] : pong_storage_data_61 ^ i_input_data[276 % IN_WIDTH];
                774 / IN_WIDTH: pong_storage_data_61 <= (fillup_transition == 1'b1) ? i_input_data[774 % IN_WIDTH] : pong_storage_data_61 ^ i_input_data[774 % IN_WIDTH];
                938 / IN_WIDTH: pong_storage_data_61 <= (fillup_transition == 1'b1) ? i_input_data[938 % IN_WIDTH] : pong_storage_data_61 ^ i_input_data[938 % IN_WIDTH];
                default: pong_storage_data_61 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_61;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_61 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_61;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_61 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_61;
            end
        end
    end
end

logic ping_storage_data_62;
logic pong_storage_data_62;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_62 <= 1'b0;
        pong_storage_data_62 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                160 / IN_WIDTH: ping_storage_data_62 <= (fillup_transition == 1'b1) ? i_input_data[160 % IN_WIDTH] : ping_storage_data_62 ^ i_input_data[160 % IN_WIDTH];
                277 / IN_WIDTH: ping_storage_data_62 <= (fillup_transition == 1'b1) ? i_input_data[277 % IN_WIDTH] : ping_storage_data_62 ^ i_input_data[277 % IN_WIDTH];
                775 / IN_WIDTH: ping_storage_data_62 <= (fillup_transition == 1'b1) ? i_input_data[775 % IN_WIDTH] : ping_storage_data_62 ^ i_input_data[775 % IN_WIDTH];
                939 / IN_WIDTH: ping_storage_data_62 <= (fillup_transition == 1'b1) ? i_input_data[939 % IN_WIDTH] : ping_storage_data_62 ^ i_input_data[939 % IN_WIDTH];
                default: ping_storage_data_62 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_62;
                endcase
            end else begin
                case (input_count)
                160 / IN_WIDTH: pong_storage_data_62 <= (fillup_transition == 1'b1) ? i_input_data[160 % IN_WIDTH] : pong_storage_data_62 ^ i_input_data[160 % IN_WIDTH];
                277 / IN_WIDTH: pong_storage_data_62 <= (fillup_transition == 1'b1) ? i_input_data[277 % IN_WIDTH] : pong_storage_data_62 ^ i_input_data[277 % IN_WIDTH];
                775 / IN_WIDTH: pong_storage_data_62 <= (fillup_transition == 1'b1) ? i_input_data[775 % IN_WIDTH] : pong_storage_data_62 ^ i_input_data[775 % IN_WIDTH];
                939 / IN_WIDTH: pong_storage_data_62 <= (fillup_transition == 1'b1) ? i_input_data[939 % IN_WIDTH] : pong_storage_data_62 ^ i_input_data[939 % IN_WIDTH];
                default: pong_storage_data_62 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_62;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_62 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_62;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_62 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_62;
            end
        end
    end
end

logic ping_storage_data_63;
logic pong_storage_data_63;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_63 <= 1'b0;
        pong_storage_data_63 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                161 / IN_WIDTH: ping_storage_data_63 <= (fillup_transition == 1'b1) ? i_input_data[161 % IN_WIDTH] : ping_storage_data_63 ^ i_input_data[161 % IN_WIDTH];
                278 / IN_WIDTH: ping_storage_data_63 <= (fillup_transition == 1'b1) ? i_input_data[278 % IN_WIDTH] : ping_storage_data_63 ^ i_input_data[278 % IN_WIDTH];
                776 / IN_WIDTH: ping_storage_data_63 <= (fillup_transition == 1'b1) ? i_input_data[776 % IN_WIDTH] : ping_storage_data_63 ^ i_input_data[776 % IN_WIDTH];
                940 / IN_WIDTH: ping_storage_data_63 <= (fillup_transition == 1'b1) ? i_input_data[940 % IN_WIDTH] : ping_storage_data_63 ^ i_input_data[940 % IN_WIDTH];
                default: ping_storage_data_63 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_63;
                endcase
            end else begin
                case (input_count)
                161 / IN_WIDTH: pong_storage_data_63 <= (fillup_transition == 1'b1) ? i_input_data[161 % IN_WIDTH] : pong_storage_data_63 ^ i_input_data[161 % IN_WIDTH];
                278 / IN_WIDTH: pong_storage_data_63 <= (fillup_transition == 1'b1) ? i_input_data[278 % IN_WIDTH] : pong_storage_data_63 ^ i_input_data[278 % IN_WIDTH];
                776 / IN_WIDTH: pong_storage_data_63 <= (fillup_transition == 1'b1) ? i_input_data[776 % IN_WIDTH] : pong_storage_data_63 ^ i_input_data[776 % IN_WIDTH];
                940 / IN_WIDTH: pong_storage_data_63 <= (fillup_transition == 1'b1) ? i_input_data[940 % IN_WIDTH] : pong_storage_data_63 ^ i_input_data[940 % IN_WIDTH];
                default: pong_storage_data_63 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_63;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_63 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_63;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_63 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_63;
            end
        end
    end
end

logic ping_storage_data_64;
logic pong_storage_data_64;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_64 <= 1'b0;
        pong_storage_data_64 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                162 / IN_WIDTH: ping_storage_data_64 <= (fillup_transition == 1'b1) ? i_input_data[162 % IN_WIDTH] : ping_storage_data_64 ^ i_input_data[162 % IN_WIDTH];
                279 / IN_WIDTH: ping_storage_data_64 <= (fillup_transition == 1'b1) ? i_input_data[279 % IN_WIDTH] : ping_storage_data_64 ^ i_input_data[279 % IN_WIDTH];
                777 / IN_WIDTH: ping_storage_data_64 <= (fillup_transition == 1'b1) ? i_input_data[777 % IN_WIDTH] : ping_storage_data_64 ^ i_input_data[777 % IN_WIDTH];
                941 / IN_WIDTH: ping_storage_data_64 <= (fillup_transition == 1'b1) ? i_input_data[941 % IN_WIDTH] : ping_storage_data_64 ^ i_input_data[941 % IN_WIDTH];
                default: ping_storage_data_64 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_64;
                endcase
            end else begin
                case (input_count)
                162 / IN_WIDTH: pong_storage_data_64 <= (fillup_transition == 1'b1) ? i_input_data[162 % IN_WIDTH] : pong_storage_data_64 ^ i_input_data[162 % IN_WIDTH];
                279 / IN_WIDTH: pong_storage_data_64 <= (fillup_transition == 1'b1) ? i_input_data[279 % IN_WIDTH] : pong_storage_data_64 ^ i_input_data[279 % IN_WIDTH];
                777 / IN_WIDTH: pong_storage_data_64 <= (fillup_transition == 1'b1) ? i_input_data[777 % IN_WIDTH] : pong_storage_data_64 ^ i_input_data[777 % IN_WIDTH];
                941 / IN_WIDTH: pong_storage_data_64 <= (fillup_transition == 1'b1) ? i_input_data[941 % IN_WIDTH] : pong_storage_data_64 ^ i_input_data[941 % IN_WIDTH];
                default: pong_storage_data_64 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_64;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_64 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_64;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_64 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_64;
            end
        end
    end
end

logic ping_storage_data_65;
logic pong_storage_data_65;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_65 <= 1'b0;
        pong_storage_data_65 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                163 / IN_WIDTH: ping_storage_data_65 <= (fillup_transition == 1'b1) ? i_input_data[163 % IN_WIDTH] : ping_storage_data_65 ^ i_input_data[163 % IN_WIDTH];
                280 / IN_WIDTH: ping_storage_data_65 <= (fillup_transition == 1'b1) ? i_input_data[280 % IN_WIDTH] : ping_storage_data_65 ^ i_input_data[280 % IN_WIDTH];
                778 / IN_WIDTH: ping_storage_data_65 <= (fillup_transition == 1'b1) ? i_input_data[778 % IN_WIDTH] : ping_storage_data_65 ^ i_input_data[778 % IN_WIDTH];
                942 / IN_WIDTH: ping_storage_data_65 <= (fillup_transition == 1'b1) ? i_input_data[942 % IN_WIDTH] : ping_storage_data_65 ^ i_input_data[942 % IN_WIDTH];
                default: ping_storage_data_65 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_65;
                endcase
            end else begin
                case (input_count)
                163 / IN_WIDTH: pong_storage_data_65 <= (fillup_transition == 1'b1) ? i_input_data[163 % IN_WIDTH] : pong_storage_data_65 ^ i_input_data[163 % IN_WIDTH];
                280 / IN_WIDTH: pong_storage_data_65 <= (fillup_transition == 1'b1) ? i_input_data[280 % IN_WIDTH] : pong_storage_data_65 ^ i_input_data[280 % IN_WIDTH];
                778 / IN_WIDTH: pong_storage_data_65 <= (fillup_transition == 1'b1) ? i_input_data[778 % IN_WIDTH] : pong_storage_data_65 ^ i_input_data[778 % IN_WIDTH];
                942 / IN_WIDTH: pong_storage_data_65 <= (fillup_transition == 1'b1) ? i_input_data[942 % IN_WIDTH] : pong_storage_data_65 ^ i_input_data[942 % IN_WIDTH];
                default: pong_storage_data_65 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_65;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_65 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_65;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_65 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_65;
            end
        end
    end
end

logic ping_storage_data_66;
logic pong_storage_data_66;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_66 <= 1'b0;
        pong_storage_data_66 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                164 / IN_WIDTH: ping_storage_data_66 <= (fillup_transition == 1'b1) ? i_input_data[164 % IN_WIDTH] : ping_storage_data_66 ^ i_input_data[164 % IN_WIDTH];
                281 / IN_WIDTH: ping_storage_data_66 <= (fillup_transition == 1'b1) ? i_input_data[281 % IN_WIDTH] : ping_storage_data_66 ^ i_input_data[281 % IN_WIDTH];
                779 / IN_WIDTH: ping_storage_data_66 <= (fillup_transition == 1'b1) ? i_input_data[779 % IN_WIDTH] : ping_storage_data_66 ^ i_input_data[779 % IN_WIDTH];
                943 / IN_WIDTH: ping_storage_data_66 <= (fillup_transition == 1'b1) ? i_input_data[943 % IN_WIDTH] : ping_storage_data_66 ^ i_input_data[943 % IN_WIDTH];
                default: ping_storage_data_66 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_66;
                endcase
            end else begin
                case (input_count)
                164 / IN_WIDTH: pong_storage_data_66 <= (fillup_transition == 1'b1) ? i_input_data[164 % IN_WIDTH] : pong_storage_data_66 ^ i_input_data[164 % IN_WIDTH];
                281 / IN_WIDTH: pong_storage_data_66 <= (fillup_transition == 1'b1) ? i_input_data[281 % IN_WIDTH] : pong_storage_data_66 ^ i_input_data[281 % IN_WIDTH];
                779 / IN_WIDTH: pong_storage_data_66 <= (fillup_transition == 1'b1) ? i_input_data[779 % IN_WIDTH] : pong_storage_data_66 ^ i_input_data[779 % IN_WIDTH];
                943 / IN_WIDTH: pong_storage_data_66 <= (fillup_transition == 1'b1) ? i_input_data[943 % IN_WIDTH] : pong_storage_data_66 ^ i_input_data[943 % IN_WIDTH];
                default: pong_storage_data_66 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_66;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_66 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_66;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_66 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_66;
            end
        end
    end
end

logic ping_storage_data_67;
logic pong_storage_data_67;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_67 <= 1'b0;
        pong_storage_data_67 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                165 / IN_WIDTH: ping_storage_data_67 <= (fillup_transition == 1'b1) ? i_input_data[165 % IN_WIDTH] : ping_storage_data_67 ^ i_input_data[165 % IN_WIDTH];
                282 / IN_WIDTH: ping_storage_data_67 <= (fillup_transition == 1'b1) ? i_input_data[282 % IN_WIDTH] : ping_storage_data_67 ^ i_input_data[282 % IN_WIDTH];
                780 / IN_WIDTH: ping_storage_data_67 <= (fillup_transition == 1'b1) ? i_input_data[780 % IN_WIDTH] : ping_storage_data_67 ^ i_input_data[780 % IN_WIDTH];
                944 / IN_WIDTH: ping_storage_data_67 <= (fillup_transition == 1'b1) ? i_input_data[944 % IN_WIDTH] : ping_storage_data_67 ^ i_input_data[944 % IN_WIDTH];
                default: ping_storage_data_67 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_67;
                endcase
            end else begin
                case (input_count)
                165 / IN_WIDTH: pong_storage_data_67 <= (fillup_transition == 1'b1) ? i_input_data[165 % IN_WIDTH] : pong_storage_data_67 ^ i_input_data[165 % IN_WIDTH];
                282 / IN_WIDTH: pong_storage_data_67 <= (fillup_transition == 1'b1) ? i_input_data[282 % IN_WIDTH] : pong_storage_data_67 ^ i_input_data[282 % IN_WIDTH];
                780 / IN_WIDTH: pong_storage_data_67 <= (fillup_transition == 1'b1) ? i_input_data[780 % IN_WIDTH] : pong_storage_data_67 ^ i_input_data[780 % IN_WIDTH];
                944 / IN_WIDTH: pong_storage_data_67 <= (fillup_transition == 1'b1) ? i_input_data[944 % IN_WIDTH] : pong_storage_data_67 ^ i_input_data[944 % IN_WIDTH];
                default: pong_storage_data_67 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_67;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_67 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_67;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_67 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_67;
            end
        end
    end
end

logic ping_storage_data_68;
logic pong_storage_data_68;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_68 <= 1'b0;
        pong_storage_data_68 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                166 / IN_WIDTH: ping_storage_data_68 <= (fillup_transition == 1'b1) ? i_input_data[166 % IN_WIDTH] : ping_storage_data_68 ^ i_input_data[166 % IN_WIDTH];
                283 / IN_WIDTH: ping_storage_data_68 <= (fillup_transition == 1'b1) ? i_input_data[283 % IN_WIDTH] : ping_storage_data_68 ^ i_input_data[283 % IN_WIDTH];
                781 / IN_WIDTH: ping_storage_data_68 <= (fillup_transition == 1'b1) ? i_input_data[781 % IN_WIDTH] : ping_storage_data_68 ^ i_input_data[781 % IN_WIDTH];
                945 / IN_WIDTH: ping_storage_data_68 <= (fillup_transition == 1'b1) ? i_input_data[945 % IN_WIDTH] : ping_storage_data_68 ^ i_input_data[945 % IN_WIDTH];
                default: ping_storage_data_68 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_68;
                endcase
            end else begin
                case (input_count)
                166 / IN_WIDTH: pong_storage_data_68 <= (fillup_transition == 1'b1) ? i_input_data[166 % IN_WIDTH] : pong_storage_data_68 ^ i_input_data[166 % IN_WIDTH];
                283 / IN_WIDTH: pong_storage_data_68 <= (fillup_transition == 1'b1) ? i_input_data[283 % IN_WIDTH] : pong_storage_data_68 ^ i_input_data[283 % IN_WIDTH];
                781 / IN_WIDTH: pong_storage_data_68 <= (fillup_transition == 1'b1) ? i_input_data[781 % IN_WIDTH] : pong_storage_data_68 ^ i_input_data[781 % IN_WIDTH];
                945 / IN_WIDTH: pong_storage_data_68 <= (fillup_transition == 1'b1) ? i_input_data[945 % IN_WIDTH] : pong_storage_data_68 ^ i_input_data[945 % IN_WIDTH];
                default: pong_storage_data_68 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_68;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_68 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_68;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_68 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_68;
            end
        end
    end
end

logic ping_storage_data_69;
logic pong_storage_data_69;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_69 <= 1'b0;
        pong_storage_data_69 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                167 / IN_WIDTH: ping_storage_data_69 <= (fillup_transition == 1'b1) ? i_input_data[167 % IN_WIDTH] : ping_storage_data_69 ^ i_input_data[167 % IN_WIDTH];
                284 / IN_WIDTH: ping_storage_data_69 <= (fillup_transition == 1'b1) ? i_input_data[284 % IN_WIDTH] : ping_storage_data_69 ^ i_input_data[284 % IN_WIDTH];
                782 / IN_WIDTH: ping_storage_data_69 <= (fillup_transition == 1'b1) ? i_input_data[782 % IN_WIDTH] : ping_storage_data_69 ^ i_input_data[782 % IN_WIDTH];
                946 / IN_WIDTH: ping_storage_data_69 <= (fillup_transition == 1'b1) ? i_input_data[946 % IN_WIDTH] : ping_storage_data_69 ^ i_input_data[946 % IN_WIDTH];
                default: ping_storage_data_69 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_69;
                endcase
            end else begin
                case (input_count)
                167 / IN_WIDTH: pong_storage_data_69 <= (fillup_transition == 1'b1) ? i_input_data[167 % IN_WIDTH] : pong_storage_data_69 ^ i_input_data[167 % IN_WIDTH];
                284 / IN_WIDTH: pong_storage_data_69 <= (fillup_transition == 1'b1) ? i_input_data[284 % IN_WIDTH] : pong_storage_data_69 ^ i_input_data[284 % IN_WIDTH];
                782 / IN_WIDTH: pong_storage_data_69 <= (fillup_transition == 1'b1) ? i_input_data[782 % IN_WIDTH] : pong_storage_data_69 ^ i_input_data[782 % IN_WIDTH];
                946 / IN_WIDTH: pong_storage_data_69 <= (fillup_transition == 1'b1) ? i_input_data[946 % IN_WIDTH] : pong_storage_data_69 ^ i_input_data[946 % IN_WIDTH];
                default: pong_storage_data_69 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_69;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_69 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_69;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_69 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_69;
            end
        end
    end
end

logic ping_storage_data_70;
logic pong_storage_data_70;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_70 <= 1'b0;
        pong_storage_data_70 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                168 / IN_WIDTH: ping_storage_data_70 <= (fillup_transition == 1'b1) ? i_input_data[168 % IN_WIDTH] : ping_storage_data_70 ^ i_input_data[168 % IN_WIDTH];
                285 / IN_WIDTH: ping_storage_data_70 <= (fillup_transition == 1'b1) ? i_input_data[285 % IN_WIDTH] : ping_storage_data_70 ^ i_input_data[285 % IN_WIDTH];
                783 / IN_WIDTH: ping_storage_data_70 <= (fillup_transition == 1'b1) ? i_input_data[783 % IN_WIDTH] : ping_storage_data_70 ^ i_input_data[783 % IN_WIDTH];
                947 / IN_WIDTH: ping_storage_data_70 <= (fillup_transition == 1'b1) ? i_input_data[947 % IN_WIDTH] : ping_storage_data_70 ^ i_input_data[947 % IN_WIDTH];
                default: ping_storage_data_70 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_70;
                endcase
            end else begin
                case (input_count)
                168 / IN_WIDTH: pong_storage_data_70 <= (fillup_transition == 1'b1) ? i_input_data[168 % IN_WIDTH] : pong_storage_data_70 ^ i_input_data[168 % IN_WIDTH];
                285 / IN_WIDTH: pong_storage_data_70 <= (fillup_transition == 1'b1) ? i_input_data[285 % IN_WIDTH] : pong_storage_data_70 ^ i_input_data[285 % IN_WIDTH];
                783 / IN_WIDTH: pong_storage_data_70 <= (fillup_transition == 1'b1) ? i_input_data[783 % IN_WIDTH] : pong_storage_data_70 ^ i_input_data[783 % IN_WIDTH];
                947 / IN_WIDTH: pong_storage_data_70 <= (fillup_transition == 1'b1) ? i_input_data[947 % IN_WIDTH] : pong_storage_data_70 ^ i_input_data[947 % IN_WIDTH];
                default: pong_storage_data_70 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_70;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_70 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_70;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_70 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_70;
            end
        end
    end
end

logic ping_storage_data_71;
logic pong_storage_data_71;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_71 <= 1'b0;
        pong_storage_data_71 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                169 / IN_WIDTH: ping_storage_data_71 <= (fillup_transition == 1'b1) ? i_input_data[169 % IN_WIDTH] : ping_storage_data_71 ^ i_input_data[169 % IN_WIDTH];
                286 / IN_WIDTH: ping_storage_data_71 <= (fillup_transition == 1'b1) ? i_input_data[286 % IN_WIDTH] : ping_storage_data_71 ^ i_input_data[286 % IN_WIDTH];
                784 / IN_WIDTH: ping_storage_data_71 <= (fillup_transition == 1'b1) ? i_input_data[784 % IN_WIDTH] : ping_storage_data_71 ^ i_input_data[784 % IN_WIDTH];
                948 / IN_WIDTH: ping_storage_data_71 <= (fillup_transition == 1'b1) ? i_input_data[948 % IN_WIDTH] : ping_storage_data_71 ^ i_input_data[948 % IN_WIDTH];
                default: ping_storage_data_71 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_71;
                endcase
            end else begin
                case (input_count)
                169 / IN_WIDTH: pong_storage_data_71 <= (fillup_transition == 1'b1) ? i_input_data[169 % IN_WIDTH] : pong_storage_data_71 ^ i_input_data[169 % IN_WIDTH];
                286 / IN_WIDTH: pong_storage_data_71 <= (fillup_transition == 1'b1) ? i_input_data[286 % IN_WIDTH] : pong_storage_data_71 ^ i_input_data[286 % IN_WIDTH];
                784 / IN_WIDTH: pong_storage_data_71 <= (fillup_transition == 1'b1) ? i_input_data[784 % IN_WIDTH] : pong_storage_data_71 ^ i_input_data[784 % IN_WIDTH];
                948 / IN_WIDTH: pong_storage_data_71 <= (fillup_transition == 1'b1) ? i_input_data[948 % IN_WIDTH] : pong_storage_data_71 ^ i_input_data[948 % IN_WIDTH];
                default: pong_storage_data_71 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_71;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_71 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_71;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_71 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_71;
            end
        end
    end
end

logic ping_storage_data_72;
logic pong_storage_data_72;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_72 <= 1'b0;
        pong_storage_data_72 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                170 / IN_WIDTH: ping_storage_data_72 <= (fillup_transition == 1'b1) ? i_input_data[170 % IN_WIDTH] : ping_storage_data_72 ^ i_input_data[170 % IN_WIDTH];
                287 / IN_WIDTH: ping_storage_data_72 <= (fillup_transition == 1'b1) ? i_input_data[287 % IN_WIDTH] : ping_storage_data_72 ^ i_input_data[287 % IN_WIDTH];
                785 / IN_WIDTH: ping_storage_data_72 <= (fillup_transition == 1'b1) ? i_input_data[785 % IN_WIDTH] : ping_storage_data_72 ^ i_input_data[785 % IN_WIDTH];
                949 / IN_WIDTH: ping_storage_data_72 <= (fillup_transition == 1'b1) ? i_input_data[949 % IN_WIDTH] : ping_storage_data_72 ^ i_input_data[949 % IN_WIDTH];
                default: ping_storage_data_72 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_72;
                endcase
            end else begin
                case (input_count)
                170 / IN_WIDTH: pong_storage_data_72 <= (fillup_transition == 1'b1) ? i_input_data[170 % IN_WIDTH] : pong_storage_data_72 ^ i_input_data[170 % IN_WIDTH];
                287 / IN_WIDTH: pong_storage_data_72 <= (fillup_transition == 1'b1) ? i_input_data[287 % IN_WIDTH] : pong_storage_data_72 ^ i_input_data[287 % IN_WIDTH];
                785 / IN_WIDTH: pong_storage_data_72 <= (fillup_transition == 1'b1) ? i_input_data[785 % IN_WIDTH] : pong_storage_data_72 ^ i_input_data[785 % IN_WIDTH];
                949 / IN_WIDTH: pong_storage_data_72 <= (fillup_transition == 1'b1) ? i_input_data[949 % IN_WIDTH] : pong_storage_data_72 ^ i_input_data[949 % IN_WIDTH];
                default: pong_storage_data_72 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_72;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_72 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_72;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_72 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_72;
            end
        end
    end
end

logic ping_storage_data_73;
logic pong_storage_data_73;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_73 <= 1'b0;
        pong_storage_data_73 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                171 / IN_WIDTH: ping_storage_data_73 <= (fillup_transition == 1'b1) ? i_input_data[171 % IN_WIDTH] : ping_storage_data_73 ^ i_input_data[171 % IN_WIDTH];
                192 / IN_WIDTH: ping_storage_data_73 <= (fillup_transition == 1'b1) ? i_input_data[192 % IN_WIDTH] : ping_storage_data_73 ^ i_input_data[192 % IN_WIDTH];
                786 / IN_WIDTH: ping_storage_data_73 <= (fillup_transition == 1'b1) ? i_input_data[786 % IN_WIDTH] : ping_storage_data_73 ^ i_input_data[786 % IN_WIDTH];
                950 / IN_WIDTH: ping_storage_data_73 <= (fillup_transition == 1'b1) ? i_input_data[950 % IN_WIDTH] : ping_storage_data_73 ^ i_input_data[950 % IN_WIDTH];
                default: ping_storage_data_73 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_73;
                endcase
            end else begin
                case (input_count)
                171 / IN_WIDTH: pong_storage_data_73 <= (fillup_transition == 1'b1) ? i_input_data[171 % IN_WIDTH] : pong_storage_data_73 ^ i_input_data[171 % IN_WIDTH];
                192 / IN_WIDTH: pong_storage_data_73 <= (fillup_transition == 1'b1) ? i_input_data[192 % IN_WIDTH] : pong_storage_data_73 ^ i_input_data[192 % IN_WIDTH];
                786 / IN_WIDTH: pong_storage_data_73 <= (fillup_transition == 1'b1) ? i_input_data[786 % IN_WIDTH] : pong_storage_data_73 ^ i_input_data[786 % IN_WIDTH];
                950 / IN_WIDTH: pong_storage_data_73 <= (fillup_transition == 1'b1) ? i_input_data[950 % IN_WIDTH] : pong_storage_data_73 ^ i_input_data[950 % IN_WIDTH];
                default: pong_storage_data_73 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_73;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_73 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_73;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_73 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_73;
            end
        end
    end
end

logic ping_storage_data_74;
logic pong_storage_data_74;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_74 <= 1'b0;
        pong_storage_data_74 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                172 / IN_WIDTH: ping_storage_data_74 <= (fillup_transition == 1'b1) ? i_input_data[172 % IN_WIDTH] : ping_storage_data_74 ^ i_input_data[172 % IN_WIDTH];
                193 / IN_WIDTH: ping_storage_data_74 <= (fillup_transition == 1'b1) ? i_input_data[193 % IN_WIDTH] : ping_storage_data_74 ^ i_input_data[193 % IN_WIDTH];
                787 / IN_WIDTH: ping_storage_data_74 <= (fillup_transition == 1'b1) ? i_input_data[787 % IN_WIDTH] : ping_storage_data_74 ^ i_input_data[787 % IN_WIDTH];
                951 / IN_WIDTH: ping_storage_data_74 <= (fillup_transition == 1'b1) ? i_input_data[951 % IN_WIDTH] : ping_storage_data_74 ^ i_input_data[951 % IN_WIDTH];
                default: ping_storage_data_74 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_74;
                endcase
            end else begin
                case (input_count)
                172 / IN_WIDTH: pong_storage_data_74 <= (fillup_transition == 1'b1) ? i_input_data[172 % IN_WIDTH] : pong_storage_data_74 ^ i_input_data[172 % IN_WIDTH];
                193 / IN_WIDTH: pong_storage_data_74 <= (fillup_transition == 1'b1) ? i_input_data[193 % IN_WIDTH] : pong_storage_data_74 ^ i_input_data[193 % IN_WIDTH];
                787 / IN_WIDTH: pong_storage_data_74 <= (fillup_transition == 1'b1) ? i_input_data[787 % IN_WIDTH] : pong_storage_data_74 ^ i_input_data[787 % IN_WIDTH];
                951 / IN_WIDTH: pong_storage_data_74 <= (fillup_transition == 1'b1) ? i_input_data[951 % IN_WIDTH] : pong_storage_data_74 ^ i_input_data[951 % IN_WIDTH];
                default: pong_storage_data_74 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_74;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_74 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_74;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_74 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_74;
            end
        end
    end
end

logic ping_storage_data_75;
logic pong_storage_data_75;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_75 <= 1'b0;
        pong_storage_data_75 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                173 / IN_WIDTH: ping_storage_data_75 <= (fillup_transition == 1'b1) ? i_input_data[173 % IN_WIDTH] : ping_storage_data_75 ^ i_input_data[173 % IN_WIDTH];
                194 / IN_WIDTH: ping_storage_data_75 <= (fillup_transition == 1'b1) ? i_input_data[194 % IN_WIDTH] : ping_storage_data_75 ^ i_input_data[194 % IN_WIDTH];
                788 / IN_WIDTH: ping_storage_data_75 <= (fillup_transition == 1'b1) ? i_input_data[788 % IN_WIDTH] : ping_storage_data_75 ^ i_input_data[788 % IN_WIDTH];
                952 / IN_WIDTH: ping_storage_data_75 <= (fillup_transition == 1'b1) ? i_input_data[952 % IN_WIDTH] : ping_storage_data_75 ^ i_input_data[952 % IN_WIDTH];
                default: ping_storage_data_75 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_75;
                endcase
            end else begin
                case (input_count)
                173 / IN_WIDTH: pong_storage_data_75 <= (fillup_transition == 1'b1) ? i_input_data[173 % IN_WIDTH] : pong_storage_data_75 ^ i_input_data[173 % IN_WIDTH];
                194 / IN_WIDTH: pong_storage_data_75 <= (fillup_transition == 1'b1) ? i_input_data[194 % IN_WIDTH] : pong_storage_data_75 ^ i_input_data[194 % IN_WIDTH];
                788 / IN_WIDTH: pong_storage_data_75 <= (fillup_transition == 1'b1) ? i_input_data[788 % IN_WIDTH] : pong_storage_data_75 ^ i_input_data[788 % IN_WIDTH];
                952 / IN_WIDTH: pong_storage_data_75 <= (fillup_transition == 1'b1) ? i_input_data[952 % IN_WIDTH] : pong_storage_data_75 ^ i_input_data[952 % IN_WIDTH];
                default: pong_storage_data_75 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_75;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_75 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_75;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_75 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_75;
            end
        end
    end
end

logic ping_storage_data_76;
logic pong_storage_data_76;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_76 <= 1'b0;
        pong_storage_data_76 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                174 / IN_WIDTH: ping_storage_data_76 <= (fillup_transition == 1'b1) ? i_input_data[174 % IN_WIDTH] : ping_storage_data_76 ^ i_input_data[174 % IN_WIDTH];
                195 / IN_WIDTH: ping_storage_data_76 <= (fillup_transition == 1'b1) ? i_input_data[195 % IN_WIDTH] : ping_storage_data_76 ^ i_input_data[195 % IN_WIDTH];
                789 / IN_WIDTH: ping_storage_data_76 <= (fillup_transition == 1'b1) ? i_input_data[789 % IN_WIDTH] : ping_storage_data_76 ^ i_input_data[789 % IN_WIDTH];
                953 / IN_WIDTH: ping_storage_data_76 <= (fillup_transition == 1'b1) ? i_input_data[953 % IN_WIDTH] : ping_storage_data_76 ^ i_input_data[953 % IN_WIDTH];
                default: ping_storage_data_76 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_76;
                endcase
            end else begin
                case (input_count)
                174 / IN_WIDTH: pong_storage_data_76 <= (fillup_transition == 1'b1) ? i_input_data[174 % IN_WIDTH] : pong_storage_data_76 ^ i_input_data[174 % IN_WIDTH];
                195 / IN_WIDTH: pong_storage_data_76 <= (fillup_transition == 1'b1) ? i_input_data[195 % IN_WIDTH] : pong_storage_data_76 ^ i_input_data[195 % IN_WIDTH];
                789 / IN_WIDTH: pong_storage_data_76 <= (fillup_transition == 1'b1) ? i_input_data[789 % IN_WIDTH] : pong_storage_data_76 ^ i_input_data[789 % IN_WIDTH];
                953 / IN_WIDTH: pong_storage_data_76 <= (fillup_transition == 1'b1) ? i_input_data[953 % IN_WIDTH] : pong_storage_data_76 ^ i_input_data[953 % IN_WIDTH];
                default: pong_storage_data_76 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_76;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_76 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_76;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_76 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_76;
            end
        end
    end
end

logic ping_storage_data_77;
logic pong_storage_data_77;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_77 <= 1'b0;
        pong_storage_data_77 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                175 / IN_WIDTH: ping_storage_data_77 <= (fillup_transition == 1'b1) ? i_input_data[175 % IN_WIDTH] : ping_storage_data_77 ^ i_input_data[175 % IN_WIDTH];
                196 / IN_WIDTH: ping_storage_data_77 <= (fillup_transition == 1'b1) ? i_input_data[196 % IN_WIDTH] : ping_storage_data_77 ^ i_input_data[196 % IN_WIDTH];
                790 / IN_WIDTH: ping_storage_data_77 <= (fillup_transition == 1'b1) ? i_input_data[790 % IN_WIDTH] : ping_storage_data_77 ^ i_input_data[790 % IN_WIDTH];
                954 / IN_WIDTH: ping_storage_data_77 <= (fillup_transition == 1'b1) ? i_input_data[954 % IN_WIDTH] : ping_storage_data_77 ^ i_input_data[954 % IN_WIDTH];
                default: ping_storage_data_77 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_77;
                endcase
            end else begin
                case (input_count)
                175 / IN_WIDTH: pong_storage_data_77 <= (fillup_transition == 1'b1) ? i_input_data[175 % IN_WIDTH] : pong_storage_data_77 ^ i_input_data[175 % IN_WIDTH];
                196 / IN_WIDTH: pong_storage_data_77 <= (fillup_transition == 1'b1) ? i_input_data[196 % IN_WIDTH] : pong_storage_data_77 ^ i_input_data[196 % IN_WIDTH];
                790 / IN_WIDTH: pong_storage_data_77 <= (fillup_transition == 1'b1) ? i_input_data[790 % IN_WIDTH] : pong_storage_data_77 ^ i_input_data[790 % IN_WIDTH];
                954 / IN_WIDTH: pong_storage_data_77 <= (fillup_transition == 1'b1) ? i_input_data[954 % IN_WIDTH] : pong_storage_data_77 ^ i_input_data[954 % IN_WIDTH];
                default: pong_storage_data_77 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_77;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_77 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_77;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_77 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_77;
            end
        end
    end
end

logic ping_storage_data_78;
logic pong_storage_data_78;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_78 <= 1'b0;
        pong_storage_data_78 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                176 / IN_WIDTH: ping_storage_data_78 <= (fillup_transition == 1'b1) ? i_input_data[176 % IN_WIDTH] : ping_storage_data_78 ^ i_input_data[176 % IN_WIDTH];
                197 / IN_WIDTH: ping_storage_data_78 <= (fillup_transition == 1'b1) ? i_input_data[197 % IN_WIDTH] : ping_storage_data_78 ^ i_input_data[197 % IN_WIDTH];
                791 / IN_WIDTH: ping_storage_data_78 <= (fillup_transition == 1'b1) ? i_input_data[791 % IN_WIDTH] : ping_storage_data_78 ^ i_input_data[791 % IN_WIDTH];
                955 / IN_WIDTH: ping_storage_data_78 <= (fillup_transition == 1'b1) ? i_input_data[955 % IN_WIDTH] : ping_storage_data_78 ^ i_input_data[955 % IN_WIDTH];
                default: ping_storage_data_78 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_78;
                endcase
            end else begin
                case (input_count)
                176 / IN_WIDTH: pong_storage_data_78 <= (fillup_transition == 1'b1) ? i_input_data[176 % IN_WIDTH] : pong_storage_data_78 ^ i_input_data[176 % IN_WIDTH];
                197 / IN_WIDTH: pong_storage_data_78 <= (fillup_transition == 1'b1) ? i_input_data[197 % IN_WIDTH] : pong_storage_data_78 ^ i_input_data[197 % IN_WIDTH];
                791 / IN_WIDTH: pong_storage_data_78 <= (fillup_transition == 1'b1) ? i_input_data[791 % IN_WIDTH] : pong_storage_data_78 ^ i_input_data[791 % IN_WIDTH];
                955 / IN_WIDTH: pong_storage_data_78 <= (fillup_transition == 1'b1) ? i_input_data[955 % IN_WIDTH] : pong_storage_data_78 ^ i_input_data[955 % IN_WIDTH];
                default: pong_storage_data_78 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_78;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_78 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_78;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_78 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_78;
            end
        end
    end
end

logic ping_storage_data_79;
logic pong_storage_data_79;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_79 <= 1'b0;
        pong_storage_data_79 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                177 / IN_WIDTH: ping_storage_data_79 <= (fillup_transition == 1'b1) ? i_input_data[177 % IN_WIDTH] : ping_storage_data_79 ^ i_input_data[177 % IN_WIDTH];
                198 / IN_WIDTH: ping_storage_data_79 <= (fillup_transition == 1'b1) ? i_input_data[198 % IN_WIDTH] : ping_storage_data_79 ^ i_input_data[198 % IN_WIDTH];
                792 / IN_WIDTH: ping_storage_data_79 <= (fillup_transition == 1'b1) ? i_input_data[792 % IN_WIDTH] : ping_storage_data_79 ^ i_input_data[792 % IN_WIDTH];
                956 / IN_WIDTH: ping_storage_data_79 <= (fillup_transition == 1'b1) ? i_input_data[956 % IN_WIDTH] : ping_storage_data_79 ^ i_input_data[956 % IN_WIDTH];
                default: ping_storage_data_79 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_79;
                endcase
            end else begin
                case (input_count)
                177 / IN_WIDTH: pong_storage_data_79 <= (fillup_transition == 1'b1) ? i_input_data[177 % IN_WIDTH] : pong_storage_data_79 ^ i_input_data[177 % IN_WIDTH];
                198 / IN_WIDTH: pong_storage_data_79 <= (fillup_transition == 1'b1) ? i_input_data[198 % IN_WIDTH] : pong_storage_data_79 ^ i_input_data[198 % IN_WIDTH];
                792 / IN_WIDTH: pong_storage_data_79 <= (fillup_transition == 1'b1) ? i_input_data[792 % IN_WIDTH] : pong_storage_data_79 ^ i_input_data[792 % IN_WIDTH];
                956 / IN_WIDTH: pong_storage_data_79 <= (fillup_transition == 1'b1) ? i_input_data[956 % IN_WIDTH] : pong_storage_data_79 ^ i_input_data[956 % IN_WIDTH];
                default: pong_storage_data_79 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_79;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_79 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_79;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_79 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_79;
            end
        end
    end
end

logic ping_storage_data_80;
logic pong_storage_data_80;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_80 <= 1'b0;
        pong_storage_data_80 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                178 / IN_WIDTH: ping_storage_data_80 <= (fillup_transition == 1'b1) ? i_input_data[178 % IN_WIDTH] : ping_storage_data_80 ^ i_input_data[178 % IN_WIDTH];
                199 / IN_WIDTH: ping_storage_data_80 <= (fillup_transition == 1'b1) ? i_input_data[199 % IN_WIDTH] : ping_storage_data_80 ^ i_input_data[199 % IN_WIDTH];
                793 / IN_WIDTH: ping_storage_data_80 <= (fillup_transition == 1'b1) ? i_input_data[793 % IN_WIDTH] : ping_storage_data_80 ^ i_input_data[793 % IN_WIDTH];
                957 / IN_WIDTH: ping_storage_data_80 <= (fillup_transition == 1'b1) ? i_input_data[957 % IN_WIDTH] : ping_storage_data_80 ^ i_input_data[957 % IN_WIDTH];
                default: ping_storage_data_80 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_80;
                endcase
            end else begin
                case (input_count)
                178 / IN_WIDTH: pong_storage_data_80 <= (fillup_transition == 1'b1) ? i_input_data[178 % IN_WIDTH] : pong_storage_data_80 ^ i_input_data[178 % IN_WIDTH];
                199 / IN_WIDTH: pong_storage_data_80 <= (fillup_transition == 1'b1) ? i_input_data[199 % IN_WIDTH] : pong_storage_data_80 ^ i_input_data[199 % IN_WIDTH];
                793 / IN_WIDTH: pong_storage_data_80 <= (fillup_transition == 1'b1) ? i_input_data[793 % IN_WIDTH] : pong_storage_data_80 ^ i_input_data[793 % IN_WIDTH];
                957 / IN_WIDTH: pong_storage_data_80 <= (fillup_transition == 1'b1) ? i_input_data[957 % IN_WIDTH] : pong_storage_data_80 ^ i_input_data[957 % IN_WIDTH];
                default: pong_storage_data_80 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_80;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_80 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_80;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_80 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_80;
            end
        end
    end
end

logic ping_storage_data_81;
logic pong_storage_data_81;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_81 <= 1'b0;
        pong_storage_data_81 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                179 / IN_WIDTH: ping_storage_data_81 <= (fillup_transition == 1'b1) ? i_input_data[179 % IN_WIDTH] : ping_storage_data_81 ^ i_input_data[179 % IN_WIDTH];
                200 / IN_WIDTH: ping_storage_data_81 <= (fillup_transition == 1'b1) ? i_input_data[200 % IN_WIDTH] : ping_storage_data_81 ^ i_input_data[200 % IN_WIDTH];
                794 / IN_WIDTH: ping_storage_data_81 <= (fillup_transition == 1'b1) ? i_input_data[794 % IN_WIDTH] : ping_storage_data_81 ^ i_input_data[794 % IN_WIDTH];
                958 / IN_WIDTH: ping_storage_data_81 <= (fillup_transition == 1'b1) ? i_input_data[958 % IN_WIDTH] : ping_storage_data_81 ^ i_input_data[958 % IN_WIDTH];
                default: ping_storage_data_81 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_81;
                endcase
            end else begin
                case (input_count)
                179 / IN_WIDTH: pong_storage_data_81 <= (fillup_transition == 1'b1) ? i_input_data[179 % IN_WIDTH] : pong_storage_data_81 ^ i_input_data[179 % IN_WIDTH];
                200 / IN_WIDTH: pong_storage_data_81 <= (fillup_transition == 1'b1) ? i_input_data[200 % IN_WIDTH] : pong_storage_data_81 ^ i_input_data[200 % IN_WIDTH];
                794 / IN_WIDTH: pong_storage_data_81 <= (fillup_transition == 1'b1) ? i_input_data[794 % IN_WIDTH] : pong_storage_data_81 ^ i_input_data[794 % IN_WIDTH];
                958 / IN_WIDTH: pong_storage_data_81 <= (fillup_transition == 1'b1) ? i_input_data[958 % IN_WIDTH] : pong_storage_data_81 ^ i_input_data[958 % IN_WIDTH];
                default: pong_storage_data_81 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_81;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_81 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_81;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_81 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_81;
            end
        end
    end
end

logic ping_storage_data_82;
logic pong_storage_data_82;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_82 <= 1'b0;
        pong_storage_data_82 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                180 / IN_WIDTH: ping_storage_data_82 <= (fillup_transition == 1'b1) ? i_input_data[180 % IN_WIDTH] : ping_storage_data_82 ^ i_input_data[180 % IN_WIDTH];
                201 / IN_WIDTH: ping_storage_data_82 <= (fillup_transition == 1'b1) ? i_input_data[201 % IN_WIDTH] : ping_storage_data_82 ^ i_input_data[201 % IN_WIDTH];
                795 / IN_WIDTH: ping_storage_data_82 <= (fillup_transition == 1'b1) ? i_input_data[795 % IN_WIDTH] : ping_storage_data_82 ^ i_input_data[795 % IN_WIDTH];
                959 / IN_WIDTH: ping_storage_data_82 <= (fillup_transition == 1'b1) ? i_input_data[959 % IN_WIDTH] : ping_storage_data_82 ^ i_input_data[959 % IN_WIDTH];
                default: ping_storage_data_82 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_82;
                endcase
            end else begin
                case (input_count)
                180 / IN_WIDTH: pong_storage_data_82 <= (fillup_transition == 1'b1) ? i_input_data[180 % IN_WIDTH] : pong_storage_data_82 ^ i_input_data[180 % IN_WIDTH];
                201 / IN_WIDTH: pong_storage_data_82 <= (fillup_transition == 1'b1) ? i_input_data[201 % IN_WIDTH] : pong_storage_data_82 ^ i_input_data[201 % IN_WIDTH];
                795 / IN_WIDTH: pong_storage_data_82 <= (fillup_transition == 1'b1) ? i_input_data[795 % IN_WIDTH] : pong_storage_data_82 ^ i_input_data[795 % IN_WIDTH];
                959 / IN_WIDTH: pong_storage_data_82 <= (fillup_transition == 1'b1) ? i_input_data[959 % IN_WIDTH] : pong_storage_data_82 ^ i_input_data[959 % IN_WIDTH];
                default: pong_storage_data_82 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_82;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_82 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_82;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_82 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_82;
            end
        end
    end
end

logic ping_storage_data_83;
logic pong_storage_data_83;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_83 <= 1'b0;
        pong_storage_data_83 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                181 / IN_WIDTH: ping_storage_data_83 <= (fillup_transition == 1'b1) ? i_input_data[181 % IN_WIDTH] : ping_storage_data_83 ^ i_input_data[181 % IN_WIDTH];
                202 / IN_WIDTH: ping_storage_data_83 <= (fillup_transition == 1'b1) ? i_input_data[202 % IN_WIDTH] : ping_storage_data_83 ^ i_input_data[202 % IN_WIDTH];
                796 / IN_WIDTH: ping_storage_data_83 <= (fillup_transition == 1'b1) ? i_input_data[796 % IN_WIDTH] : ping_storage_data_83 ^ i_input_data[796 % IN_WIDTH];
                864 / IN_WIDTH: ping_storage_data_83 <= (fillup_transition == 1'b1) ? i_input_data[864 % IN_WIDTH] : ping_storage_data_83 ^ i_input_data[864 % IN_WIDTH];
                default: ping_storage_data_83 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_83;
                endcase
            end else begin
                case (input_count)
                181 / IN_WIDTH: pong_storage_data_83 <= (fillup_transition == 1'b1) ? i_input_data[181 % IN_WIDTH] : pong_storage_data_83 ^ i_input_data[181 % IN_WIDTH];
                202 / IN_WIDTH: pong_storage_data_83 <= (fillup_transition == 1'b1) ? i_input_data[202 % IN_WIDTH] : pong_storage_data_83 ^ i_input_data[202 % IN_WIDTH];
                796 / IN_WIDTH: pong_storage_data_83 <= (fillup_transition == 1'b1) ? i_input_data[796 % IN_WIDTH] : pong_storage_data_83 ^ i_input_data[796 % IN_WIDTH];
                864 / IN_WIDTH: pong_storage_data_83 <= (fillup_transition == 1'b1) ? i_input_data[864 % IN_WIDTH] : pong_storage_data_83 ^ i_input_data[864 % IN_WIDTH];
                default: pong_storage_data_83 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_83;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_83 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_83;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_83 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_83;
            end
        end
    end
end

logic ping_storage_data_84;
logic pong_storage_data_84;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_84 <= 1'b0;
        pong_storage_data_84 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                182 / IN_WIDTH: ping_storage_data_84 <= (fillup_transition == 1'b1) ? i_input_data[182 % IN_WIDTH] : ping_storage_data_84 ^ i_input_data[182 % IN_WIDTH];
                203 / IN_WIDTH: ping_storage_data_84 <= (fillup_transition == 1'b1) ? i_input_data[203 % IN_WIDTH] : ping_storage_data_84 ^ i_input_data[203 % IN_WIDTH];
                797 / IN_WIDTH: ping_storage_data_84 <= (fillup_transition == 1'b1) ? i_input_data[797 % IN_WIDTH] : ping_storage_data_84 ^ i_input_data[797 % IN_WIDTH];
                865 / IN_WIDTH: ping_storage_data_84 <= (fillup_transition == 1'b1) ? i_input_data[865 % IN_WIDTH] : ping_storage_data_84 ^ i_input_data[865 % IN_WIDTH];
                default: ping_storage_data_84 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_84;
                endcase
            end else begin
                case (input_count)
                182 / IN_WIDTH: pong_storage_data_84 <= (fillup_transition == 1'b1) ? i_input_data[182 % IN_WIDTH] : pong_storage_data_84 ^ i_input_data[182 % IN_WIDTH];
                203 / IN_WIDTH: pong_storage_data_84 <= (fillup_transition == 1'b1) ? i_input_data[203 % IN_WIDTH] : pong_storage_data_84 ^ i_input_data[203 % IN_WIDTH];
                797 / IN_WIDTH: pong_storage_data_84 <= (fillup_transition == 1'b1) ? i_input_data[797 % IN_WIDTH] : pong_storage_data_84 ^ i_input_data[797 % IN_WIDTH];
                865 / IN_WIDTH: pong_storage_data_84 <= (fillup_transition == 1'b1) ? i_input_data[865 % IN_WIDTH] : pong_storage_data_84 ^ i_input_data[865 % IN_WIDTH];
                default: pong_storage_data_84 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_84;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_84 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_84;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_84 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_84;
            end
        end
    end
end

logic ping_storage_data_85;
logic pong_storage_data_85;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_85 <= 1'b0;
        pong_storage_data_85 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                183 / IN_WIDTH: ping_storage_data_85 <= (fillup_transition == 1'b1) ? i_input_data[183 % IN_WIDTH] : ping_storage_data_85 ^ i_input_data[183 % IN_WIDTH];
                204 / IN_WIDTH: ping_storage_data_85 <= (fillup_transition == 1'b1) ? i_input_data[204 % IN_WIDTH] : ping_storage_data_85 ^ i_input_data[204 % IN_WIDTH];
                798 / IN_WIDTH: ping_storage_data_85 <= (fillup_transition == 1'b1) ? i_input_data[798 % IN_WIDTH] : ping_storage_data_85 ^ i_input_data[798 % IN_WIDTH];
                866 / IN_WIDTH: ping_storage_data_85 <= (fillup_transition == 1'b1) ? i_input_data[866 % IN_WIDTH] : ping_storage_data_85 ^ i_input_data[866 % IN_WIDTH];
                default: ping_storage_data_85 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_85;
                endcase
            end else begin
                case (input_count)
                183 / IN_WIDTH: pong_storage_data_85 <= (fillup_transition == 1'b1) ? i_input_data[183 % IN_WIDTH] : pong_storage_data_85 ^ i_input_data[183 % IN_WIDTH];
                204 / IN_WIDTH: pong_storage_data_85 <= (fillup_transition == 1'b1) ? i_input_data[204 % IN_WIDTH] : pong_storage_data_85 ^ i_input_data[204 % IN_WIDTH];
                798 / IN_WIDTH: pong_storage_data_85 <= (fillup_transition == 1'b1) ? i_input_data[798 % IN_WIDTH] : pong_storage_data_85 ^ i_input_data[798 % IN_WIDTH];
                866 / IN_WIDTH: pong_storage_data_85 <= (fillup_transition == 1'b1) ? i_input_data[866 % IN_WIDTH] : pong_storage_data_85 ^ i_input_data[866 % IN_WIDTH];
                default: pong_storage_data_85 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_85;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_85 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_85;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_85 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_85;
            end
        end
    end
end

logic ping_storage_data_86;
logic pong_storage_data_86;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_86 <= 1'b0;
        pong_storage_data_86 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                184 / IN_WIDTH: ping_storage_data_86 <= (fillup_transition == 1'b1) ? i_input_data[184 % IN_WIDTH] : ping_storage_data_86 ^ i_input_data[184 % IN_WIDTH];
                205 / IN_WIDTH: ping_storage_data_86 <= (fillup_transition == 1'b1) ? i_input_data[205 % IN_WIDTH] : ping_storage_data_86 ^ i_input_data[205 % IN_WIDTH];
                799 / IN_WIDTH: ping_storage_data_86 <= (fillup_transition == 1'b1) ? i_input_data[799 % IN_WIDTH] : ping_storage_data_86 ^ i_input_data[799 % IN_WIDTH];
                867 / IN_WIDTH: ping_storage_data_86 <= (fillup_transition == 1'b1) ? i_input_data[867 % IN_WIDTH] : ping_storage_data_86 ^ i_input_data[867 % IN_WIDTH];
                default: ping_storage_data_86 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_86;
                endcase
            end else begin
                case (input_count)
                184 / IN_WIDTH: pong_storage_data_86 <= (fillup_transition == 1'b1) ? i_input_data[184 % IN_WIDTH] : pong_storage_data_86 ^ i_input_data[184 % IN_WIDTH];
                205 / IN_WIDTH: pong_storage_data_86 <= (fillup_transition == 1'b1) ? i_input_data[205 % IN_WIDTH] : pong_storage_data_86 ^ i_input_data[205 % IN_WIDTH];
                799 / IN_WIDTH: pong_storage_data_86 <= (fillup_transition == 1'b1) ? i_input_data[799 % IN_WIDTH] : pong_storage_data_86 ^ i_input_data[799 % IN_WIDTH];
                867 / IN_WIDTH: pong_storage_data_86 <= (fillup_transition == 1'b1) ? i_input_data[867 % IN_WIDTH] : pong_storage_data_86 ^ i_input_data[867 % IN_WIDTH];
                default: pong_storage_data_86 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_86;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_86 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_86;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_86 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_86;
            end
        end
    end
end

logic ping_storage_data_87;
logic pong_storage_data_87;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_87 <= 1'b0;
        pong_storage_data_87 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                185 / IN_WIDTH: ping_storage_data_87 <= (fillup_transition == 1'b1) ? i_input_data[185 % IN_WIDTH] : ping_storage_data_87 ^ i_input_data[185 % IN_WIDTH];
                206 / IN_WIDTH: ping_storage_data_87 <= (fillup_transition == 1'b1) ? i_input_data[206 % IN_WIDTH] : ping_storage_data_87 ^ i_input_data[206 % IN_WIDTH];
                800 / IN_WIDTH: ping_storage_data_87 <= (fillup_transition == 1'b1) ? i_input_data[800 % IN_WIDTH] : ping_storage_data_87 ^ i_input_data[800 % IN_WIDTH];
                868 / IN_WIDTH: ping_storage_data_87 <= (fillup_transition == 1'b1) ? i_input_data[868 % IN_WIDTH] : ping_storage_data_87 ^ i_input_data[868 % IN_WIDTH];
                default: ping_storage_data_87 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_87;
                endcase
            end else begin
                case (input_count)
                185 / IN_WIDTH: pong_storage_data_87 <= (fillup_transition == 1'b1) ? i_input_data[185 % IN_WIDTH] : pong_storage_data_87 ^ i_input_data[185 % IN_WIDTH];
                206 / IN_WIDTH: pong_storage_data_87 <= (fillup_transition == 1'b1) ? i_input_data[206 % IN_WIDTH] : pong_storage_data_87 ^ i_input_data[206 % IN_WIDTH];
                800 / IN_WIDTH: pong_storage_data_87 <= (fillup_transition == 1'b1) ? i_input_data[800 % IN_WIDTH] : pong_storage_data_87 ^ i_input_data[800 % IN_WIDTH];
                868 / IN_WIDTH: pong_storage_data_87 <= (fillup_transition == 1'b1) ? i_input_data[868 % IN_WIDTH] : pong_storage_data_87 ^ i_input_data[868 % IN_WIDTH];
                default: pong_storage_data_87 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_87;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_87 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_87;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_87 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_87;
            end
        end
    end
end

logic ping_storage_data_88;
logic pong_storage_data_88;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_88 <= 1'b0;
        pong_storage_data_88 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                186 / IN_WIDTH: ping_storage_data_88 <= (fillup_transition == 1'b1) ? i_input_data[186 % IN_WIDTH] : ping_storage_data_88 ^ i_input_data[186 % IN_WIDTH];
                207 / IN_WIDTH: ping_storage_data_88 <= (fillup_transition == 1'b1) ? i_input_data[207 % IN_WIDTH] : ping_storage_data_88 ^ i_input_data[207 % IN_WIDTH];
                801 / IN_WIDTH: ping_storage_data_88 <= (fillup_transition == 1'b1) ? i_input_data[801 % IN_WIDTH] : ping_storage_data_88 ^ i_input_data[801 % IN_WIDTH];
                869 / IN_WIDTH: ping_storage_data_88 <= (fillup_transition == 1'b1) ? i_input_data[869 % IN_WIDTH] : ping_storage_data_88 ^ i_input_data[869 % IN_WIDTH];
                default: ping_storage_data_88 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_88;
                endcase
            end else begin
                case (input_count)
                186 / IN_WIDTH: pong_storage_data_88 <= (fillup_transition == 1'b1) ? i_input_data[186 % IN_WIDTH] : pong_storage_data_88 ^ i_input_data[186 % IN_WIDTH];
                207 / IN_WIDTH: pong_storage_data_88 <= (fillup_transition == 1'b1) ? i_input_data[207 % IN_WIDTH] : pong_storage_data_88 ^ i_input_data[207 % IN_WIDTH];
                801 / IN_WIDTH: pong_storage_data_88 <= (fillup_transition == 1'b1) ? i_input_data[801 % IN_WIDTH] : pong_storage_data_88 ^ i_input_data[801 % IN_WIDTH];
                869 / IN_WIDTH: pong_storage_data_88 <= (fillup_transition == 1'b1) ? i_input_data[869 % IN_WIDTH] : pong_storage_data_88 ^ i_input_data[869 % IN_WIDTH];
                default: pong_storage_data_88 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_88;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_88 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_88;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_88 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_88;
            end
        end
    end
end

logic ping_storage_data_89;
logic pong_storage_data_89;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_89 <= 1'b0;
        pong_storage_data_89 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                187 / IN_WIDTH: ping_storage_data_89 <= (fillup_transition == 1'b1) ? i_input_data[187 % IN_WIDTH] : ping_storage_data_89 ^ i_input_data[187 % IN_WIDTH];
                208 / IN_WIDTH: ping_storage_data_89 <= (fillup_transition == 1'b1) ? i_input_data[208 % IN_WIDTH] : ping_storage_data_89 ^ i_input_data[208 % IN_WIDTH];
                802 / IN_WIDTH: ping_storage_data_89 <= (fillup_transition == 1'b1) ? i_input_data[802 % IN_WIDTH] : ping_storage_data_89 ^ i_input_data[802 % IN_WIDTH];
                870 / IN_WIDTH: ping_storage_data_89 <= (fillup_transition == 1'b1) ? i_input_data[870 % IN_WIDTH] : ping_storage_data_89 ^ i_input_data[870 % IN_WIDTH];
                default: ping_storage_data_89 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_89;
                endcase
            end else begin
                case (input_count)
                187 / IN_WIDTH: pong_storage_data_89 <= (fillup_transition == 1'b1) ? i_input_data[187 % IN_WIDTH] : pong_storage_data_89 ^ i_input_data[187 % IN_WIDTH];
                208 / IN_WIDTH: pong_storage_data_89 <= (fillup_transition == 1'b1) ? i_input_data[208 % IN_WIDTH] : pong_storage_data_89 ^ i_input_data[208 % IN_WIDTH];
                802 / IN_WIDTH: pong_storage_data_89 <= (fillup_transition == 1'b1) ? i_input_data[802 % IN_WIDTH] : pong_storage_data_89 ^ i_input_data[802 % IN_WIDTH];
                870 / IN_WIDTH: pong_storage_data_89 <= (fillup_transition == 1'b1) ? i_input_data[870 % IN_WIDTH] : pong_storage_data_89 ^ i_input_data[870 % IN_WIDTH];
                default: pong_storage_data_89 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_89;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_89 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_89;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_89 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_89;
            end
        end
    end
end

logic ping_storage_data_90;
logic pong_storage_data_90;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_90 <= 1'b0;
        pong_storage_data_90 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                188 / IN_WIDTH: ping_storage_data_90 <= (fillup_transition == 1'b1) ? i_input_data[188 % IN_WIDTH] : ping_storage_data_90 ^ i_input_data[188 % IN_WIDTH];
                209 / IN_WIDTH: ping_storage_data_90 <= (fillup_transition == 1'b1) ? i_input_data[209 % IN_WIDTH] : ping_storage_data_90 ^ i_input_data[209 % IN_WIDTH];
                803 / IN_WIDTH: ping_storage_data_90 <= (fillup_transition == 1'b1) ? i_input_data[803 % IN_WIDTH] : ping_storage_data_90 ^ i_input_data[803 % IN_WIDTH];
                871 / IN_WIDTH: ping_storage_data_90 <= (fillup_transition == 1'b1) ? i_input_data[871 % IN_WIDTH] : ping_storage_data_90 ^ i_input_data[871 % IN_WIDTH];
                default: ping_storage_data_90 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_90;
                endcase
            end else begin
                case (input_count)
                188 / IN_WIDTH: pong_storage_data_90 <= (fillup_transition == 1'b1) ? i_input_data[188 % IN_WIDTH] : pong_storage_data_90 ^ i_input_data[188 % IN_WIDTH];
                209 / IN_WIDTH: pong_storage_data_90 <= (fillup_transition == 1'b1) ? i_input_data[209 % IN_WIDTH] : pong_storage_data_90 ^ i_input_data[209 % IN_WIDTH];
                803 / IN_WIDTH: pong_storage_data_90 <= (fillup_transition == 1'b1) ? i_input_data[803 % IN_WIDTH] : pong_storage_data_90 ^ i_input_data[803 % IN_WIDTH];
                871 / IN_WIDTH: pong_storage_data_90 <= (fillup_transition == 1'b1) ? i_input_data[871 % IN_WIDTH] : pong_storage_data_90 ^ i_input_data[871 % IN_WIDTH];
                default: pong_storage_data_90 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_90;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_90 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_90;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_90 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_90;
            end
        end
    end
end

logic ping_storage_data_91;
logic pong_storage_data_91;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_91 <= 1'b0;
        pong_storage_data_91 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                189 / IN_WIDTH: ping_storage_data_91 <= (fillup_transition == 1'b1) ? i_input_data[189 % IN_WIDTH] : ping_storage_data_91 ^ i_input_data[189 % IN_WIDTH];
                210 / IN_WIDTH: ping_storage_data_91 <= (fillup_transition == 1'b1) ? i_input_data[210 % IN_WIDTH] : ping_storage_data_91 ^ i_input_data[210 % IN_WIDTH];
                804 / IN_WIDTH: ping_storage_data_91 <= (fillup_transition == 1'b1) ? i_input_data[804 % IN_WIDTH] : ping_storage_data_91 ^ i_input_data[804 % IN_WIDTH];
                872 / IN_WIDTH: ping_storage_data_91 <= (fillup_transition == 1'b1) ? i_input_data[872 % IN_WIDTH] : ping_storage_data_91 ^ i_input_data[872 % IN_WIDTH];
                default: ping_storage_data_91 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_91;
                endcase
            end else begin
                case (input_count)
                189 / IN_WIDTH: pong_storage_data_91 <= (fillup_transition == 1'b1) ? i_input_data[189 % IN_WIDTH] : pong_storage_data_91 ^ i_input_data[189 % IN_WIDTH];
                210 / IN_WIDTH: pong_storage_data_91 <= (fillup_transition == 1'b1) ? i_input_data[210 % IN_WIDTH] : pong_storage_data_91 ^ i_input_data[210 % IN_WIDTH];
                804 / IN_WIDTH: pong_storage_data_91 <= (fillup_transition == 1'b1) ? i_input_data[804 % IN_WIDTH] : pong_storage_data_91 ^ i_input_data[804 % IN_WIDTH];
                872 / IN_WIDTH: pong_storage_data_91 <= (fillup_transition == 1'b1) ? i_input_data[872 % IN_WIDTH] : pong_storage_data_91 ^ i_input_data[872 % IN_WIDTH];
                default: pong_storage_data_91 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_91;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_91 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_91;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_91 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_91;
            end
        end
    end
end

logic ping_storage_data_92;
logic pong_storage_data_92;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_92 <= 1'b0;
        pong_storage_data_92 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                190 / IN_WIDTH: ping_storage_data_92 <= (fillup_transition == 1'b1) ? i_input_data[190 % IN_WIDTH] : ping_storage_data_92 ^ i_input_data[190 % IN_WIDTH];
                211 / IN_WIDTH: ping_storage_data_92 <= (fillup_transition == 1'b1) ? i_input_data[211 % IN_WIDTH] : ping_storage_data_92 ^ i_input_data[211 % IN_WIDTH];
                805 / IN_WIDTH: ping_storage_data_92 <= (fillup_transition == 1'b1) ? i_input_data[805 % IN_WIDTH] : ping_storage_data_92 ^ i_input_data[805 % IN_WIDTH];
                873 / IN_WIDTH: ping_storage_data_92 <= (fillup_transition == 1'b1) ? i_input_data[873 % IN_WIDTH] : ping_storage_data_92 ^ i_input_data[873 % IN_WIDTH];
                default: ping_storage_data_92 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_92;
                endcase
            end else begin
                case (input_count)
                190 / IN_WIDTH: pong_storage_data_92 <= (fillup_transition == 1'b1) ? i_input_data[190 % IN_WIDTH] : pong_storage_data_92 ^ i_input_data[190 % IN_WIDTH];
                211 / IN_WIDTH: pong_storage_data_92 <= (fillup_transition == 1'b1) ? i_input_data[211 % IN_WIDTH] : pong_storage_data_92 ^ i_input_data[211 % IN_WIDTH];
                805 / IN_WIDTH: pong_storage_data_92 <= (fillup_transition == 1'b1) ? i_input_data[805 % IN_WIDTH] : pong_storage_data_92 ^ i_input_data[805 % IN_WIDTH];
                873 / IN_WIDTH: pong_storage_data_92 <= (fillup_transition == 1'b1) ? i_input_data[873 % IN_WIDTH] : pong_storage_data_92 ^ i_input_data[873 % IN_WIDTH];
                default: pong_storage_data_92 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_92;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_92 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_92;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_92 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_92;
            end
        end
    end
end

logic ping_storage_data_93;
logic pong_storage_data_93;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_93 <= 1'b0;
        pong_storage_data_93 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                191 / IN_WIDTH: ping_storage_data_93 <= (fillup_transition == 1'b1) ? i_input_data[191 % IN_WIDTH] : ping_storage_data_93 ^ i_input_data[191 % IN_WIDTH];
                212 / IN_WIDTH: ping_storage_data_93 <= (fillup_transition == 1'b1) ? i_input_data[212 % IN_WIDTH] : ping_storage_data_93 ^ i_input_data[212 % IN_WIDTH];
                806 / IN_WIDTH: ping_storage_data_93 <= (fillup_transition == 1'b1) ? i_input_data[806 % IN_WIDTH] : ping_storage_data_93 ^ i_input_data[806 % IN_WIDTH];
                874 / IN_WIDTH: ping_storage_data_93 <= (fillup_transition == 1'b1) ? i_input_data[874 % IN_WIDTH] : ping_storage_data_93 ^ i_input_data[874 % IN_WIDTH];
                default: ping_storage_data_93 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_93;
                endcase
            end else begin
                case (input_count)
                191 / IN_WIDTH: pong_storage_data_93 <= (fillup_transition == 1'b1) ? i_input_data[191 % IN_WIDTH] : pong_storage_data_93 ^ i_input_data[191 % IN_WIDTH];
                212 / IN_WIDTH: pong_storage_data_93 <= (fillup_transition == 1'b1) ? i_input_data[212 % IN_WIDTH] : pong_storage_data_93 ^ i_input_data[212 % IN_WIDTH];
                806 / IN_WIDTH: pong_storage_data_93 <= (fillup_transition == 1'b1) ? i_input_data[806 % IN_WIDTH] : pong_storage_data_93 ^ i_input_data[806 % IN_WIDTH];
                874 / IN_WIDTH: pong_storage_data_93 <= (fillup_transition == 1'b1) ? i_input_data[874 % IN_WIDTH] : pong_storage_data_93 ^ i_input_data[874 % IN_WIDTH];
                default: pong_storage_data_93 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_93;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_93 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_93;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_93 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_93;
            end
        end
    end
end

logic ping_storage_data_94;
logic pong_storage_data_94;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_94 <= 1'b0;
        pong_storage_data_94 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                96 / IN_WIDTH: ping_storage_data_94 <= (fillup_transition == 1'b1) ? i_input_data[96 % IN_WIDTH] : ping_storage_data_94 ^ i_input_data[96 % IN_WIDTH];
                213 / IN_WIDTH: ping_storage_data_94 <= (fillup_transition == 1'b1) ? i_input_data[213 % IN_WIDTH] : ping_storage_data_94 ^ i_input_data[213 % IN_WIDTH];
                807 / IN_WIDTH: ping_storage_data_94 <= (fillup_transition == 1'b1) ? i_input_data[807 % IN_WIDTH] : ping_storage_data_94 ^ i_input_data[807 % IN_WIDTH];
                875 / IN_WIDTH: ping_storage_data_94 <= (fillup_transition == 1'b1) ? i_input_data[875 % IN_WIDTH] : ping_storage_data_94 ^ i_input_data[875 % IN_WIDTH];
                default: ping_storage_data_94 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_94;
                endcase
            end else begin
                case (input_count)
                96 / IN_WIDTH: pong_storage_data_94 <= (fillup_transition == 1'b1) ? i_input_data[96 % IN_WIDTH] : pong_storage_data_94 ^ i_input_data[96 % IN_WIDTH];
                213 / IN_WIDTH: pong_storage_data_94 <= (fillup_transition == 1'b1) ? i_input_data[213 % IN_WIDTH] : pong_storage_data_94 ^ i_input_data[213 % IN_WIDTH];
                807 / IN_WIDTH: pong_storage_data_94 <= (fillup_transition == 1'b1) ? i_input_data[807 % IN_WIDTH] : pong_storage_data_94 ^ i_input_data[807 % IN_WIDTH];
                875 / IN_WIDTH: pong_storage_data_94 <= (fillup_transition == 1'b1) ? i_input_data[875 % IN_WIDTH] : pong_storage_data_94 ^ i_input_data[875 % IN_WIDTH];
                default: pong_storage_data_94 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_94;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_94 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_94;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_94 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_94;
            end
        end
    end
end

logic ping_storage_data_95;
logic pong_storage_data_95;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_95 <= 1'b0;
        pong_storage_data_95 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                97 / IN_WIDTH: ping_storage_data_95 <= (fillup_transition == 1'b1) ? i_input_data[97 % IN_WIDTH] : ping_storage_data_95 ^ i_input_data[97 % IN_WIDTH];
                214 / IN_WIDTH: ping_storage_data_95 <= (fillup_transition == 1'b1) ? i_input_data[214 % IN_WIDTH] : ping_storage_data_95 ^ i_input_data[214 % IN_WIDTH];
                808 / IN_WIDTH: ping_storage_data_95 <= (fillup_transition == 1'b1) ? i_input_data[808 % IN_WIDTH] : ping_storage_data_95 ^ i_input_data[808 % IN_WIDTH];
                876 / IN_WIDTH: ping_storage_data_95 <= (fillup_transition == 1'b1) ? i_input_data[876 % IN_WIDTH] : ping_storage_data_95 ^ i_input_data[876 % IN_WIDTH];
                default: ping_storage_data_95 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_95;
                endcase
            end else begin
                case (input_count)
                97 / IN_WIDTH: pong_storage_data_95 <= (fillup_transition == 1'b1) ? i_input_data[97 % IN_WIDTH] : pong_storage_data_95 ^ i_input_data[97 % IN_WIDTH];
                214 / IN_WIDTH: pong_storage_data_95 <= (fillup_transition == 1'b1) ? i_input_data[214 % IN_WIDTH] : pong_storage_data_95 ^ i_input_data[214 % IN_WIDTH];
                808 / IN_WIDTH: pong_storage_data_95 <= (fillup_transition == 1'b1) ? i_input_data[808 % IN_WIDTH] : pong_storage_data_95 ^ i_input_data[808 % IN_WIDTH];
                876 / IN_WIDTH: pong_storage_data_95 <= (fillup_transition == 1'b1) ? i_input_data[876 % IN_WIDTH] : pong_storage_data_95 ^ i_input_data[876 % IN_WIDTH];
                default: pong_storage_data_95 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_95;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_95 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_95;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_95 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_95;
            end
        end
    end
end

logic ping_storage_data_96;
logic pong_storage_data_96;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_96 <= 1'b0;
        pong_storage_data_96 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                165 / IN_WIDTH: ping_storage_data_96 <= (fillup_transition == 1'b1) ? i_input_data[165 % IN_WIDTH] : ping_storage_data_96 ^ i_input_data[165 % IN_WIDTH];
                554 / IN_WIDTH: ping_storage_data_96 <= (fillup_transition == 1'b1) ? i_input_data[554 % IN_WIDTH] : ping_storage_data_96 ^ i_input_data[554 % IN_WIDTH];
                593 / IN_WIDTH: ping_storage_data_96 <= (fillup_transition == 1'b1) ? i_input_data[593 % IN_WIDTH] : ping_storage_data_96 ^ i_input_data[593 % IN_WIDTH];
                759 / IN_WIDTH: ping_storage_data_96 <= (fillup_transition == 1'b1) ? i_input_data[759 % IN_WIDTH] : ping_storage_data_96 ^ i_input_data[759 % IN_WIDTH];
                1140 / IN_WIDTH: ping_storage_data_96 <= (fillup_transition == 1'b1) ? i_input_data[1140 % IN_WIDTH] : ping_storage_data_96 ^ i_input_data[1140 % IN_WIDTH];
                default: ping_storage_data_96 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_96;
                endcase
            end else begin
                case (input_count)
                165 / IN_WIDTH: pong_storage_data_96 <= (fillup_transition == 1'b1) ? i_input_data[165 % IN_WIDTH] : pong_storage_data_96 ^ i_input_data[165 % IN_WIDTH];
                554 / IN_WIDTH: pong_storage_data_96 <= (fillup_transition == 1'b1) ? i_input_data[554 % IN_WIDTH] : pong_storage_data_96 ^ i_input_data[554 % IN_WIDTH];
                593 / IN_WIDTH: pong_storage_data_96 <= (fillup_transition == 1'b1) ? i_input_data[593 % IN_WIDTH] : pong_storage_data_96 ^ i_input_data[593 % IN_WIDTH];
                759 / IN_WIDTH: pong_storage_data_96 <= (fillup_transition == 1'b1) ? i_input_data[759 % IN_WIDTH] : pong_storage_data_96 ^ i_input_data[759 % IN_WIDTH];
                1140 / IN_WIDTH: pong_storage_data_96 <= (fillup_transition == 1'b1) ? i_input_data[1140 % IN_WIDTH] : pong_storage_data_96 ^ i_input_data[1140 % IN_WIDTH];
                default: pong_storage_data_96 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_96;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_96 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_96;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_96 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_96;
            end
        end
    end
end

logic ping_storage_data_97;
logic pong_storage_data_97;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_97 <= 1'b0;
        pong_storage_data_97 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                166 / IN_WIDTH: ping_storage_data_97 <= (fillup_transition == 1'b1) ? i_input_data[166 % IN_WIDTH] : ping_storage_data_97 ^ i_input_data[166 % IN_WIDTH];
                555 / IN_WIDTH: ping_storage_data_97 <= (fillup_transition == 1'b1) ? i_input_data[555 % IN_WIDTH] : ping_storage_data_97 ^ i_input_data[555 % IN_WIDTH];
                594 / IN_WIDTH: ping_storage_data_97 <= (fillup_transition == 1'b1) ? i_input_data[594 % IN_WIDTH] : ping_storage_data_97 ^ i_input_data[594 % IN_WIDTH];
                760 / IN_WIDTH: ping_storage_data_97 <= (fillup_transition == 1'b1) ? i_input_data[760 % IN_WIDTH] : ping_storage_data_97 ^ i_input_data[760 % IN_WIDTH];
                1141 / IN_WIDTH: ping_storage_data_97 <= (fillup_transition == 1'b1) ? i_input_data[1141 % IN_WIDTH] : ping_storage_data_97 ^ i_input_data[1141 % IN_WIDTH];
                default: ping_storage_data_97 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_97;
                endcase
            end else begin
                case (input_count)
                166 / IN_WIDTH: pong_storage_data_97 <= (fillup_transition == 1'b1) ? i_input_data[166 % IN_WIDTH] : pong_storage_data_97 ^ i_input_data[166 % IN_WIDTH];
                555 / IN_WIDTH: pong_storage_data_97 <= (fillup_transition == 1'b1) ? i_input_data[555 % IN_WIDTH] : pong_storage_data_97 ^ i_input_data[555 % IN_WIDTH];
                594 / IN_WIDTH: pong_storage_data_97 <= (fillup_transition == 1'b1) ? i_input_data[594 % IN_WIDTH] : pong_storage_data_97 ^ i_input_data[594 % IN_WIDTH];
                760 / IN_WIDTH: pong_storage_data_97 <= (fillup_transition == 1'b1) ? i_input_data[760 % IN_WIDTH] : pong_storage_data_97 ^ i_input_data[760 % IN_WIDTH];
                1141 / IN_WIDTH: pong_storage_data_97 <= (fillup_transition == 1'b1) ? i_input_data[1141 % IN_WIDTH] : pong_storage_data_97 ^ i_input_data[1141 % IN_WIDTH];
                default: pong_storage_data_97 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_97;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_97 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_97;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_97 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_97;
            end
        end
    end
end

logic ping_storage_data_98;
logic pong_storage_data_98;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_98 <= 1'b0;
        pong_storage_data_98 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                167 / IN_WIDTH: ping_storage_data_98 <= (fillup_transition == 1'b1) ? i_input_data[167 % IN_WIDTH] : ping_storage_data_98 ^ i_input_data[167 % IN_WIDTH];
                556 / IN_WIDTH: ping_storage_data_98 <= (fillup_transition == 1'b1) ? i_input_data[556 % IN_WIDTH] : ping_storage_data_98 ^ i_input_data[556 % IN_WIDTH];
                595 / IN_WIDTH: ping_storage_data_98 <= (fillup_transition == 1'b1) ? i_input_data[595 % IN_WIDTH] : ping_storage_data_98 ^ i_input_data[595 % IN_WIDTH];
                761 / IN_WIDTH: ping_storage_data_98 <= (fillup_transition == 1'b1) ? i_input_data[761 % IN_WIDTH] : ping_storage_data_98 ^ i_input_data[761 % IN_WIDTH];
                1142 / IN_WIDTH: ping_storage_data_98 <= (fillup_transition == 1'b1) ? i_input_data[1142 % IN_WIDTH] : ping_storage_data_98 ^ i_input_data[1142 % IN_WIDTH];
                default: ping_storage_data_98 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_98;
                endcase
            end else begin
                case (input_count)
                167 / IN_WIDTH: pong_storage_data_98 <= (fillup_transition == 1'b1) ? i_input_data[167 % IN_WIDTH] : pong_storage_data_98 ^ i_input_data[167 % IN_WIDTH];
                556 / IN_WIDTH: pong_storage_data_98 <= (fillup_transition == 1'b1) ? i_input_data[556 % IN_WIDTH] : pong_storage_data_98 ^ i_input_data[556 % IN_WIDTH];
                595 / IN_WIDTH: pong_storage_data_98 <= (fillup_transition == 1'b1) ? i_input_data[595 % IN_WIDTH] : pong_storage_data_98 ^ i_input_data[595 % IN_WIDTH];
                761 / IN_WIDTH: pong_storage_data_98 <= (fillup_transition == 1'b1) ? i_input_data[761 % IN_WIDTH] : pong_storage_data_98 ^ i_input_data[761 % IN_WIDTH];
                1142 / IN_WIDTH: pong_storage_data_98 <= (fillup_transition == 1'b1) ? i_input_data[1142 % IN_WIDTH] : pong_storage_data_98 ^ i_input_data[1142 % IN_WIDTH];
                default: pong_storage_data_98 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_98;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_98 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_98;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_98 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_98;
            end
        end
    end
end

logic ping_storage_data_99;
logic pong_storage_data_99;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_99 <= 1'b0;
        pong_storage_data_99 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                168 / IN_WIDTH: ping_storage_data_99 <= (fillup_transition == 1'b1) ? i_input_data[168 % IN_WIDTH] : ping_storage_data_99 ^ i_input_data[168 % IN_WIDTH];
                557 / IN_WIDTH: ping_storage_data_99 <= (fillup_transition == 1'b1) ? i_input_data[557 % IN_WIDTH] : ping_storage_data_99 ^ i_input_data[557 % IN_WIDTH];
                596 / IN_WIDTH: ping_storage_data_99 <= (fillup_transition == 1'b1) ? i_input_data[596 % IN_WIDTH] : ping_storage_data_99 ^ i_input_data[596 % IN_WIDTH];
                762 / IN_WIDTH: ping_storage_data_99 <= (fillup_transition == 1'b1) ? i_input_data[762 % IN_WIDTH] : ping_storage_data_99 ^ i_input_data[762 % IN_WIDTH];
                1143 / IN_WIDTH: ping_storage_data_99 <= (fillup_transition == 1'b1) ? i_input_data[1143 % IN_WIDTH] : ping_storage_data_99 ^ i_input_data[1143 % IN_WIDTH];
                default: ping_storage_data_99 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_99;
                endcase
            end else begin
                case (input_count)
                168 / IN_WIDTH: pong_storage_data_99 <= (fillup_transition == 1'b1) ? i_input_data[168 % IN_WIDTH] : pong_storage_data_99 ^ i_input_data[168 % IN_WIDTH];
                557 / IN_WIDTH: pong_storage_data_99 <= (fillup_transition == 1'b1) ? i_input_data[557 % IN_WIDTH] : pong_storage_data_99 ^ i_input_data[557 % IN_WIDTH];
                596 / IN_WIDTH: pong_storage_data_99 <= (fillup_transition == 1'b1) ? i_input_data[596 % IN_WIDTH] : pong_storage_data_99 ^ i_input_data[596 % IN_WIDTH];
                762 / IN_WIDTH: pong_storage_data_99 <= (fillup_transition == 1'b1) ? i_input_data[762 % IN_WIDTH] : pong_storage_data_99 ^ i_input_data[762 % IN_WIDTH];
                1143 / IN_WIDTH: pong_storage_data_99 <= (fillup_transition == 1'b1) ? i_input_data[1143 % IN_WIDTH] : pong_storage_data_99 ^ i_input_data[1143 % IN_WIDTH];
                default: pong_storage_data_99 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_99;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_99 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_99;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_99 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_99;
            end
        end
    end
end

logic ping_storage_data_100;
logic pong_storage_data_100;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_100 <= 1'b0;
        pong_storage_data_100 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                169 / IN_WIDTH: ping_storage_data_100 <= (fillup_transition == 1'b1) ? i_input_data[169 % IN_WIDTH] : ping_storage_data_100 ^ i_input_data[169 % IN_WIDTH];
                558 / IN_WIDTH: ping_storage_data_100 <= (fillup_transition == 1'b1) ? i_input_data[558 % IN_WIDTH] : ping_storage_data_100 ^ i_input_data[558 % IN_WIDTH];
                597 / IN_WIDTH: ping_storage_data_100 <= (fillup_transition == 1'b1) ? i_input_data[597 % IN_WIDTH] : ping_storage_data_100 ^ i_input_data[597 % IN_WIDTH];
                763 / IN_WIDTH: ping_storage_data_100 <= (fillup_transition == 1'b1) ? i_input_data[763 % IN_WIDTH] : ping_storage_data_100 ^ i_input_data[763 % IN_WIDTH];
                1144 / IN_WIDTH: ping_storage_data_100 <= (fillup_transition == 1'b1) ? i_input_data[1144 % IN_WIDTH] : ping_storage_data_100 ^ i_input_data[1144 % IN_WIDTH];
                default: ping_storage_data_100 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_100;
                endcase
            end else begin
                case (input_count)
                169 / IN_WIDTH: pong_storage_data_100 <= (fillup_transition == 1'b1) ? i_input_data[169 % IN_WIDTH] : pong_storage_data_100 ^ i_input_data[169 % IN_WIDTH];
                558 / IN_WIDTH: pong_storage_data_100 <= (fillup_transition == 1'b1) ? i_input_data[558 % IN_WIDTH] : pong_storage_data_100 ^ i_input_data[558 % IN_WIDTH];
                597 / IN_WIDTH: pong_storage_data_100 <= (fillup_transition == 1'b1) ? i_input_data[597 % IN_WIDTH] : pong_storage_data_100 ^ i_input_data[597 % IN_WIDTH];
                763 / IN_WIDTH: pong_storage_data_100 <= (fillup_transition == 1'b1) ? i_input_data[763 % IN_WIDTH] : pong_storage_data_100 ^ i_input_data[763 % IN_WIDTH];
                1144 / IN_WIDTH: pong_storage_data_100 <= (fillup_transition == 1'b1) ? i_input_data[1144 % IN_WIDTH] : pong_storage_data_100 ^ i_input_data[1144 % IN_WIDTH];
                default: pong_storage_data_100 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_100;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_100 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_100;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_100 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_100;
            end
        end
    end
end

logic ping_storage_data_101;
logic pong_storage_data_101;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_101 <= 1'b0;
        pong_storage_data_101 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                170 / IN_WIDTH: ping_storage_data_101 <= (fillup_transition == 1'b1) ? i_input_data[170 % IN_WIDTH] : ping_storage_data_101 ^ i_input_data[170 % IN_WIDTH];
                559 / IN_WIDTH: ping_storage_data_101 <= (fillup_transition == 1'b1) ? i_input_data[559 % IN_WIDTH] : ping_storage_data_101 ^ i_input_data[559 % IN_WIDTH];
                598 / IN_WIDTH: ping_storage_data_101 <= (fillup_transition == 1'b1) ? i_input_data[598 % IN_WIDTH] : ping_storage_data_101 ^ i_input_data[598 % IN_WIDTH];
                764 / IN_WIDTH: ping_storage_data_101 <= (fillup_transition == 1'b1) ? i_input_data[764 % IN_WIDTH] : ping_storage_data_101 ^ i_input_data[764 % IN_WIDTH];
                1145 / IN_WIDTH: ping_storage_data_101 <= (fillup_transition == 1'b1) ? i_input_data[1145 % IN_WIDTH] : ping_storage_data_101 ^ i_input_data[1145 % IN_WIDTH];
                default: ping_storage_data_101 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_101;
                endcase
            end else begin
                case (input_count)
                170 / IN_WIDTH: pong_storage_data_101 <= (fillup_transition == 1'b1) ? i_input_data[170 % IN_WIDTH] : pong_storage_data_101 ^ i_input_data[170 % IN_WIDTH];
                559 / IN_WIDTH: pong_storage_data_101 <= (fillup_transition == 1'b1) ? i_input_data[559 % IN_WIDTH] : pong_storage_data_101 ^ i_input_data[559 % IN_WIDTH];
                598 / IN_WIDTH: pong_storage_data_101 <= (fillup_transition == 1'b1) ? i_input_data[598 % IN_WIDTH] : pong_storage_data_101 ^ i_input_data[598 % IN_WIDTH];
                764 / IN_WIDTH: pong_storage_data_101 <= (fillup_transition == 1'b1) ? i_input_data[764 % IN_WIDTH] : pong_storage_data_101 ^ i_input_data[764 % IN_WIDTH];
                1145 / IN_WIDTH: pong_storage_data_101 <= (fillup_transition == 1'b1) ? i_input_data[1145 % IN_WIDTH] : pong_storage_data_101 ^ i_input_data[1145 % IN_WIDTH];
                default: pong_storage_data_101 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_101;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_101 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_101;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_101 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_101;
            end
        end
    end
end

logic ping_storage_data_102;
logic pong_storage_data_102;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_102 <= 1'b0;
        pong_storage_data_102 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                171 / IN_WIDTH: ping_storage_data_102 <= (fillup_transition == 1'b1) ? i_input_data[171 % IN_WIDTH] : ping_storage_data_102 ^ i_input_data[171 % IN_WIDTH];
                560 / IN_WIDTH: ping_storage_data_102 <= (fillup_transition == 1'b1) ? i_input_data[560 % IN_WIDTH] : ping_storage_data_102 ^ i_input_data[560 % IN_WIDTH];
                599 / IN_WIDTH: ping_storage_data_102 <= (fillup_transition == 1'b1) ? i_input_data[599 % IN_WIDTH] : ping_storage_data_102 ^ i_input_data[599 % IN_WIDTH];
                765 / IN_WIDTH: ping_storage_data_102 <= (fillup_transition == 1'b1) ? i_input_data[765 % IN_WIDTH] : ping_storage_data_102 ^ i_input_data[765 % IN_WIDTH];
                1146 / IN_WIDTH: ping_storage_data_102 <= (fillup_transition == 1'b1) ? i_input_data[1146 % IN_WIDTH] : ping_storage_data_102 ^ i_input_data[1146 % IN_WIDTH];
                default: ping_storage_data_102 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_102;
                endcase
            end else begin
                case (input_count)
                171 / IN_WIDTH: pong_storage_data_102 <= (fillup_transition == 1'b1) ? i_input_data[171 % IN_WIDTH] : pong_storage_data_102 ^ i_input_data[171 % IN_WIDTH];
                560 / IN_WIDTH: pong_storage_data_102 <= (fillup_transition == 1'b1) ? i_input_data[560 % IN_WIDTH] : pong_storage_data_102 ^ i_input_data[560 % IN_WIDTH];
                599 / IN_WIDTH: pong_storage_data_102 <= (fillup_transition == 1'b1) ? i_input_data[599 % IN_WIDTH] : pong_storage_data_102 ^ i_input_data[599 % IN_WIDTH];
                765 / IN_WIDTH: pong_storage_data_102 <= (fillup_transition == 1'b1) ? i_input_data[765 % IN_WIDTH] : pong_storage_data_102 ^ i_input_data[765 % IN_WIDTH];
                1146 / IN_WIDTH: pong_storage_data_102 <= (fillup_transition == 1'b1) ? i_input_data[1146 % IN_WIDTH] : pong_storage_data_102 ^ i_input_data[1146 % IN_WIDTH];
                default: pong_storage_data_102 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_102;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_102 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_102;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_102 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_102;
            end
        end
    end
end

logic ping_storage_data_103;
logic pong_storage_data_103;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_103 <= 1'b0;
        pong_storage_data_103 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                172 / IN_WIDTH: ping_storage_data_103 <= (fillup_transition == 1'b1) ? i_input_data[172 % IN_WIDTH] : ping_storage_data_103 ^ i_input_data[172 % IN_WIDTH];
                561 / IN_WIDTH: ping_storage_data_103 <= (fillup_transition == 1'b1) ? i_input_data[561 % IN_WIDTH] : ping_storage_data_103 ^ i_input_data[561 % IN_WIDTH];
                600 / IN_WIDTH: ping_storage_data_103 <= (fillup_transition == 1'b1) ? i_input_data[600 % IN_WIDTH] : ping_storage_data_103 ^ i_input_data[600 % IN_WIDTH];
                766 / IN_WIDTH: ping_storage_data_103 <= (fillup_transition == 1'b1) ? i_input_data[766 % IN_WIDTH] : ping_storage_data_103 ^ i_input_data[766 % IN_WIDTH];
                1147 / IN_WIDTH: ping_storage_data_103 <= (fillup_transition == 1'b1) ? i_input_data[1147 % IN_WIDTH] : ping_storage_data_103 ^ i_input_data[1147 % IN_WIDTH];
                default: ping_storage_data_103 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_103;
                endcase
            end else begin
                case (input_count)
                172 / IN_WIDTH: pong_storage_data_103 <= (fillup_transition == 1'b1) ? i_input_data[172 % IN_WIDTH] : pong_storage_data_103 ^ i_input_data[172 % IN_WIDTH];
                561 / IN_WIDTH: pong_storage_data_103 <= (fillup_transition == 1'b1) ? i_input_data[561 % IN_WIDTH] : pong_storage_data_103 ^ i_input_data[561 % IN_WIDTH];
                600 / IN_WIDTH: pong_storage_data_103 <= (fillup_transition == 1'b1) ? i_input_data[600 % IN_WIDTH] : pong_storage_data_103 ^ i_input_data[600 % IN_WIDTH];
                766 / IN_WIDTH: pong_storage_data_103 <= (fillup_transition == 1'b1) ? i_input_data[766 % IN_WIDTH] : pong_storage_data_103 ^ i_input_data[766 % IN_WIDTH];
                1147 / IN_WIDTH: pong_storage_data_103 <= (fillup_transition == 1'b1) ? i_input_data[1147 % IN_WIDTH] : pong_storage_data_103 ^ i_input_data[1147 % IN_WIDTH];
                default: pong_storage_data_103 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_103;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_103 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_103;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_103 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_103;
            end
        end
    end
end

logic ping_storage_data_104;
logic pong_storage_data_104;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_104 <= 1'b0;
        pong_storage_data_104 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                173 / IN_WIDTH: ping_storage_data_104 <= (fillup_transition == 1'b1) ? i_input_data[173 % IN_WIDTH] : ping_storage_data_104 ^ i_input_data[173 % IN_WIDTH];
                562 / IN_WIDTH: ping_storage_data_104 <= (fillup_transition == 1'b1) ? i_input_data[562 % IN_WIDTH] : ping_storage_data_104 ^ i_input_data[562 % IN_WIDTH];
                601 / IN_WIDTH: ping_storage_data_104 <= (fillup_transition == 1'b1) ? i_input_data[601 % IN_WIDTH] : ping_storage_data_104 ^ i_input_data[601 % IN_WIDTH];
                767 / IN_WIDTH: ping_storage_data_104 <= (fillup_transition == 1'b1) ? i_input_data[767 % IN_WIDTH] : ping_storage_data_104 ^ i_input_data[767 % IN_WIDTH];
                1148 / IN_WIDTH: ping_storage_data_104 <= (fillup_transition == 1'b1) ? i_input_data[1148 % IN_WIDTH] : ping_storage_data_104 ^ i_input_data[1148 % IN_WIDTH];
                default: ping_storage_data_104 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_104;
                endcase
            end else begin
                case (input_count)
                173 / IN_WIDTH: pong_storage_data_104 <= (fillup_transition == 1'b1) ? i_input_data[173 % IN_WIDTH] : pong_storage_data_104 ^ i_input_data[173 % IN_WIDTH];
                562 / IN_WIDTH: pong_storage_data_104 <= (fillup_transition == 1'b1) ? i_input_data[562 % IN_WIDTH] : pong_storage_data_104 ^ i_input_data[562 % IN_WIDTH];
                601 / IN_WIDTH: pong_storage_data_104 <= (fillup_transition == 1'b1) ? i_input_data[601 % IN_WIDTH] : pong_storage_data_104 ^ i_input_data[601 % IN_WIDTH];
                767 / IN_WIDTH: pong_storage_data_104 <= (fillup_transition == 1'b1) ? i_input_data[767 % IN_WIDTH] : pong_storage_data_104 ^ i_input_data[767 % IN_WIDTH];
                1148 / IN_WIDTH: pong_storage_data_104 <= (fillup_transition == 1'b1) ? i_input_data[1148 % IN_WIDTH] : pong_storage_data_104 ^ i_input_data[1148 % IN_WIDTH];
                default: pong_storage_data_104 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_104;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_104 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_104;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_104 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_104;
            end
        end
    end
end

logic ping_storage_data_105;
logic pong_storage_data_105;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_105 <= 1'b0;
        pong_storage_data_105 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                174 / IN_WIDTH: ping_storage_data_105 <= (fillup_transition == 1'b1) ? i_input_data[174 % IN_WIDTH] : ping_storage_data_105 ^ i_input_data[174 % IN_WIDTH];
                563 / IN_WIDTH: ping_storage_data_105 <= (fillup_transition == 1'b1) ? i_input_data[563 % IN_WIDTH] : ping_storage_data_105 ^ i_input_data[563 % IN_WIDTH];
                602 / IN_WIDTH: ping_storage_data_105 <= (fillup_transition == 1'b1) ? i_input_data[602 % IN_WIDTH] : ping_storage_data_105 ^ i_input_data[602 % IN_WIDTH];
                672 / IN_WIDTH: ping_storage_data_105 <= (fillup_transition == 1'b1) ? i_input_data[672 % IN_WIDTH] : ping_storage_data_105 ^ i_input_data[672 % IN_WIDTH];
                1149 / IN_WIDTH: ping_storage_data_105 <= (fillup_transition == 1'b1) ? i_input_data[1149 % IN_WIDTH] : ping_storage_data_105 ^ i_input_data[1149 % IN_WIDTH];
                default: ping_storage_data_105 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_105;
                endcase
            end else begin
                case (input_count)
                174 / IN_WIDTH: pong_storage_data_105 <= (fillup_transition == 1'b1) ? i_input_data[174 % IN_WIDTH] : pong_storage_data_105 ^ i_input_data[174 % IN_WIDTH];
                563 / IN_WIDTH: pong_storage_data_105 <= (fillup_transition == 1'b1) ? i_input_data[563 % IN_WIDTH] : pong_storage_data_105 ^ i_input_data[563 % IN_WIDTH];
                602 / IN_WIDTH: pong_storage_data_105 <= (fillup_transition == 1'b1) ? i_input_data[602 % IN_WIDTH] : pong_storage_data_105 ^ i_input_data[602 % IN_WIDTH];
                672 / IN_WIDTH: pong_storage_data_105 <= (fillup_transition == 1'b1) ? i_input_data[672 % IN_WIDTH] : pong_storage_data_105 ^ i_input_data[672 % IN_WIDTH];
                1149 / IN_WIDTH: pong_storage_data_105 <= (fillup_transition == 1'b1) ? i_input_data[1149 % IN_WIDTH] : pong_storage_data_105 ^ i_input_data[1149 % IN_WIDTH];
                default: pong_storage_data_105 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_105;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_105 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_105;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_105 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_105;
            end
        end
    end
end

logic ping_storage_data_106;
logic pong_storage_data_106;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_106 <= 1'b0;
        pong_storage_data_106 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                175 / IN_WIDTH: ping_storage_data_106 <= (fillup_transition == 1'b1) ? i_input_data[175 % IN_WIDTH] : ping_storage_data_106 ^ i_input_data[175 % IN_WIDTH];
                564 / IN_WIDTH: ping_storage_data_106 <= (fillup_transition == 1'b1) ? i_input_data[564 % IN_WIDTH] : ping_storage_data_106 ^ i_input_data[564 % IN_WIDTH];
                603 / IN_WIDTH: ping_storage_data_106 <= (fillup_transition == 1'b1) ? i_input_data[603 % IN_WIDTH] : ping_storage_data_106 ^ i_input_data[603 % IN_WIDTH];
                673 / IN_WIDTH: ping_storage_data_106 <= (fillup_transition == 1'b1) ? i_input_data[673 % IN_WIDTH] : ping_storage_data_106 ^ i_input_data[673 % IN_WIDTH];
                1150 / IN_WIDTH: ping_storage_data_106 <= (fillup_transition == 1'b1) ? i_input_data[1150 % IN_WIDTH] : ping_storage_data_106 ^ i_input_data[1150 % IN_WIDTH];
                default: ping_storage_data_106 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_106;
                endcase
            end else begin
                case (input_count)
                175 / IN_WIDTH: pong_storage_data_106 <= (fillup_transition == 1'b1) ? i_input_data[175 % IN_WIDTH] : pong_storage_data_106 ^ i_input_data[175 % IN_WIDTH];
                564 / IN_WIDTH: pong_storage_data_106 <= (fillup_transition == 1'b1) ? i_input_data[564 % IN_WIDTH] : pong_storage_data_106 ^ i_input_data[564 % IN_WIDTH];
                603 / IN_WIDTH: pong_storage_data_106 <= (fillup_transition == 1'b1) ? i_input_data[603 % IN_WIDTH] : pong_storage_data_106 ^ i_input_data[603 % IN_WIDTH];
                673 / IN_WIDTH: pong_storage_data_106 <= (fillup_transition == 1'b1) ? i_input_data[673 % IN_WIDTH] : pong_storage_data_106 ^ i_input_data[673 % IN_WIDTH];
                1150 / IN_WIDTH: pong_storage_data_106 <= (fillup_transition == 1'b1) ? i_input_data[1150 % IN_WIDTH] : pong_storage_data_106 ^ i_input_data[1150 % IN_WIDTH];
                default: pong_storage_data_106 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_106;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_106 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_106;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_106 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_106;
            end
        end
    end
end

logic ping_storage_data_107;
logic pong_storage_data_107;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_107 <= 1'b0;
        pong_storage_data_107 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                176 / IN_WIDTH: ping_storage_data_107 <= (fillup_transition == 1'b1) ? i_input_data[176 % IN_WIDTH] : ping_storage_data_107 ^ i_input_data[176 % IN_WIDTH];
                565 / IN_WIDTH: ping_storage_data_107 <= (fillup_transition == 1'b1) ? i_input_data[565 % IN_WIDTH] : ping_storage_data_107 ^ i_input_data[565 % IN_WIDTH];
                604 / IN_WIDTH: ping_storage_data_107 <= (fillup_transition == 1'b1) ? i_input_data[604 % IN_WIDTH] : ping_storage_data_107 ^ i_input_data[604 % IN_WIDTH];
                674 / IN_WIDTH: ping_storage_data_107 <= (fillup_transition == 1'b1) ? i_input_data[674 % IN_WIDTH] : ping_storage_data_107 ^ i_input_data[674 % IN_WIDTH];
                1151 / IN_WIDTH: ping_storage_data_107 <= (fillup_transition == 1'b1) ? i_input_data[1151 % IN_WIDTH] : ping_storage_data_107 ^ i_input_data[1151 % IN_WIDTH];
                default: ping_storage_data_107 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_107;
                endcase
            end else begin
                case (input_count)
                176 / IN_WIDTH: pong_storage_data_107 <= (fillup_transition == 1'b1) ? i_input_data[176 % IN_WIDTH] : pong_storage_data_107 ^ i_input_data[176 % IN_WIDTH];
                565 / IN_WIDTH: pong_storage_data_107 <= (fillup_transition == 1'b1) ? i_input_data[565 % IN_WIDTH] : pong_storage_data_107 ^ i_input_data[565 % IN_WIDTH];
                604 / IN_WIDTH: pong_storage_data_107 <= (fillup_transition == 1'b1) ? i_input_data[604 % IN_WIDTH] : pong_storage_data_107 ^ i_input_data[604 % IN_WIDTH];
                674 / IN_WIDTH: pong_storage_data_107 <= (fillup_transition == 1'b1) ? i_input_data[674 % IN_WIDTH] : pong_storage_data_107 ^ i_input_data[674 % IN_WIDTH];
                1151 / IN_WIDTH: pong_storage_data_107 <= (fillup_transition == 1'b1) ? i_input_data[1151 % IN_WIDTH] : pong_storage_data_107 ^ i_input_data[1151 % IN_WIDTH];
                default: pong_storage_data_107 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_107;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_107 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_107;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_107 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_107;
            end
        end
    end
end

logic ping_storage_data_108;
logic pong_storage_data_108;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_108 <= 1'b0;
        pong_storage_data_108 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                177 / IN_WIDTH: ping_storage_data_108 <= (fillup_transition == 1'b1) ? i_input_data[177 % IN_WIDTH] : ping_storage_data_108 ^ i_input_data[177 % IN_WIDTH];
                566 / IN_WIDTH: ping_storage_data_108 <= (fillup_transition == 1'b1) ? i_input_data[566 % IN_WIDTH] : ping_storage_data_108 ^ i_input_data[566 % IN_WIDTH];
                605 / IN_WIDTH: ping_storage_data_108 <= (fillup_transition == 1'b1) ? i_input_data[605 % IN_WIDTH] : ping_storage_data_108 ^ i_input_data[605 % IN_WIDTH];
                675 / IN_WIDTH: ping_storage_data_108 <= (fillup_transition == 1'b1) ? i_input_data[675 % IN_WIDTH] : ping_storage_data_108 ^ i_input_data[675 % IN_WIDTH];
                1056 / IN_WIDTH: ping_storage_data_108 <= (fillup_transition == 1'b1) ? i_input_data[1056 % IN_WIDTH] : ping_storage_data_108 ^ i_input_data[1056 % IN_WIDTH];
                default: ping_storage_data_108 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_108;
                endcase
            end else begin
                case (input_count)
                177 / IN_WIDTH: pong_storage_data_108 <= (fillup_transition == 1'b1) ? i_input_data[177 % IN_WIDTH] : pong_storage_data_108 ^ i_input_data[177 % IN_WIDTH];
                566 / IN_WIDTH: pong_storage_data_108 <= (fillup_transition == 1'b1) ? i_input_data[566 % IN_WIDTH] : pong_storage_data_108 ^ i_input_data[566 % IN_WIDTH];
                605 / IN_WIDTH: pong_storage_data_108 <= (fillup_transition == 1'b1) ? i_input_data[605 % IN_WIDTH] : pong_storage_data_108 ^ i_input_data[605 % IN_WIDTH];
                675 / IN_WIDTH: pong_storage_data_108 <= (fillup_transition == 1'b1) ? i_input_data[675 % IN_WIDTH] : pong_storage_data_108 ^ i_input_data[675 % IN_WIDTH];
                1056 / IN_WIDTH: pong_storage_data_108 <= (fillup_transition == 1'b1) ? i_input_data[1056 % IN_WIDTH] : pong_storage_data_108 ^ i_input_data[1056 % IN_WIDTH];
                default: pong_storage_data_108 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_108;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_108 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_108;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_108 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_108;
            end
        end
    end
end

logic ping_storage_data_109;
logic pong_storage_data_109;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_109 <= 1'b0;
        pong_storage_data_109 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                178 / IN_WIDTH: ping_storage_data_109 <= (fillup_transition == 1'b1) ? i_input_data[178 % IN_WIDTH] : ping_storage_data_109 ^ i_input_data[178 % IN_WIDTH];
                567 / IN_WIDTH: ping_storage_data_109 <= (fillup_transition == 1'b1) ? i_input_data[567 % IN_WIDTH] : ping_storage_data_109 ^ i_input_data[567 % IN_WIDTH];
                606 / IN_WIDTH: ping_storage_data_109 <= (fillup_transition == 1'b1) ? i_input_data[606 % IN_WIDTH] : ping_storage_data_109 ^ i_input_data[606 % IN_WIDTH];
                676 / IN_WIDTH: ping_storage_data_109 <= (fillup_transition == 1'b1) ? i_input_data[676 % IN_WIDTH] : ping_storage_data_109 ^ i_input_data[676 % IN_WIDTH];
                1057 / IN_WIDTH: ping_storage_data_109 <= (fillup_transition == 1'b1) ? i_input_data[1057 % IN_WIDTH] : ping_storage_data_109 ^ i_input_data[1057 % IN_WIDTH];
                default: ping_storage_data_109 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_109;
                endcase
            end else begin
                case (input_count)
                178 / IN_WIDTH: pong_storage_data_109 <= (fillup_transition == 1'b1) ? i_input_data[178 % IN_WIDTH] : pong_storage_data_109 ^ i_input_data[178 % IN_WIDTH];
                567 / IN_WIDTH: pong_storage_data_109 <= (fillup_transition == 1'b1) ? i_input_data[567 % IN_WIDTH] : pong_storage_data_109 ^ i_input_data[567 % IN_WIDTH];
                606 / IN_WIDTH: pong_storage_data_109 <= (fillup_transition == 1'b1) ? i_input_data[606 % IN_WIDTH] : pong_storage_data_109 ^ i_input_data[606 % IN_WIDTH];
                676 / IN_WIDTH: pong_storage_data_109 <= (fillup_transition == 1'b1) ? i_input_data[676 % IN_WIDTH] : pong_storage_data_109 ^ i_input_data[676 % IN_WIDTH];
                1057 / IN_WIDTH: pong_storage_data_109 <= (fillup_transition == 1'b1) ? i_input_data[1057 % IN_WIDTH] : pong_storage_data_109 ^ i_input_data[1057 % IN_WIDTH];
                default: pong_storage_data_109 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_109;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_109 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_109;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_109 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_109;
            end
        end
    end
end

logic ping_storage_data_110;
logic pong_storage_data_110;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_110 <= 1'b0;
        pong_storage_data_110 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                179 / IN_WIDTH: ping_storage_data_110 <= (fillup_transition == 1'b1) ? i_input_data[179 % IN_WIDTH] : ping_storage_data_110 ^ i_input_data[179 % IN_WIDTH];
                568 / IN_WIDTH: ping_storage_data_110 <= (fillup_transition == 1'b1) ? i_input_data[568 % IN_WIDTH] : ping_storage_data_110 ^ i_input_data[568 % IN_WIDTH];
                607 / IN_WIDTH: ping_storage_data_110 <= (fillup_transition == 1'b1) ? i_input_data[607 % IN_WIDTH] : ping_storage_data_110 ^ i_input_data[607 % IN_WIDTH];
                677 / IN_WIDTH: ping_storage_data_110 <= (fillup_transition == 1'b1) ? i_input_data[677 % IN_WIDTH] : ping_storage_data_110 ^ i_input_data[677 % IN_WIDTH];
                1058 / IN_WIDTH: ping_storage_data_110 <= (fillup_transition == 1'b1) ? i_input_data[1058 % IN_WIDTH] : ping_storage_data_110 ^ i_input_data[1058 % IN_WIDTH];
                default: ping_storage_data_110 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_110;
                endcase
            end else begin
                case (input_count)
                179 / IN_WIDTH: pong_storage_data_110 <= (fillup_transition == 1'b1) ? i_input_data[179 % IN_WIDTH] : pong_storage_data_110 ^ i_input_data[179 % IN_WIDTH];
                568 / IN_WIDTH: pong_storage_data_110 <= (fillup_transition == 1'b1) ? i_input_data[568 % IN_WIDTH] : pong_storage_data_110 ^ i_input_data[568 % IN_WIDTH];
                607 / IN_WIDTH: pong_storage_data_110 <= (fillup_transition == 1'b1) ? i_input_data[607 % IN_WIDTH] : pong_storage_data_110 ^ i_input_data[607 % IN_WIDTH];
                677 / IN_WIDTH: pong_storage_data_110 <= (fillup_transition == 1'b1) ? i_input_data[677 % IN_WIDTH] : pong_storage_data_110 ^ i_input_data[677 % IN_WIDTH];
                1058 / IN_WIDTH: pong_storage_data_110 <= (fillup_transition == 1'b1) ? i_input_data[1058 % IN_WIDTH] : pong_storage_data_110 ^ i_input_data[1058 % IN_WIDTH];
                default: pong_storage_data_110 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_110;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_110 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_110;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_110 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_110;
            end
        end
    end
end

logic ping_storage_data_111;
logic pong_storage_data_111;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_111 <= 1'b0;
        pong_storage_data_111 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                180 / IN_WIDTH: ping_storage_data_111 <= (fillup_transition == 1'b1) ? i_input_data[180 % IN_WIDTH] : ping_storage_data_111 ^ i_input_data[180 % IN_WIDTH];
                569 / IN_WIDTH: ping_storage_data_111 <= (fillup_transition == 1'b1) ? i_input_data[569 % IN_WIDTH] : ping_storage_data_111 ^ i_input_data[569 % IN_WIDTH];
                608 / IN_WIDTH: ping_storage_data_111 <= (fillup_transition == 1'b1) ? i_input_data[608 % IN_WIDTH] : ping_storage_data_111 ^ i_input_data[608 % IN_WIDTH];
                678 / IN_WIDTH: ping_storage_data_111 <= (fillup_transition == 1'b1) ? i_input_data[678 % IN_WIDTH] : ping_storage_data_111 ^ i_input_data[678 % IN_WIDTH];
                1059 / IN_WIDTH: ping_storage_data_111 <= (fillup_transition == 1'b1) ? i_input_data[1059 % IN_WIDTH] : ping_storage_data_111 ^ i_input_data[1059 % IN_WIDTH];
                default: ping_storage_data_111 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_111;
                endcase
            end else begin
                case (input_count)
                180 / IN_WIDTH: pong_storage_data_111 <= (fillup_transition == 1'b1) ? i_input_data[180 % IN_WIDTH] : pong_storage_data_111 ^ i_input_data[180 % IN_WIDTH];
                569 / IN_WIDTH: pong_storage_data_111 <= (fillup_transition == 1'b1) ? i_input_data[569 % IN_WIDTH] : pong_storage_data_111 ^ i_input_data[569 % IN_WIDTH];
                608 / IN_WIDTH: pong_storage_data_111 <= (fillup_transition == 1'b1) ? i_input_data[608 % IN_WIDTH] : pong_storage_data_111 ^ i_input_data[608 % IN_WIDTH];
                678 / IN_WIDTH: pong_storage_data_111 <= (fillup_transition == 1'b1) ? i_input_data[678 % IN_WIDTH] : pong_storage_data_111 ^ i_input_data[678 % IN_WIDTH];
                1059 / IN_WIDTH: pong_storage_data_111 <= (fillup_transition == 1'b1) ? i_input_data[1059 % IN_WIDTH] : pong_storage_data_111 ^ i_input_data[1059 % IN_WIDTH];
                default: pong_storage_data_111 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_111;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_111 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_111;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_111 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_111;
            end
        end
    end
end

logic ping_storage_data_112;
logic pong_storage_data_112;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_112 <= 1'b0;
        pong_storage_data_112 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                181 / IN_WIDTH: ping_storage_data_112 <= (fillup_transition == 1'b1) ? i_input_data[181 % IN_WIDTH] : ping_storage_data_112 ^ i_input_data[181 % IN_WIDTH];
                570 / IN_WIDTH: ping_storage_data_112 <= (fillup_transition == 1'b1) ? i_input_data[570 % IN_WIDTH] : ping_storage_data_112 ^ i_input_data[570 % IN_WIDTH];
                609 / IN_WIDTH: ping_storage_data_112 <= (fillup_transition == 1'b1) ? i_input_data[609 % IN_WIDTH] : ping_storage_data_112 ^ i_input_data[609 % IN_WIDTH];
                679 / IN_WIDTH: ping_storage_data_112 <= (fillup_transition == 1'b1) ? i_input_data[679 % IN_WIDTH] : ping_storage_data_112 ^ i_input_data[679 % IN_WIDTH];
                1060 / IN_WIDTH: ping_storage_data_112 <= (fillup_transition == 1'b1) ? i_input_data[1060 % IN_WIDTH] : ping_storage_data_112 ^ i_input_data[1060 % IN_WIDTH];
                default: ping_storage_data_112 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_112;
                endcase
            end else begin
                case (input_count)
                181 / IN_WIDTH: pong_storage_data_112 <= (fillup_transition == 1'b1) ? i_input_data[181 % IN_WIDTH] : pong_storage_data_112 ^ i_input_data[181 % IN_WIDTH];
                570 / IN_WIDTH: pong_storage_data_112 <= (fillup_transition == 1'b1) ? i_input_data[570 % IN_WIDTH] : pong_storage_data_112 ^ i_input_data[570 % IN_WIDTH];
                609 / IN_WIDTH: pong_storage_data_112 <= (fillup_transition == 1'b1) ? i_input_data[609 % IN_WIDTH] : pong_storage_data_112 ^ i_input_data[609 % IN_WIDTH];
                679 / IN_WIDTH: pong_storage_data_112 <= (fillup_transition == 1'b1) ? i_input_data[679 % IN_WIDTH] : pong_storage_data_112 ^ i_input_data[679 % IN_WIDTH];
                1060 / IN_WIDTH: pong_storage_data_112 <= (fillup_transition == 1'b1) ? i_input_data[1060 % IN_WIDTH] : pong_storage_data_112 ^ i_input_data[1060 % IN_WIDTH];
                default: pong_storage_data_112 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_112;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_112 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_112;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_112 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_112;
            end
        end
    end
end

logic ping_storage_data_113;
logic pong_storage_data_113;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_113 <= 1'b0;
        pong_storage_data_113 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                182 / IN_WIDTH: ping_storage_data_113 <= (fillup_transition == 1'b1) ? i_input_data[182 % IN_WIDTH] : ping_storage_data_113 ^ i_input_data[182 % IN_WIDTH];
                571 / IN_WIDTH: ping_storage_data_113 <= (fillup_transition == 1'b1) ? i_input_data[571 % IN_WIDTH] : ping_storage_data_113 ^ i_input_data[571 % IN_WIDTH];
                610 / IN_WIDTH: ping_storage_data_113 <= (fillup_transition == 1'b1) ? i_input_data[610 % IN_WIDTH] : ping_storage_data_113 ^ i_input_data[610 % IN_WIDTH];
                680 / IN_WIDTH: ping_storage_data_113 <= (fillup_transition == 1'b1) ? i_input_data[680 % IN_WIDTH] : ping_storage_data_113 ^ i_input_data[680 % IN_WIDTH];
                1061 / IN_WIDTH: ping_storage_data_113 <= (fillup_transition == 1'b1) ? i_input_data[1061 % IN_WIDTH] : ping_storage_data_113 ^ i_input_data[1061 % IN_WIDTH];
                default: ping_storage_data_113 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_113;
                endcase
            end else begin
                case (input_count)
                182 / IN_WIDTH: pong_storage_data_113 <= (fillup_transition == 1'b1) ? i_input_data[182 % IN_WIDTH] : pong_storage_data_113 ^ i_input_data[182 % IN_WIDTH];
                571 / IN_WIDTH: pong_storage_data_113 <= (fillup_transition == 1'b1) ? i_input_data[571 % IN_WIDTH] : pong_storage_data_113 ^ i_input_data[571 % IN_WIDTH];
                610 / IN_WIDTH: pong_storage_data_113 <= (fillup_transition == 1'b1) ? i_input_data[610 % IN_WIDTH] : pong_storage_data_113 ^ i_input_data[610 % IN_WIDTH];
                680 / IN_WIDTH: pong_storage_data_113 <= (fillup_transition == 1'b1) ? i_input_data[680 % IN_WIDTH] : pong_storage_data_113 ^ i_input_data[680 % IN_WIDTH];
                1061 / IN_WIDTH: pong_storage_data_113 <= (fillup_transition == 1'b1) ? i_input_data[1061 % IN_WIDTH] : pong_storage_data_113 ^ i_input_data[1061 % IN_WIDTH];
                default: pong_storage_data_113 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_113;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_113 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_113;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_113 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_113;
            end
        end
    end
end

logic ping_storage_data_114;
logic pong_storage_data_114;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_114 <= 1'b0;
        pong_storage_data_114 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                183 / IN_WIDTH: ping_storage_data_114 <= (fillup_transition == 1'b1) ? i_input_data[183 % IN_WIDTH] : ping_storage_data_114 ^ i_input_data[183 % IN_WIDTH];
                572 / IN_WIDTH: ping_storage_data_114 <= (fillup_transition == 1'b1) ? i_input_data[572 % IN_WIDTH] : ping_storage_data_114 ^ i_input_data[572 % IN_WIDTH];
                611 / IN_WIDTH: ping_storage_data_114 <= (fillup_transition == 1'b1) ? i_input_data[611 % IN_WIDTH] : ping_storage_data_114 ^ i_input_data[611 % IN_WIDTH];
                681 / IN_WIDTH: ping_storage_data_114 <= (fillup_transition == 1'b1) ? i_input_data[681 % IN_WIDTH] : ping_storage_data_114 ^ i_input_data[681 % IN_WIDTH];
                1062 / IN_WIDTH: ping_storage_data_114 <= (fillup_transition == 1'b1) ? i_input_data[1062 % IN_WIDTH] : ping_storage_data_114 ^ i_input_data[1062 % IN_WIDTH];
                default: ping_storage_data_114 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_114;
                endcase
            end else begin
                case (input_count)
                183 / IN_WIDTH: pong_storage_data_114 <= (fillup_transition == 1'b1) ? i_input_data[183 % IN_WIDTH] : pong_storage_data_114 ^ i_input_data[183 % IN_WIDTH];
                572 / IN_WIDTH: pong_storage_data_114 <= (fillup_transition == 1'b1) ? i_input_data[572 % IN_WIDTH] : pong_storage_data_114 ^ i_input_data[572 % IN_WIDTH];
                611 / IN_WIDTH: pong_storage_data_114 <= (fillup_transition == 1'b1) ? i_input_data[611 % IN_WIDTH] : pong_storage_data_114 ^ i_input_data[611 % IN_WIDTH];
                681 / IN_WIDTH: pong_storage_data_114 <= (fillup_transition == 1'b1) ? i_input_data[681 % IN_WIDTH] : pong_storage_data_114 ^ i_input_data[681 % IN_WIDTH];
                1062 / IN_WIDTH: pong_storage_data_114 <= (fillup_transition == 1'b1) ? i_input_data[1062 % IN_WIDTH] : pong_storage_data_114 ^ i_input_data[1062 % IN_WIDTH];
                default: pong_storage_data_114 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_114;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_114 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_114;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_114 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_114;
            end
        end
    end
end

logic ping_storage_data_115;
logic pong_storage_data_115;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_115 <= 1'b0;
        pong_storage_data_115 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                184 / IN_WIDTH: ping_storage_data_115 <= (fillup_transition == 1'b1) ? i_input_data[184 % IN_WIDTH] : ping_storage_data_115 ^ i_input_data[184 % IN_WIDTH];
                573 / IN_WIDTH: ping_storage_data_115 <= (fillup_transition == 1'b1) ? i_input_data[573 % IN_WIDTH] : ping_storage_data_115 ^ i_input_data[573 % IN_WIDTH];
                612 / IN_WIDTH: ping_storage_data_115 <= (fillup_transition == 1'b1) ? i_input_data[612 % IN_WIDTH] : ping_storage_data_115 ^ i_input_data[612 % IN_WIDTH];
                682 / IN_WIDTH: ping_storage_data_115 <= (fillup_transition == 1'b1) ? i_input_data[682 % IN_WIDTH] : ping_storage_data_115 ^ i_input_data[682 % IN_WIDTH];
                1063 / IN_WIDTH: ping_storage_data_115 <= (fillup_transition == 1'b1) ? i_input_data[1063 % IN_WIDTH] : ping_storage_data_115 ^ i_input_data[1063 % IN_WIDTH];
                default: ping_storage_data_115 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_115;
                endcase
            end else begin
                case (input_count)
                184 / IN_WIDTH: pong_storage_data_115 <= (fillup_transition == 1'b1) ? i_input_data[184 % IN_WIDTH] : pong_storage_data_115 ^ i_input_data[184 % IN_WIDTH];
                573 / IN_WIDTH: pong_storage_data_115 <= (fillup_transition == 1'b1) ? i_input_data[573 % IN_WIDTH] : pong_storage_data_115 ^ i_input_data[573 % IN_WIDTH];
                612 / IN_WIDTH: pong_storage_data_115 <= (fillup_transition == 1'b1) ? i_input_data[612 % IN_WIDTH] : pong_storage_data_115 ^ i_input_data[612 % IN_WIDTH];
                682 / IN_WIDTH: pong_storage_data_115 <= (fillup_transition == 1'b1) ? i_input_data[682 % IN_WIDTH] : pong_storage_data_115 ^ i_input_data[682 % IN_WIDTH];
                1063 / IN_WIDTH: pong_storage_data_115 <= (fillup_transition == 1'b1) ? i_input_data[1063 % IN_WIDTH] : pong_storage_data_115 ^ i_input_data[1063 % IN_WIDTH];
                default: pong_storage_data_115 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_115;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_115 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_115;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_115 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_115;
            end
        end
    end
end

logic ping_storage_data_116;
logic pong_storage_data_116;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_116 <= 1'b0;
        pong_storage_data_116 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                185 / IN_WIDTH: ping_storage_data_116 <= (fillup_transition == 1'b1) ? i_input_data[185 % IN_WIDTH] : ping_storage_data_116 ^ i_input_data[185 % IN_WIDTH];
                574 / IN_WIDTH: ping_storage_data_116 <= (fillup_transition == 1'b1) ? i_input_data[574 % IN_WIDTH] : ping_storage_data_116 ^ i_input_data[574 % IN_WIDTH];
                613 / IN_WIDTH: ping_storage_data_116 <= (fillup_transition == 1'b1) ? i_input_data[613 % IN_WIDTH] : ping_storage_data_116 ^ i_input_data[613 % IN_WIDTH];
                683 / IN_WIDTH: ping_storage_data_116 <= (fillup_transition == 1'b1) ? i_input_data[683 % IN_WIDTH] : ping_storage_data_116 ^ i_input_data[683 % IN_WIDTH];
                1064 / IN_WIDTH: ping_storage_data_116 <= (fillup_transition == 1'b1) ? i_input_data[1064 % IN_WIDTH] : ping_storage_data_116 ^ i_input_data[1064 % IN_WIDTH];
                default: ping_storage_data_116 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_116;
                endcase
            end else begin
                case (input_count)
                185 / IN_WIDTH: pong_storage_data_116 <= (fillup_transition == 1'b1) ? i_input_data[185 % IN_WIDTH] : pong_storage_data_116 ^ i_input_data[185 % IN_WIDTH];
                574 / IN_WIDTH: pong_storage_data_116 <= (fillup_transition == 1'b1) ? i_input_data[574 % IN_WIDTH] : pong_storage_data_116 ^ i_input_data[574 % IN_WIDTH];
                613 / IN_WIDTH: pong_storage_data_116 <= (fillup_transition == 1'b1) ? i_input_data[613 % IN_WIDTH] : pong_storage_data_116 ^ i_input_data[613 % IN_WIDTH];
                683 / IN_WIDTH: pong_storage_data_116 <= (fillup_transition == 1'b1) ? i_input_data[683 % IN_WIDTH] : pong_storage_data_116 ^ i_input_data[683 % IN_WIDTH];
                1064 / IN_WIDTH: pong_storage_data_116 <= (fillup_transition == 1'b1) ? i_input_data[1064 % IN_WIDTH] : pong_storage_data_116 ^ i_input_data[1064 % IN_WIDTH];
                default: pong_storage_data_116 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_116;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_116 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_116;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_116 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_116;
            end
        end
    end
end

logic ping_storage_data_117;
logic pong_storage_data_117;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_117 <= 1'b0;
        pong_storage_data_117 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                186 / IN_WIDTH: ping_storage_data_117 <= (fillup_transition == 1'b1) ? i_input_data[186 % IN_WIDTH] : ping_storage_data_117 ^ i_input_data[186 % IN_WIDTH];
                575 / IN_WIDTH: ping_storage_data_117 <= (fillup_transition == 1'b1) ? i_input_data[575 % IN_WIDTH] : ping_storage_data_117 ^ i_input_data[575 % IN_WIDTH];
                614 / IN_WIDTH: ping_storage_data_117 <= (fillup_transition == 1'b1) ? i_input_data[614 % IN_WIDTH] : ping_storage_data_117 ^ i_input_data[614 % IN_WIDTH];
                684 / IN_WIDTH: ping_storage_data_117 <= (fillup_transition == 1'b1) ? i_input_data[684 % IN_WIDTH] : ping_storage_data_117 ^ i_input_data[684 % IN_WIDTH];
                1065 / IN_WIDTH: ping_storage_data_117 <= (fillup_transition == 1'b1) ? i_input_data[1065 % IN_WIDTH] : ping_storage_data_117 ^ i_input_data[1065 % IN_WIDTH];
                default: ping_storage_data_117 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_117;
                endcase
            end else begin
                case (input_count)
                186 / IN_WIDTH: pong_storage_data_117 <= (fillup_transition == 1'b1) ? i_input_data[186 % IN_WIDTH] : pong_storage_data_117 ^ i_input_data[186 % IN_WIDTH];
                575 / IN_WIDTH: pong_storage_data_117 <= (fillup_transition == 1'b1) ? i_input_data[575 % IN_WIDTH] : pong_storage_data_117 ^ i_input_data[575 % IN_WIDTH];
                614 / IN_WIDTH: pong_storage_data_117 <= (fillup_transition == 1'b1) ? i_input_data[614 % IN_WIDTH] : pong_storage_data_117 ^ i_input_data[614 % IN_WIDTH];
                684 / IN_WIDTH: pong_storage_data_117 <= (fillup_transition == 1'b1) ? i_input_data[684 % IN_WIDTH] : pong_storage_data_117 ^ i_input_data[684 % IN_WIDTH];
                1065 / IN_WIDTH: pong_storage_data_117 <= (fillup_transition == 1'b1) ? i_input_data[1065 % IN_WIDTH] : pong_storage_data_117 ^ i_input_data[1065 % IN_WIDTH];
                default: pong_storage_data_117 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_117;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_117 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_117;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_117 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_117;
            end
        end
    end
end

logic ping_storage_data_118;
logic pong_storage_data_118;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_118 <= 1'b0;
        pong_storage_data_118 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                187 / IN_WIDTH: ping_storage_data_118 <= (fillup_transition == 1'b1) ? i_input_data[187 % IN_WIDTH] : ping_storage_data_118 ^ i_input_data[187 % IN_WIDTH];
                480 / IN_WIDTH: ping_storage_data_118 <= (fillup_transition == 1'b1) ? i_input_data[480 % IN_WIDTH] : ping_storage_data_118 ^ i_input_data[480 % IN_WIDTH];
                615 / IN_WIDTH: ping_storage_data_118 <= (fillup_transition == 1'b1) ? i_input_data[615 % IN_WIDTH] : ping_storage_data_118 ^ i_input_data[615 % IN_WIDTH];
                685 / IN_WIDTH: ping_storage_data_118 <= (fillup_transition == 1'b1) ? i_input_data[685 % IN_WIDTH] : ping_storage_data_118 ^ i_input_data[685 % IN_WIDTH];
                1066 / IN_WIDTH: ping_storage_data_118 <= (fillup_transition == 1'b1) ? i_input_data[1066 % IN_WIDTH] : ping_storage_data_118 ^ i_input_data[1066 % IN_WIDTH];
                default: ping_storage_data_118 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_118;
                endcase
            end else begin
                case (input_count)
                187 / IN_WIDTH: pong_storage_data_118 <= (fillup_transition == 1'b1) ? i_input_data[187 % IN_WIDTH] : pong_storage_data_118 ^ i_input_data[187 % IN_WIDTH];
                480 / IN_WIDTH: pong_storage_data_118 <= (fillup_transition == 1'b1) ? i_input_data[480 % IN_WIDTH] : pong_storage_data_118 ^ i_input_data[480 % IN_WIDTH];
                615 / IN_WIDTH: pong_storage_data_118 <= (fillup_transition == 1'b1) ? i_input_data[615 % IN_WIDTH] : pong_storage_data_118 ^ i_input_data[615 % IN_WIDTH];
                685 / IN_WIDTH: pong_storage_data_118 <= (fillup_transition == 1'b1) ? i_input_data[685 % IN_WIDTH] : pong_storage_data_118 ^ i_input_data[685 % IN_WIDTH];
                1066 / IN_WIDTH: pong_storage_data_118 <= (fillup_transition == 1'b1) ? i_input_data[1066 % IN_WIDTH] : pong_storage_data_118 ^ i_input_data[1066 % IN_WIDTH];
                default: pong_storage_data_118 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_118;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_118 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_118;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_118 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_118;
            end
        end
    end
end

logic ping_storage_data_119;
logic pong_storage_data_119;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_119 <= 1'b0;
        pong_storage_data_119 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                188 / IN_WIDTH: ping_storage_data_119 <= (fillup_transition == 1'b1) ? i_input_data[188 % IN_WIDTH] : ping_storage_data_119 ^ i_input_data[188 % IN_WIDTH];
                481 / IN_WIDTH: ping_storage_data_119 <= (fillup_transition == 1'b1) ? i_input_data[481 % IN_WIDTH] : ping_storage_data_119 ^ i_input_data[481 % IN_WIDTH];
                616 / IN_WIDTH: ping_storage_data_119 <= (fillup_transition == 1'b1) ? i_input_data[616 % IN_WIDTH] : ping_storage_data_119 ^ i_input_data[616 % IN_WIDTH];
                686 / IN_WIDTH: ping_storage_data_119 <= (fillup_transition == 1'b1) ? i_input_data[686 % IN_WIDTH] : ping_storage_data_119 ^ i_input_data[686 % IN_WIDTH];
                1067 / IN_WIDTH: ping_storage_data_119 <= (fillup_transition == 1'b1) ? i_input_data[1067 % IN_WIDTH] : ping_storage_data_119 ^ i_input_data[1067 % IN_WIDTH];
                default: ping_storage_data_119 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_119;
                endcase
            end else begin
                case (input_count)
                188 / IN_WIDTH: pong_storage_data_119 <= (fillup_transition == 1'b1) ? i_input_data[188 % IN_WIDTH] : pong_storage_data_119 ^ i_input_data[188 % IN_WIDTH];
                481 / IN_WIDTH: pong_storage_data_119 <= (fillup_transition == 1'b1) ? i_input_data[481 % IN_WIDTH] : pong_storage_data_119 ^ i_input_data[481 % IN_WIDTH];
                616 / IN_WIDTH: pong_storage_data_119 <= (fillup_transition == 1'b1) ? i_input_data[616 % IN_WIDTH] : pong_storage_data_119 ^ i_input_data[616 % IN_WIDTH];
                686 / IN_WIDTH: pong_storage_data_119 <= (fillup_transition == 1'b1) ? i_input_data[686 % IN_WIDTH] : pong_storage_data_119 ^ i_input_data[686 % IN_WIDTH];
                1067 / IN_WIDTH: pong_storage_data_119 <= (fillup_transition == 1'b1) ? i_input_data[1067 % IN_WIDTH] : pong_storage_data_119 ^ i_input_data[1067 % IN_WIDTH];
                default: pong_storage_data_119 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_119;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_119 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_119;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_119 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_119;
            end
        end
    end
end

logic ping_storage_data_120;
logic pong_storage_data_120;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_120 <= 1'b0;
        pong_storage_data_120 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                189 / IN_WIDTH: ping_storage_data_120 <= (fillup_transition == 1'b1) ? i_input_data[189 % IN_WIDTH] : ping_storage_data_120 ^ i_input_data[189 % IN_WIDTH];
                482 / IN_WIDTH: ping_storage_data_120 <= (fillup_transition == 1'b1) ? i_input_data[482 % IN_WIDTH] : ping_storage_data_120 ^ i_input_data[482 % IN_WIDTH];
                617 / IN_WIDTH: ping_storage_data_120 <= (fillup_transition == 1'b1) ? i_input_data[617 % IN_WIDTH] : ping_storage_data_120 ^ i_input_data[617 % IN_WIDTH];
                687 / IN_WIDTH: ping_storage_data_120 <= (fillup_transition == 1'b1) ? i_input_data[687 % IN_WIDTH] : ping_storage_data_120 ^ i_input_data[687 % IN_WIDTH];
                1068 / IN_WIDTH: ping_storage_data_120 <= (fillup_transition == 1'b1) ? i_input_data[1068 % IN_WIDTH] : ping_storage_data_120 ^ i_input_data[1068 % IN_WIDTH];
                default: ping_storage_data_120 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_120;
                endcase
            end else begin
                case (input_count)
                189 / IN_WIDTH: pong_storage_data_120 <= (fillup_transition == 1'b1) ? i_input_data[189 % IN_WIDTH] : pong_storage_data_120 ^ i_input_data[189 % IN_WIDTH];
                482 / IN_WIDTH: pong_storage_data_120 <= (fillup_transition == 1'b1) ? i_input_data[482 % IN_WIDTH] : pong_storage_data_120 ^ i_input_data[482 % IN_WIDTH];
                617 / IN_WIDTH: pong_storage_data_120 <= (fillup_transition == 1'b1) ? i_input_data[617 % IN_WIDTH] : pong_storage_data_120 ^ i_input_data[617 % IN_WIDTH];
                687 / IN_WIDTH: pong_storage_data_120 <= (fillup_transition == 1'b1) ? i_input_data[687 % IN_WIDTH] : pong_storage_data_120 ^ i_input_data[687 % IN_WIDTH];
                1068 / IN_WIDTH: pong_storage_data_120 <= (fillup_transition == 1'b1) ? i_input_data[1068 % IN_WIDTH] : pong_storage_data_120 ^ i_input_data[1068 % IN_WIDTH];
                default: pong_storage_data_120 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_120;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_120 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_120;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_120 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_120;
            end
        end
    end
end

logic ping_storage_data_121;
logic pong_storage_data_121;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_121 <= 1'b0;
        pong_storage_data_121 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                190 / IN_WIDTH: ping_storage_data_121 <= (fillup_transition == 1'b1) ? i_input_data[190 % IN_WIDTH] : ping_storage_data_121 ^ i_input_data[190 % IN_WIDTH];
                483 / IN_WIDTH: ping_storage_data_121 <= (fillup_transition == 1'b1) ? i_input_data[483 % IN_WIDTH] : ping_storage_data_121 ^ i_input_data[483 % IN_WIDTH];
                618 / IN_WIDTH: ping_storage_data_121 <= (fillup_transition == 1'b1) ? i_input_data[618 % IN_WIDTH] : ping_storage_data_121 ^ i_input_data[618 % IN_WIDTH];
                688 / IN_WIDTH: ping_storage_data_121 <= (fillup_transition == 1'b1) ? i_input_data[688 % IN_WIDTH] : ping_storage_data_121 ^ i_input_data[688 % IN_WIDTH];
                1069 / IN_WIDTH: ping_storage_data_121 <= (fillup_transition == 1'b1) ? i_input_data[1069 % IN_WIDTH] : ping_storage_data_121 ^ i_input_data[1069 % IN_WIDTH];
                default: ping_storage_data_121 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_121;
                endcase
            end else begin
                case (input_count)
                190 / IN_WIDTH: pong_storage_data_121 <= (fillup_transition == 1'b1) ? i_input_data[190 % IN_WIDTH] : pong_storage_data_121 ^ i_input_data[190 % IN_WIDTH];
                483 / IN_WIDTH: pong_storage_data_121 <= (fillup_transition == 1'b1) ? i_input_data[483 % IN_WIDTH] : pong_storage_data_121 ^ i_input_data[483 % IN_WIDTH];
                618 / IN_WIDTH: pong_storage_data_121 <= (fillup_transition == 1'b1) ? i_input_data[618 % IN_WIDTH] : pong_storage_data_121 ^ i_input_data[618 % IN_WIDTH];
                688 / IN_WIDTH: pong_storage_data_121 <= (fillup_transition == 1'b1) ? i_input_data[688 % IN_WIDTH] : pong_storage_data_121 ^ i_input_data[688 % IN_WIDTH];
                1069 / IN_WIDTH: pong_storage_data_121 <= (fillup_transition == 1'b1) ? i_input_data[1069 % IN_WIDTH] : pong_storage_data_121 ^ i_input_data[1069 % IN_WIDTH];
                default: pong_storage_data_121 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_121;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_121 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_121;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_121 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_121;
            end
        end
    end
end

logic ping_storage_data_122;
logic pong_storage_data_122;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_122 <= 1'b0;
        pong_storage_data_122 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                191 / IN_WIDTH: ping_storage_data_122 <= (fillup_transition == 1'b1) ? i_input_data[191 % IN_WIDTH] : ping_storage_data_122 ^ i_input_data[191 % IN_WIDTH];
                484 / IN_WIDTH: ping_storage_data_122 <= (fillup_transition == 1'b1) ? i_input_data[484 % IN_WIDTH] : ping_storage_data_122 ^ i_input_data[484 % IN_WIDTH];
                619 / IN_WIDTH: ping_storage_data_122 <= (fillup_transition == 1'b1) ? i_input_data[619 % IN_WIDTH] : ping_storage_data_122 ^ i_input_data[619 % IN_WIDTH];
                689 / IN_WIDTH: ping_storage_data_122 <= (fillup_transition == 1'b1) ? i_input_data[689 % IN_WIDTH] : ping_storage_data_122 ^ i_input_data[689 % IN_WIDTH];
                1070 / IN_WIDTH: ping_storage_data_122 <= (fillup_transition == 1'b1) ? i_input_data[1070 % IN_WIDTH] : ping_storage_data_122 ^ i_input_data[1070 % IN_WIDTH];
                default: ping_storage_data_122 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_122;
                endcase
            end else begin
                case (input_count)
                191 / IN_WIDTH: pong_storage_data_122 <= (fillup_transition == 1'b1) ? i_input_data[191 % IN_WIDTH] : pong_storage_data_122 ^ i_input_data[191 % IN_WIDTH];
                484 / IN_WIDTH: pong_storage_data_122 <= (fillup_transition == 1'b1) ? i_input_data[484 % IN_WIDTH] : pong_storage_data_122 ^ i_input_data[484 % IN_WIDTH];
                619 / IN_WIDTH: pong_storage_data_122 <= (fillup_transition == 1'b1) ? i_input_data[619 % IN_WIDTH] : pong_storage_data_122 ^ i_input_data[619 % IN_WIDTH];
                689 / IN_WIDTH: pong_storage_data_122 <= (fillup_transition == 1'b1) ? i_input_data[689 % IN_WIDTH] : pong_storage_data_122 ^ i_input_data[689 % IN_WIDTH];
                1070 / IN_WIDTH: pong_storage_data_122 <= (fillup_transition == 1'b1) ? i_input_data[1070 % IN_WIDTH] : pong_storage_data_122 ^ i_input_data[1070 % IN_WIDTH];
                default: pong_storage_data_122 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_122;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_122 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_122;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_122 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_122;
            end
        end
    end
end

logic ping_storage_data_123;
logic pong_storage_data_123;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_123 <= 1'b0;
        pong_storage_data_123 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                96 / IN_WIDTH: ping_storage_data_123 <= (fillup_transition == 1'b1) ? i_input_data[96 % IN_WIDTH] : ping_storage_data_123 ^ i_input_data[96 % IN_WIDTH];
                485 / IN_WIDTH: ping_storage_data_123 <= (fillup_transition == 1'b1) ? i_input_data[485 % IN_WIDTH] : ping_storage_data_123 ^ i_input_data[485 % IN_WIDTH];
                620 / IN_WIDTH: ping_storage_data_123 <= (fillup_transition == 1'b1) ? i_input_data[620 % IN_WIDTH] : ping_storage_data_123 ^ i_input_data[620 % IN_WIDTH];
                690 / IN_WIDTH: ping_storage_data_123 <= (fillup_transition == 1'b1) ? i_input_data[690 % IN_WIDTH] : ping_storage_data_123 ^ i_input_data[690 % IN_WIDTH];
                1071 / IN_WIDTH: ping_storage_data_123 <= (fillup_transition == 1'b1) ? i_input_data[1071 % IN_WIDTH] : ping_storage_data_123 ^ i_input_data[1071 % IN_WIDTH];
                default: ping_storage_data_123 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_123;
                endcase
            end else begin
                case (input_count)
                96 / IN_WIDTH: pong_storage_data_123 <= (fillup_transition == 1'b1) ? i_input_data[96 % IN_WIDTH] : pong_storage_data_123 ^ i_input_data[96 % IN_WIDTH];
                485 / IN_WIDTH: pong_storage_data_123 <= (fillup_transition == 1'b1) ? i_input_data[485 % IN_WIDTH] : pong_storage_data_123 ^ i_input_data[485 % IN_WIDTH];
                620 / IN_WIDTH: pong_storage_data_123 <= (fillup_transition == 1'b1) ? i_input_data[620 % IN_WIDTH] : pong_storage_data_123 ^ i_input_data[620 % IN_WIDTH];
                690 / IN_WIDTH: pong_storage_data_123 <= (fillup_transition == 1'b1) ? i_input_data[690 % IN_WIDTH] : pong_storage_data_123 ^ i_input_data[690 % IN_WIDTH];
                1071 / IN_WIDTH: pong_storage_data_123 <= (fillup_transition == 1'b1) ? i_input_data[1071 % IN_WIDTH] : pong_storage_data_123 ^ i_input_data[1071 % IN_WIDTH];
                default: pong_storage_data_123 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_123;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_123 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_123;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_123 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_123;
            end
        end
    end
end

logic ping_storage_data_124;
logic pong_storage_data_124;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_124 <= 1'b0;
        pong_storage_data_124 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                97 / IN_WIDTH: ping_storage_data_124 <= (fillup_transition == 1'b1) ? i_input_data[97 % IN_WIDTH] : ping_storage_data_124 ^ i_input_data[97 % IN_WIDTH];
                486 / IN_WIDTH: ping_storage_data_124 <= (fillup_transition == 1'b1) ? i_input_data[486 % IN_WIDTH] : ping_storage_data_124 ^ i_input_data[486 % IN_WIDTH];
                621 / IN_WIDTH: ping_storage_data_124 <= (fillup_transition == 1'b1) ? i_input_data[621 % IN_WIDTH] : ping_storage_data_124 ^ i_input_data[621 % IN_WIDTH];
                691 / IN_WIDTH: ping_storage_data_124 <= (fillup_transition == 1'b1) ? i_input_data[691 % IN_WIDTH] : ping_storage_data_124 ^ i_input_data[691 % IN_WIDTH];
                1072 / IN_WIDTH: ping_storage_data_124 <= (fillup_transition == 1'b1) ? i_input_data[1072 % IN_WIDTH] : ping_storage_data_124 ^ i_input_data[1072 % IN_WIDTH];
                default: ping_storage_data_124 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_124;
                endcase
            end else begin
                case (input_count)
                97 / IN_WIDTH: pong_storage_data_124 <= (fillup_transition == 1'b1) ? i_input_data[97 % IN_WIDTH] : pong_storage_data_124 ^ i_input_data[97 % IN_WIDTH];
                486 / IN_WIDTH: pong_storage_data_124 <= (fillup_transition == 1'b1) ? i_input_data[486 % IN_WIDTH] : pong_storage_data_124 ^ i_input_data[486 % IN_WIDTH];
                621 / IN_WIDTH: pong_storage_data_124 <= (fillup_transition == 1'b1) ? i_input_data[621 % IN_WIDTH] : pong_storage_data_124 ^ i_input_data[621 % IN_WIDTH];
                691 / IN_WIDTH: pong_storage_data_124 <= (fillup_transition == 1'b1) ? i_input_data[691 % IN_WIDTH] : pong_storage_data_124 ^ i_input_data[691 % IN_WIDTH];
                1072 / IN_WIDTH: pong_storage_data_124 <= (fillup_transition == 1'b1) ? i_input_data[1072 % IN_WIDTH] : pong_storage_data_124 ^ i_input_data[1072 % IN_WIDTH];
                default: pong_storage_data_124 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_124;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_124 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_124;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_124 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_124;
            end
        end
    end
end

logic ping_storage_data_125;
logic pong_storage_data_125;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_125 <= 1'b0;
        pong_storage_data_125 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                98 / IN_WIDTH: ping_storage_data_125 <= (fillup_transition == 1'b1) ? i_input_data[98 % IN_WIDTH] : ping_storage_data_125 ^ i_input_data[98 % IN_WIDTH];
                487 / IN_WIDTH: ping_storage_data_125 <= (fillup_transition == 1'b1) ? i_input_data[487 % IN_WIDTH] : ping_storage_data_125 ^ i_input_data[487 % IN_WIDTH];
                622 / IN_WIDTH: ping_storage_data_125 <= (fillup_transition == 1'b1) ? i_input_data[622 % IN_WIDTH] : ping_storage_data_125 ^ i_input_data[622 % IN_WIDTH];
                692 / IN_WIDTH: ping_storage_data_125 <= (fillup_transition == 1'b1) ? i_input_data[692 % IN_WIDTH] : ping_storage_data_125 ^ i_input_data[692 % IN_WIDTH];
                1073 / IN_WIDTH: ping_storage_data_125 <= (fillup_transition == 1'b1) ? i_input_data[1073 % IN_WIDTH] : ping_storage_data_125 ^ i_input_data[1073 % IN_WIDTH];
                default: ping_storage_data_125 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_125;
                endcase
            end else begin
                case (input_count)
                98 / IN_WIDTH: pong_storage_data_125 <= (fillup_transition == 1'b1) ? i_input_data[98 % IN_WIDTH] : pong_storage_data_125 ^ i_input_data[98 % IN_WIDTH];
                487 / IN_WIDTH: pong_storage_data_125 <= (fillup_transition == 1'b1) ? i_input_data[487 % IN_WIDTH] : pong_storage_data_125 ^ i_input_data[487 % IN_WIDTH];
                622 / IN_WIDTH: pong_storage_data_125 <= (fillup_transition == 1'b1) ? i_input_data[622 % IN_WIDTH] : pong_storage_data_125 ^ i_input_data[622 % IN_WIDTH];
                692 / IN_WIDTH: pong_storage_data_125 <= (fillup_transition == 1'b1) ? i_input_data[692 % IN_WIDTH] : pong_storage_data_125 ^ i_input_data[692 % IN_WIDTH];
                1073 / IN_WIDTH: pong_storage_data_125 <= (fillup_transition == 1'b1) ? i_input_data[1073 % IN_WIDTH] : pong_storage_data_125 ^ i_input_data[1073 % IN_WIDTH];
                default: pong_storage_data_125 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_125;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_125 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_125;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_125 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_125;
            end
        end
    end
end

logic ping_storage_data_126;
logic pong_storage_data_126;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_126 <= 1'b0;
        pong_storage_data_126 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                99 / IN_WIDTH: ping_storage_data_126 <= (fillup_transition == 1'b1) ? i_input_data[99 % IN_WIDTH] : ping_storage_data_126 ^ i_input_data[99 % IN_WIDTH];
                488 / IN_WIDTH: ping_storage_data_126 <= (fillup_transition == 1'b1) ? i_input_data[488 % IN_WIDTH] : ping_storage_data_126 ^ i_input_data[488 % IN_WIDTH];
                623 / IN_WIDTH: ping_storage_data_126 <= (fillup_transition == 1'b1) ? i_input_data[623 % IN_WIDTH] : ping_storage_data_126 ^ i_input_data[623 % IN_WIDTH];
                693 / IN_WIDTH: ping_storage_data_126 <= (fillup_transition == 1'b1) ? i_input_data[693 % IN_WIDTH] : ping_storage_data_126 ^ i_input_data[693 % IN_WIDTH];
                1074 / IN_WIDTH: ping_storage_data_126 <= (fillup_transition == 1'b1) ? i_input_data[1074 % IN_WIDTH] : ping_storage_data_126 ^ i_input_data[1074 % IN_WIDTH];
                default: ping_storage_data_126 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_126;
                endcase
            end else begin
                case (input_count)
                99 / IN_WIDTH: pong_storage_data_126 <= (fillup_transition == 1'b1) ? i_input_data[99 % IN_WIDTH] : pong_storage_data_126 ^ i_input_data[99 % IN_WIDTH];
                488 / IN_WIDTH: pong_storage_data_126 <= (fillup_transition == 1'b1) ? i_input_data[488 % IN_WIDTH] : pong_storage_data_126 ^ i_input_data[488 % IN_WIDTH];
                623 / IN_WIDTH: pong_storage_data_126 <= (fillup_transition == 1'b1) ? i_input_data[623 % IN_WIDTH] : pong_storage_data_126 ^ i_input_data[623 % IN_WIDTH];
                693 / IN_WIDTH: pong_storage_data_126 <= (fillup_transition == 1'b1) ? i_input_data[693 % IN_WIDTH] : pong_storage_data_126 ^ i_input_data[693 % IN_WIDTH];
                1074 / IN_WIDTH: pong_storage_data_126 <= (fillup_transition == 1'b1) ? i_input_data[1074 % IN_WIDTH] : pong_storage_data_126 ^ i_input_data[1074 % IN_WIDTH];
                default: pong_storage_data_126 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_126;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_126 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_126;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_126 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_126;
            end
        end
    end
end

logic ping_storage_data_127;
logic pong_storage_data_127;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_127 <= 1'b0;
        pong_storage_data_127 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                100 / IN_WIDTH: ping_storage_data_127 <= (fillup_transition == 1'b1) ? i_input_data[100 % IN_WIDTH] : ping_storage_data_127 ^ i_input_data[100 % IN_WIDTH];
                489 / IN_WIDTH: ping_storage_data_127 <= (fillup_transition == 1'b1) ? i_input_data[489 % IN_WIDTH] : ping_storage_data_127 ^ i_input_data[489 % IN_WIDTH];
                624 / IN_WIDTH: ping_storage_data_127 <= (fillup_transition == 1'b1) ? i_input_data[624 % IN_WIDTH] : ping_storage_data_127 ^ i_input_data[624 % IN_WIDTH];
                694 / IN_WIDTH: ping_storage_data_127 <= (fillup_transition == 1'b1) ? i_input_data[694 % IN_WIDTH] : ping_storage_data_127 ^ i_input_data[694 % IN_WIDTH];
                1075 / IN_WIDTH: ping_storage_data_127 <= (fillup_transition == 1'b1) ? i_input_data[1075 % IN_WIDTH] : ping_storage_data_127 ^ i_input_data[1075 % IN_WIDTH];
                default: ping_storage_data_127 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_127;
                endcase
            end else begin
                case (input_count)
                100 / IN_WIDTH: pong_storage_data_127 <= (fillup_transition == 1'b1) ? i_input_data[100 % IN_WIDTH] : pong_storage_data_127 ^ i_input_data[100 % IN_WIDTH];
                489 / IN_WIDTH: pong_storage_data_127 <= (fillup_transition == 1'b1) ? i_input_data[489 % IN_WIDTH] : pong_storage_data_127 ^ i_input_data[489 % IN_WIDTH];
                624 / IN_WIDTH: pong_storage_data_127 <= (fillup_transition == 1'b1) ? i_input_data[624 % IN_WIDTH] : pong_storage_data_127 ^ i_input_data[624 % IN_WIDTH];
                694 / IN_WIDTH: pong_storage_data_127 <= (fillup_transition == 1'b1) ? i_input_data[694 % IN_WIDTH] : pong_storage_data_127 ^ i_input_data[694 % IN_WIDTH];
                1075 / IN_WIDTH: pong_storage_data_127 <= (fillup_transition == 1'b1) ? i_input_data[1075 % IN_WIDTH] : pong_storage_data_127 ^ i_input_data[1075 % IN_WIDTH];
                default: pong_storage_data_127 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_127;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_127 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_127;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_127 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_127;
            end
        end
    end
end

logic ping_storage_data_128;
logic pong_storage_data_128;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_128 <= 1'b0;
        pong_storage_data_128 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                101 / IN_WIDTH: ping_storage_data_128 <= (fillup_transition == 1'b1) ? i_input_data[101 % IN_WIDTH] : ping_storage_data_128 ^ i_input_data[101 % IN_WIDTH];
                490 / IN_WIDTH: ping_storage_data_128 <= (fillup_transition == 1'b1) ? i_input_data[490 % IN_WIDTH] : ping_storage_data_128 ^ i_input_data[490 % IN_WIDTH];
                625 / IN_WIDTH: ping_storage_data_128 <= (fillup_transition == 1'b1) ? i_input_data[625 % IN_WIDTH] : ping_storage_data_128 ^ i_input_data[625 % IN_WIDTH];
                695 / IN_WIDTH: ping_storage_data_128 <= (fillup_transition == 1'b1) ? i_input_data[695 % IN_WIDTH] : ping_storage_data_128 ^ i_input_data[695 % IN_WIDTH];
                1076 / IN_WIDTH: ping_storage_data_128 <= (fillup_transition == 1'b1) ? i_input_data[1076 % IN_WIDTH] : ping_storage_data_128 ^ i_input_data[1076 % IN_WIDTH];
                default: ping_storage_data_128 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_128;
                endcase
            end else begin
                case (input_count)
                101 / IN_WIDTH: pong_storage_data_128 <= (fillup_transition == 1'b1) ? i_input_data[101 % IN_WIDTH] : pong_storage_data_128 ^ i_input_data[101 % IN_WIDTH];
                490 / IN_WIDTH: pong_storage_data_128 <= (fillup_transition == 1'b1) ? i_input_data[490 % IN_WIDTH] : pong_storage_data_128 ^ i_input_data[490 % IN_WIDTH];
                625 / IN_WIDTH: pong_storage_data_128 <= (fillup_transition == 1'b1) ? i_input_data[625 % IN_WIDTH] : pong_storage_data_128 ^ i_input_data[625 % IN_WIDTH];
                695 / IN_WIDTH: pong_storage_data_128 <= (fillup_transition == 1'b1) ? i_input_data[695 % IN_WIDTH] : pong_storage_data_128 ^ i_input_data[695 % IN_WIDTH];
                1076 / IN_WIDTH: pong_storage_data_128 <= (fillup_transition == 1'b1) ? i_input_data[1076 % IN_WIDTH] : pong_storage_data_128 ^ i_input_data[1076 % IN_WIDTH];
                default: pong_storage_data_128 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_128;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_128 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_128;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_128 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_128;
            end
        end
    end
end

logic ping_storage_data_129;
logic pong_storage_data_129;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_129 <= 1'b0;
        pong_storage_data_129 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                102 / IN_WIDTH: ping_storage_data_129 <= (fillup_transition == 1'b1) ? i_input_data[102 % IN_WIDTH] : ping_storage_data_129 ^ i_input_data[102 % IN_WIDTH];
                491 / IN_WIDTH: ping_storage_data_129 <= (fillup_transition == 1'b1) ? i_input_data[491 % IN_WIDTH] : ping_storage_data_129 ^ i_input_data[491 % IN_WIDTH];
                626 / IN_WIDTH: ping_storage_data_129 <= (fillup_transition == 1'b1) ? i_input_data[626 % IN_WIDTH] : ping_storage_data_129 ^ i_input_data[626 % IN_WIDTH];
                696 / IN_WIDTH: ping_storage_data_129 <= (fillup_transition == 1'b1) ? i_input_data[696 % IN_WIDTH] : ping_storage_data_129 ^ i_input_data[696 % IN_WIDTH];
                1077 / IN_WIDTH: ping_storage_data_129 <= (fillup_transition == 1'b1) ? i_input_data[1077 % IN_WIDTH] : ping_storage_data_129 ^ i_input_data[1077 % IN_WIDTH];
                default: ping_storage_data_129 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_129;
                endcase
            end else begin
                case (input_count)
                102 / IN_WIDTH: pong_storage_data_129 <= (fillup_transition == 1'b1) ? i_input_data[102 % IN_WIDTH] : pong_storage_data_129 ^ i_input_data[102 % IN_WIDTH];
                491 / IN_WIDTH: pong_storage_data_129 <= (fillup_transition == 1'b1) ? i_input_data[491 % IN_WIDTH] : pong_storage_data_129 ^ i_input_data[491 % IN_WIDTH];
                626 / IN_WIDTH: pong_storage_data_129 <= (fillup_transition == 1'b1) ? i_input_data[626 % IN_WIDTH] : pong_storage_data_129 ^ i_input_data[626 % IN_WIDTH];
                696 / IN_WIDTH: pong_storage_data_129 <= (fillup_transition == 1'b1) ? i_input_data[696 % IN_WIDTH] : pong_storage_data_129 ^ i_input_data[696 % IN_WIDTH];
                1077 / IN_WIDTH: pong_storage_data_129 <= (fillup_transition == 1'b1) ? i_input_data[1077 % IN_WIDTH] : pong_storage_data_129 ^ i_input_data[1077 % IN_WIDTH];
                default: pong_storage_data_129 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_129;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_129 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_129;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_129 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_129;
            end
        end
    end
end

logic ping_storage_data_130;
logic pong_storage_data_130;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_130 <= 1'b0;
        pong_storage_data_130 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                103 / IN_WIDTH: ping_storage_data_130 <= (fillup_transition == 1'b1) ? i_input_data[103 % IN_WIDTH] : ping_storage_data_130 ^ i_input_data[103 % IN_WIDTH];
                492 / IN_WIDTH: ping_storage_data_130 <= (fillup_transition == 1'b1) ? i_input_data[492 % IN_WIDTH] : ping_storage_data_130 ^ i_input_data[492 % IN_WIDTH];
                627 / IN_WIDTH: ping_storage_data_130 <= (fillup_transition == 1'b1) ? i_input_data[627 % IN_WIDTH] : ping_storage_data_130 ^ i_input_data[627 % IN_WIDTH];
                697 / IN_WIDTH: ping_storage_data_130 <= (fillup_transition == 1'b1) ? i_input_data[697 % IN_WIDTH] : ping_storage_data_130 ^ i_input_data[697 % IN_WIDTH];
                1078 / IN_WIDTH: ping_storage_data_130 <= (fillup_transition == 1'b1) ? i_input_data[1078 % IN_WIDTH] : ping_storage_data_130 ^ i_input_data[1078 % IN_WIDTH];
                default: ping_storage_data_130 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_130;
                endcase
            end else begin
                case (input_count)
                103 / IN_WIDTH: pong_storage_data_130 <= (fillup_transition == 1'b1) ? i_input_data[103 % IN_WIDTH] : pong_storage_data_130 ^ i_input_data[103 % IN_WIDTH];
                492 / IN_WIDTH: pong_storage_data_130 <= (fillup_transition == 1'b1) ? i_input_data[492 % IN_WIDTH] : pong_storage_data_130 ^ i_input_data[492 % IN_WIDTH];
                627 / IN_WIDTH: pong_storage_data_130 <= (fillup_transition == 1'b1) ? i_input_data[627 % IN_WIDTH] : pong_storage_data_130 ^ i_input_data[627 % IN_WIDTH];
                697 / IN_WIDTH: pong_storage_data_130 <= (fillup_transition == 1'b1) ? i_input_data[697 % IN_WIDTH] : pong_storage_data_130 ^ i_input_data[697 % IN_WIDTH];
                1078 / IN_WIDTH: pong_storage_data_130 <= (fillup_transition == 1'b1) ? i_input_data[1078 % IN_WIDTH] : pong_storage_data_130 ^ i_input_data[1078 % IN_WIDTH];
                default: pong_storage_data_130 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_130;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_130 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_130;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_130 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_130;
            end
        end
    end
end

logic ping_storage_data_131;
logic pong_storage_data_131;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_131 <= 1'b0;
        pong_storage_data_131 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                104 / IN_WIDTH: ping_storage_data_131 <= (fillup_transition == 1'b1) ? i_input_data[104 % IN_WIDTH] : ping_storage_data_131 ^ i_input_data[104 % IN_WIDTH];
                493 / IN_WIDTH: ping_storage_data_131 <= (fillup_transition == 1'b1) ? i_input_data[493 % IN_WIDTH] : ping_storage_data_131 ^ i_input_data[493 % IN_WIDTH];
                628 / IN_WIDTH: ping_storage_data_131 <= (fillup_transition == 1'b1) ? i_input_data[628 % IN_WIDTH] : ping_storage_data_131 ^ i_input_data[628 % IN_WIDTH];
                698 / IN_WIDTH: ping_storage_data_131 <= (fillup_transition == 1'b1) ? i_input_data[698 % IN_WIDTH] : ping_storage_data_131 ^ i_input_data[698 % IN_WIDTH];
                1079 / IN_WIDTH: ping_storage_data_131 <= (fillup_transition == 1'b1) ? i_input_data[1079 % IN_WIDTH] : ping_storage_data_131 ^ i_input_data[1079 % IN_WIDTH];
                default: ping_storage_data_131 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_131;
                endcase
            end else begin
                case (input_count)
                104 / IN_WIDTH: pong_storage_data_131 <= (fillup_transition == 1'b1) ? i_input_data[104 % IN_WIDTH] : pong_storage_data_131 ^ i_input_data[104 % IN_WIDTH];
                493 / IN_WIDTH: pong_storage_data_131 <= (fillup_transition == 1'b1) ? i_input_data[493 % IN_WIDTH] : pong_storage_data_131 ^ i_input_data[493 % IN_WIDTH];
                628 / IN_WIDTH: pong_storage_data_131 <= (fillup_transition == 1'b1) ? i_input_data[628 % IN_WIDTH] : pong_storage_data_131 ^ i_input_data[628 % IN_WIDTH];
                698 / IN_WIDTH: pong_storage_data_131 <= (fillup_transition == 1'b1) ? i_input_data[698 % IN_WIDTH] : pong_storage_data_131 ^ i_input_data[698 % IN_WIDTH];
                1079 / IN_WIDTH: pong_storage_data_131 <= (fillup_transition == 1'b1) ? i_input_data[1079 % IN_WIDTH] : pong_storage_data_131 ^ i_input_data[1079 % IN_WIDTH];
                default: pong_storage_data_131 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_131;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_131 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_131;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_131 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_131;
            end
        end
    end
end

logic ping_storage_data_132;
logic pong_storage_data_132;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_132 <= 1'b0;
        pong_storage_data_132 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                105 / IN_WIDTH: ping_storage_data_132 <= (fillup_transition == 1'b1) ? i_input_data[105 % IN_WIDTH] : ping_storage_data_132 ^ i_input_data[105 % IN_WIDTH];
                494 / IN_WIDTH: ping_storage_data_132 <= (fillup_transition == 1'b1) ? i_input_data[494 % IN_WIDTH] : ping_storage_data_132 ^ i_input_data[494 % IN_WIDTH];
                629 / IN_WIDTH: ping_storage_data_132 <= (fillup_transition == 1'b1) ? i_input_data[629 % IN_WIDTH] : ping_storage_data_132 ^ i_input_data[629 % IN_WIDTH];
                699 / IN_WIDTH: ping_storage_data_132 <= (fillup_transition == 1'b1) ? i_input_data[699 % IN_WIDTH] : ping_storage_data_132 ^ i_input_data[699 % IN_WIDTH];
                1080 / IN_WIDTH: ping_storage_data_132 <= (fillup_transition == 1'b1) ? i_input_data[1080 % IN_WIDTH] : ping_storage_data_132 ^ i_input_data[1080 % IN_WIDTH];
                default: ping_storage_data_132 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_132;
                endcase
            end else begin
                case (input_count)
                105 / IN_WIDTH: pong_storage_data_132 <= (fillup_transition == 1'b1) ? i_input_data[105 % IN_WIDTH] : pong_storage_data_132 ^ i_input_data[105 % IN_WIDTH];
                494 / IN_WIDTH: pong_storage_data_132 <= (fillup_transition == 1'b1) ? i_input_data[494 % IN_WIDTH] : pong_storage_data_132 ^ i_input_data[494 % IN_WIDTH];
                629 / IN_WIDTH: pong_storage_data_132 <= (fillup_transition == 1'b1) ? i_input_data[629 % IN_WIDTH] : pong_storage_data_132 ^ i_input_data[629 % IN_WIDTH];
                699 / IN_WIDTH: pong_storage_data_132 <= (fillup_transition == 1'b1) ? i_input_data[699 % IN_WIDTH] : pong_storage_data_132 ^ i_input_data[699 % IN_WIDTH];
                1080 / IN_WIDTH: pong_storage_data_132 <= (fillup_transition == 1'b1) ? i_input_data[1080 % IN_WIDTH] : pong_storage_data_132 ^ i_input_data[1080 % IN_WIDTH];
                default: pong_storage_data_132 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_132;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_132 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_132;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_132 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_132;
            end
        end
    end
end

logic ping_storage_data_133;
logic pong_storage_data_133;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_133 <= 1'b0;
        pong_storage_data_133 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                106 / IN_WIDTH: ping_storage_data_133 <= (fillup_transition == 1'b1) ? i_input_data[106 % IN_WIDTH] : ping_storage_data_133 ^ i_input_data[106 % IN_WIDTH];
                495 / IN_WIDTH: ping_storage_data_133 <= (fillup_transition == 1'b1) ? i_input_data[495 % IN_WIDTH] : ping_storage_data_133 ^ i_input_data[495 % IN_WIDTH];
                630 / IN_WIDTH: ping_storage_data_133 <= (fillup_transition == 1'b1) ? i_input_data[630 % IN_WIDTH] : ping_storage_data_133 ^ i_input_data[630 % IN_WIDTH];
                700 / IN_WIDTH: ping_storage_data_133 <= (fillup_transition == 1'b1) ? i_input_data[700 % IN_WIDTH] : ping_storage_data_133 ^ i_input_data[700 % IN_WIDTH];
                1081 / IN_WIDTH: ping_storage_data_133 <= (fillup_transition == 1'b1) ? i_input_data[1081 % IN_WIDTH] : ping_storage_data_133 ^ i_input_data[1081 % IN_WIDTH];
                default: ping_storage_data_133 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_133;
                endcase
            end else begin
                case (input_count)
                106 / IN_WIDTH: pong_storage_data_133 <= (fillup_transition == 1'b1) ? i_input_data[106 % IN_WIDTH] : pong_storage_data_133 ^ i_input_data[106 % IN_WIDTH];
                495 / IN_WIDTH: pong_storage_data_133 <= (fillup_transition == 1'b1) ? i_input_data[495 % IN_WIDTH] : pong_storage_data_133 ^ i_input_data[495 % IN_WIDTH];
                630 / IN_WIDTH: pong_storage_data_133 <= (fillup_transition == 1'b1) ? i_input_data[630 % IN_WIDTH] : pong_storage_data_133 ^ i_input_data[630 % IN_WIDTH];
                700 / IN_WIDTH: pong_storage_data_133 <= (fillup_transition == 1'b1) ? i_input_data[700 % IN_WIDTH] : pong_storage_data_133 ^ i_input_data[700 % IN_WIDTH];
                1081 / IN_WIDTH: pong_storage_data_133 <= (fillup_transition == 1'b1) ? i_input_data[1081 % IN_WIDTH] : pong_storage_data_133 ^ i_input_data[1081 % IN_WIDTH];
                default: pong_storage_data_133 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_133;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_133 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_133;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_133 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_133;
            end
        end
    end
end

logic ping_storage_data_134;
logic pong_storage_data_134;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_134 <= 1'b0;
        pong_storage_data_134 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                107 / IN_WIDTH: ping_storage_data_134 <= (fillup_transition == 1'b1) ? i_input_data[107 % IN_WIDTH] : ping_storage_data_134 ^ i_input_data[107 % IN_WIDTH];
                496 / IN_WIDTH: ping_storage_data_134 <= (fillup_transition == 1'b1) ? i_input_data[496 % IN_WIDTH] : ping_storage_data_134 ^ i_input_data[496 % IN_WIDTH];
                631 / IN_WIDTH: ping_storage_data_134 <= (fillup_transition == 1'b1) ? i_input_data[631 % IN_WIDTH] : ping_storage_data_134 ^ i_input_data[631 % IN_WIDTH];
                701 / IN_WIDTH: ping_storage_data_134 <= (fillup_transition == 1'b1) ? i_input_data[701 % IN_WIDTH] : ping_storage_data_134 ^ i_input_data[701 % IN_WIDTH];
                1082 / IN_WIDTH: ping_storage_data_134 <= (fillup_transition == 1'b1) ? i_input_data[1082 % IN_WIDTH] : ping_storage_data_134 ^ i_input_data[1082 % IN_WIDTH];
                default: ping_storage_data_134 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_134;
                endcase
            end else begin
                case (input_count)
                107 / IN_WIDTH: pong_storage_data_134 <= (fillup_transition == 1'b1) ? i_input_data[107 % IN_WIDTH] : pong_storage_data_134 ^ i_input_data[107 % IN_WIDTH];
                496 / IN_WIDTH: pong_storage_data_134 <= (fillup_transition == 1'b1) ? i_input_data[496 % IN_WIDTH] : pong_storage_data_134 ^ i_input_data[496 % IN_WIDTH];
                631 / IN_WIDTH: pong_storage_data_134 <= (fillup_transition == 1'b1) ? i_input_data[631 % IN_WIDTH] : pong_storage_data_134 ^ i_input_data[631 % IN_WIDTH];
                701 / IN_WIDTH: pong_storage_data_134 <= (fillup_transition == 1'b1) ? i_input_data[701 % IN_WIDTH] : pong_storage_data_134 ^ i_input_data[701 % IN_WIDTH];
                1082 / IN_WIDTH: pong_storage_data_134 <= (fillup_transition == 1'b1) ? i_input_data[1082 % IN_WIDTH] : pong_storage_data_134 ^ i_input_data[1082 % IN_WIDTH];
                default: pong_storage_data_134 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_134;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_134 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_134;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_134 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_134;
            end
        end
    end
end

logic ping_storage_data_135;
logic pong_storage_data_135;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_135 <= 1'b0;
        pong_storage_data_135 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                108 / IN_WIDTH: ping_storage_data_135 <= (fillup_transition == 1'b1) ? i_input_data[108 % IN_WIDTH] : ping_storage_data_135 ^ i_input_data[108 % IN_WIDTH];
                497 / IN_WIDTH: ping_storage_data_135 <= (fillup_transition == 1'b1) ? i_input_data[497 % IN_WIDTH] : ping_storage_data_135 ^ i_input_data[497 % IN_WIDTH];
                632 / IN_WIDTH: ping_storage_data_135 <= (fillup_transition == 1'b1) ? i_input_data[632 % IN_WIDTH] : ping_storage_data_135 ^ i_input_data[632 % IN_WIDTH];
                702 / IN_WIDTH: ping_storage_data_135 <= (fillup_transition == 1'b1) ? i_input_data[702 % IN_WIDTH] : ping_storage_data_135 ^ i_input_data[702 % IN_WIDTH];
                1083 / IN_WIDTH: ping_storage_data_135 <= (fillup_transition == 1'b1) ? i_input_data[1083 % IN_WIDTH] : ping_storage_data_135 ^ i_input_data[1083 % IN_WIDTH];
                default: ping_storage_data_135 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_135;
                endcase
            end else begin
                case (input_count)
                108 / IN_WIDTH: pong_storage_data_135 <= (fillup_transition == 1'b1) ? i_input_data[108 % IN_WIDTH] : pong_storage_data_135 ^ i_input_data[108 % IN_WIDTH];
                497 / IN_WIDTH: pong_storage_data_135 <= (fillup_transition == 1'b1) ? i_input_data[497 % IN_WIDTH] : pong_storage_data_135 ^ i_input_data[497 % IN_WIDTH];
                632 / IN_WIDTH: pong_storage_data_135 <= (fillup_transition == 1'b1) ? i_input_data[632 % IN_WIDTH] : pong_storage_data_135 ^ i_input_data[632 % IN_WIDTH];
                702 / IN_WIDTH: pong_storage_data_135 <= (fillup_transition == 1'b1) ? i_input_data[702 % IN_WIDTH] : pong_storage_data_135 ^ i_input_data[702 % IN_WIDTH];
                1083 / IN_WIDTH: pong_storage_data_135 <= (fillup_transition == 1'b1) ? i_input_data[1083 % IN_WIDTH] : pong_storage_data_135 ^ i_input_data[1083 % IN_WIDTH];
                default: pong_storage_data_135 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_135;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_135 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_135;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_135 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_135;
            end
        end
    end
end

logic ping_storage_data_136;
logic pong_storage_data_136;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_136 <= 1'b0;
        pong_storage_data_136 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                109 / IN_WIDTH: ping_storage_data_136 <= (fillup_transition == 1'b1) ? i_input_data[109 % IN_WIDTH] : ping_storage_data_136 ^ i_input_data[109 % IN_WIDTH];
                498 / IN_WIDTH: ping_storage_data_136 <= (fillup_transition == 1'b1) ? i_input_data[498 % IN_WIDTH] : ping_storage_data_136 ^ i_input_data[498 % IN_WIDTH];
                633 / IN_WIDTH: ping_storage_data_136 <= (fillup_transition == 1'b1) ? i_input_data[633 % IN_WIDTH] : ping_storage_data_136 ^ i_input_data[633 % IN_WIDTH];
                703 / IN_WIDTH: ping_storage_data_136 <= (fillup_transition == 1'b1) ? i_input_data[703 % IN_WIDTH] : ping_storage_data_136 ^ i_input_data[703 % IN_WIDTH];
                1084 / IN_WIDTH: ping_storage_data_136 <= (fillup_transition == 1'b1) ? i_input_data[1084 % IN_WIDTH] : ping_storage_data_136 ^ i_input_data[1084 % IN_WIDTH];
                default: ping_storage_data_136 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_136;
                endcase
            end else begin
                case (input_count)
                109 / IN_WIDTH: pong_storage_data_136 <= (fillup_transition == 1'b1) ? i_input_data[109 % IN_WIDTH] : pong_storage_data_136 ^ i_input_data[109 % IN_WIDTH];
                498 / IN_WIDTH: pong_storage_data_136 <= (fillup_transition == 1'b1) ? i_input_data[498 % IN_WIDTH] : pong_storage_data_136 ^ i_input_data[498 % IN_WIDTH];
                633 / IN_WIDTH: pong_storage_data_136 <= (fillup_transition == 1'b1) ? i_input_data[633 % IN_WIDTH] : pong_storage_data_136 ^ i_input_data[633 % IN_WIDTH];
                703 / IN_WIDTH: pong_storage_data_136 <= (fillup_transition == 1'b1) ? i_input_data[703 % IN_WIDTH] : pong_storage_data_136 ^ i_input_data[703 % IN_WIDTH];
                1084 / IN_WIDTH: pong_storage_data_136 <= (fillup_transition == 1'b1) ? i_input_data[1084 % IN_WIDTH] : pong_storage_data_136 ^ i_input_data[1084 % IN_WIDTH];
                default: pong_storage_data_136 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_136;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_136 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_136;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_136 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_136;
            end
        end
    end
end

logic ping_storage_data_137;
logic pong_storage_data_137;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_137 <= 1'b0;
        pong_storage_data_137 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                110 / IN_WIDTH: ping_storage_data_137 <= (fillup_transition == 1'b1) ? i_input_data[110 % IN_WIDTH] : ping_storage_data_137 ^ i_input_data[110 % IN_WIDTH];
                499 / IN_WIDTH: ping_storage_data_137 <= (fillup_transition == 1'b1) ? i_input_data[499 % IN_WIDTH] : ping_storage_data_137 ^ i_input_data[499 % IN_WIDTH];
                634 / IN_WIDTH: ping_storage_data_137 <= (fillup_transition == 1'b1) ? i_input_data[634 % IN_WIDTH] : ping_storage_data_137 ^ i_input_data[634 % IN_WIDTH];
                704 / IN_WIDTH: ping_storage_data_137 <= (fillup_transition == 1'b1) ? i_input_data[704 % IN_WIDTH] : ping_storage_data_137 ^ i_input_data[704 % IN_WIDTH];
                1085 / IN_WIDTH: ping_storage_data_137 <= (fillup_transition == 1'b1) ? i_input_data[1085 % IN_WIDTH] : ping_storage_data_137 ^ i_input_data[1085 % IN_WIDTH];
                default: ping_storage_data_137 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_137;
                endcase
            end else begin
                case (input_count)
                110 / IN_WIDTH: pong_storage_data_137 <= (fillup_transition == 1'b1) ? i_input_data[110 % IN_WIDTH] : pong_storage_data_137 ^ i_input_data[110 % IN_WIDTH];
                499 / IN_WIDTH: pong_storage_data_137 <= (fillup_transition == 1'b1) ? i_input_data[499 % IN_WIDTH] : pong_storage_data_137 ^ i_input_data[499 % IN_WIDTH];
                634 / IN_WIDTH: pong_storage_data_137 <= (fillup_transition == 1'b1) ? i_input_data[634 % IN_WIDTH] : pong_storage_data_137 ^ i_input_data[634 % IN_WIDTH];
                704 / IN_WIDTH: pong_storage_data_137 <= (fillup_transition == 1'b1) ? i_input_data[704 % IN_WIDTH] : pong_storage_data_137 ^ i_input_data[704 % IN_WIDTH];
                1085 / IN_WIDTH: pong_storage_data_137 <= (fillup_transition == 1'b1) ? i_input_data[1085 % IN_WIDTH] : pong_storage_data_137 ^ i_input_data[1085 % IN_WIDTH];
                default: pong_storage_data_137 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_137;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_137 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_137;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_137 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_137;
            end
        end
    end
end

logic ping_storage_data_138;
logic pong_storage_data_138;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_138 <= 1'b0;
        pong_storage_data_138 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                111 / IN_WIDTH: ping_storage_data_138 <= (fillup_transition == 1'b1) ? i_input_data[111 % IN_WIDTH] : ping_storage_data_138 ^ i_input_data[111 % IN_WIDTH];
                500 / IN_WIDTH: ping_storage_data_138 <= (fillup_transition == 1'b1) ? i_input_data[500 % IN_WIDTH] : ping_storage_data_138 ^ i_input_data[500 % IN_WIDTH];
                635 / IN_WIDTH: ping_storage_data_138 <= (fillup_transition == 1'b1) ? i_input_data[635 % IN_WIDTH] : ping_storage_data_138 ^ i_input_data[635 % IN_WIDTH];
                705 / IN_WIDTH: ping_storage_data_138 <= (fillup_transition == 1'b1) ? i_input_data[705 % IN_WIDTH] : ping_storage_data_138 ^ i_input_data[705 % IN_WIDTH];
                1086 / IN_WIDTH: ping_storage_data_138 <= (fillup_transition == 1'b1) ? i_input_data[1086 % IN_WIDTH] : ping_storage_data_138 ^ i_input_data[1086 % IN_WIDTH];
                default: ping_storage_data_138 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_138;
                endcase
            end else begin
                case (input_count)
                111 / IN_WIDTH: pong_storage_data_138 <= (fillup_transition == 1'b1) ? i_input_data[111 % IN_WIDTH] : pong_storage_data_138 ^ i_input_data[111 % IN_WIDTH];
                500 / IN_WIDTH: pong_storage_data_138 <= (fillup_transition == 1'b1) ? i_input_data[500 % IN_WIDTH] : pong_storage_data_138 ^ i_input_data[500 % IN_WIDTH];
                635 / IN_WIDTH: pong_storage_data_138 <= (fillup_transition == 1'b1) ? i_input_data[635 % IN_WIDTH] : pong_storage_data_138 ^ i_input_data[635 % IN_WIDTH];
                705 / IN_WIDTH: pong_storage_data_138 <= (fillup_transition == 1'b1) ? i_input_data[705 % IN_WIDTH] : pong_storage_data_138 ^ i_input_data[705 % IN_WIDTH];
                1086 / IN_WIDTH: pong_storage_data_138 <= (fillup_transition == 1'b1) ? i_input_data[1086 % IN_WIDTH] : pong_storage_data_138 ^ i_input_data[1086 % IN_WIDTH];
                default: pong_storage_data_138 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_138;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_138 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_138;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_138 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_138;
            end
        end
    end
end

logic ping_storage_data_139;
logic pong_storage_data_139;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_139 <= 1'b0;
        pong_storage_data_139 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                112 / IN_WIDTH: ping_storage_data_139 <= (fillup_transition == 1'b1) ? i_input_data[112 % IN_WIDTH] : ping_storage_data_139 ^ i_input_data[112 % IN_WIDTH];
                501 / IN_WIDTH: ping_storage_data_139 <= (fillup_transition == 1'b1) ? i_input_data[501 % IN_WIDTH] : ping_storage_data_139 ^ i_input_data[501 % IN_WIDTH];
                636 / IN_WIDTH: ping_storage_data_139 <= (fillup_transition == 1'b1) ? i_input_data[636 % IN_WIDTH] : ping_storage_data_139 ^ i_input_data[636 % IN_WIDTH];
                706 / IN_WIDTH: ping_storage_data_139 <= (fillup_transition == 1'b1) ? i_input_data[706 % IN_WIDTH] : ping_storage_data_139 ^ i_input_data[706 % IN_WIDTH];
                1087 / IN_WIDTH: ping_storage_data_139 <= (fillup_transition == 1'b1) ? i_input_data[1087 % IN_WIDTH] : ping_storage_data_139 ^ i_input_data[1087 % IN_WIDTH];
                default: ping_storage_data_139 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_139;
                endcase
            end else begin
                case (input_count)
                112 / IN_WIDTH: pong_storage_data_139 <= (fillup_transition == 1'b1) ? i_input_data[112 % IN_WIDTH] : pong_storage_data_139 ^ i_input_data[112 % IN_WIDTH];
                501 / IN_WIDTH: pong_storage_data_139 <= (fillup_transition == 1'b1) ? i_input_data[501 % IN_WIDTH] : pong_storage_data_139 ^ i_input_data[501 % IN_WIDTH];
                636 / IN_WIDTH: pong_storage_data_139 <= (fillup_transition == 1'b1) ? i_input_data[636 % IN_WIDTH] : pong_storage_data_139 ^ i_input_data[636 % IN_WIDTH];
                706 / IN_WIDTH: pong_storage_data_139 <= (fillup_transition == 1'b1) ? i_input_data[706 % IN_WIDTH] : pong_storage_data_139 ^ i_input_data[706 % IN_WIDTH];
                1087 / IN_WIDTH: pong_storage_data_139 <= (fillup_transition == 1'b1) ? i_input_data[1087 % IN_WIDTH] : pong_storage_data_139 ^ i_input_data[1087 % IN_WIDTH];
                default: pong_storage_data_139 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_139;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_139 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_139;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_139 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_139;
            end
        end
    end
end

logic ping_storage_data_140;
logic pong_storage_data_140;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_140 <= 1'b0;
        pong_storage_data_140 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                113 / IN_WIDTH: ping_storage_data_140 <= (fillup_transition == 1'b1) ? i_input_data[113 % IN_WIDTH] : ping_storage_data_140 ^ i_input_data[113 % IN_WIDTH];
                502 / IN_WIDTH: ping_storage_data_140 <= (fillup_transition == 1'b1) ? i_input_data[502 % IN_WIDTH] : ping_storage_data_140 ^ i_input_data[502 % IN_WIDTH];
                637 / IN_WIDTH: ping_storage_data_140 <= (fillup_transition == 1'b1) ? i_input_data[637 % IN_WIDTH] : ping_storage_data_140 ^ i_input_data[637 % IN_WIDTH];
                707 / IN_WIDTH: ping_storage_data_140 <= (fillup_transition == 1'b1) ? i_input_data[707 % IN_WIDTH] : ping_storage_data_140 ^ i_input_data[707 % IN_WIDTH];
                1088 / IN_WIDTH: ping_storage_data_140 <= (fillup_transition == 1'b1) ? i_input_data[1088 % IN_WIDTH] : ping_storage_data_140 ^ i_input_data[1088 % IN_WIDTH];
                default: ping_storage_data_140 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_140;
                endcase
            end else begin
                case (input_count)
                113 / IN_WIDTH: pong_storage_data_140 <= (fillup_transition == 1'b1) ? i_input_data[113 % IN_WIDTH] : pong_storage_data_140 ^ i_input_data[113 % IN_WIDTH];
                502 / IN_WIDTH: pong_storage_data_140 <= (fillup_transition == 1'b1) ? i_input_data[502 % IN_WIDTH] : pong_storage_data_140 ^ i_input_data[502 % IN_WIDTH];
                637 / IN_WIDTH: pong_storage_data_140 <= (fillup_transition == 1'b1) ? i_input_data[637 % IN_WIDTH] : pong_storage_data_140 ^ i_input_data[637 % IN_WIDTH];
                707 / IN_WIDTH: pong_storage_data_140 <= (fillup_transition == 1'b1) ? i_input_data[707 % IN_WIDTH] : pong_storage_data_140 ^ i_input_data[707 % IN_WIDTH];
                1088 / IN_WIDTH: pong_storage_data_140 <= (fillup_transition == 1'b1) ? i_input_data[1088 % IN_WIDTH] : pong_storage_data_140 ^ i_input_data[1088 % IN_WIDTH];
                default: pong_storage_data_140 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_140;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_140 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_140;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_140 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_140;
            end
        end
    end
end

logic ping_storage_data_141;
logic pong_storage_data_141;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_141 <= 1'b0;
        pong_storage_data_141 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                114 / IN_WIDTH: ping_storage_data_141 <= (fillup_transition == 1'b1) ? i_input_data[114 % IN_WIDTH] : ping_storage_data_141 ^ i_input_data[114 % IN_WIDTH];
                503 / IN_WIDTH: ping_storage_data_141 <= (fillup_transition == 1'b1) ? i_input_data[503 % IN_WIDTH] : ping_storage_data_141 ^ i_input_data[503 % IN_WIDTH];
                638 / IN_WIDTH: ping_storage_data_141 <= (fillup_transition == 1'b1) ? i_input_data[638 % IN_WIDTH] : ping_storage_data_141 ^ i_input_data[638 % IN_WIDTH];
                708 / IN_WIDTH: ping_storage_data_141 <= (fillup_transition == 1'b1) ? i_input_data[708 % IN_WIDTH] : ping_storage_data_141 ^ i_input_data[708 % IN_WIDTH];
                1089 / IN_WIDTH: ping_storage_data_141 <= (fillup_transition == 1'b1) ? i_input_data[1089 % IN_WIDTH] : ping_storage_data_141 ^ i_input_data[1089 % IN_WIDTH];
                default: ping_storage_data_141 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_141;
                endcase
            end else begin
                case (input_count)
                114 / IN_WIDTH: pong_storage_data_141 <= (fillup_transition == 1'b1) ? i_input_data[114 % IN_WIDTH] : pong_storage_data_141 ^ i_input_data[114 % IN_WIDTH];
                503 / IN_WIDTH: pong_storage_data_141 <= (fillup_transition == 1'b1) ? i_input_data[503 % IN_WIDTH] : pong_storage_data_141 ^ i_input_data[503 % IN_WIDTH];
                638 / IN_WIDTH: pong_storage_data_141 <= (fillup_transition == 1'b1) ? i_input_data[638 % IN_WIDTH] : pong_storage_data_141 ^ i_input_data[638 % IN_WIDTH];
                708 / IN_WIDTH: pong_storage_data_141 <= (fillup_transition == 1'b1) ? i_input_data[708 % IN_WIDTH] : pong_storage_data_141 ^ i_input_data[708 % IN_WIDTH];
                1089 / IN_WIDTH: pong_storage_data_141 <= (fillup_transition == 1'b1) ? i_input_data[1089 % IN_WIDTH] : pong_storage_data_141 ^ i_input_data[1089 % IN_WIDTH];
                default: pong_storage_data_141 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_141;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_141 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_141;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_141 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_141;
            end
        end
    end
end

logic ping_storage_data_142;
logic pong_storage_data_142;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_142 <= 1'b0;
        pong_storage_data_142 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                115 / IN_WIDTH: ping_storage_data_142 <= (fillup_transition == 1'b1) ? i_input_data[115 % IN_WIDTH] : ping_storage_data_142 ^ i_input_data[115 % IN_WIDTH];
                504 / IN_WIDTH: ping_storage_data_142 <= (fillup_transition == 1'b1) ? i_input_data[504 % IN_WIDTH] : ping_storage_data_142 ^ i_input_data[504 % IN_WIDTH];
                639 / IN_WIDTH: ping_storage_data_142 <= (fillup_transition == 1'b1) ? i_input_data[639 % IN_WIDTH] : ping_storage_data_142 ^ i_input_data[639 % IN_WIDTH];
                709 / IN_WIDTH: ping_storage_data_142 <= (fillup_transition == 1'b1) ? i_input_data[709 % IN_WIDTH] : ping_storage_data_142 ^ i_input_data[709 % IN_WIDTH];
                1090 / IN_WIDTH: ping_storage_data_142 <= (fillup_transition == 1'b1) ? i_input_data[1090 % IN_WIDTH] : ping_storage_data_142 ^ i_input_data[1090 % IN_WIDTH];
                default: ping_storage_data_142 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_142;
                endcase
            end else begin
                case (input_count)
                115 / IN_WIDTH: pong_storage_data_142 <= (fillup_transition == 1'b1) ? i_input_data[115 % IN_WIDTH] : pong_storage_data_142 ^ i_input_data[115 % IN_WIDTH];
                504 / IN_WIDTH: pong_storage_data_142 <= (fillup_transition == 1'b1) ? i_input_data[504 % IN_WIDTH] : pong_storage_data_142 ^ i_input_data[504 % IN_WIDTH];
                639 / IN_WIDTH: pong_storage_data_142 <= (fillup_transition == 1'b1) ? i_input_data[639 % IN_WIDTH] : pong_storage_data_142 ^ i_input_data[639 % IN_WIDTH];
                709 / IN_WIDTH: pong_storage_data_142 <= (fillup_transition == 1'b1) ? i_input_data[709 % IN_WIDTH] : pong_storage_data_142 ^ i_input_data[709 % IN_WIDTH];
                1090 / IN_WIDTH: pong_storage_data_142 <= (fillup_transition == 1'b1) ? i_input_data[1090 % IN_WIDTH] : pong_storage_data_142 ^ i_input_data[1090 % IN_WIDTH];
                default: pong_storage_data_142 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_142;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_142 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_142;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_142 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_142;
            end
        end
    end
end

logic ping_storage_data_143;
logic pong_storage_data_143;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_143 <= 1'b0;
        pong_storage_data_143 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                116 / IN_WIDTH: ping_storage_data_143 <= (fillup_transition == 1'b1) ? i_input_data[116 % IN_WIDTH] : ping_storage_data_143 ^ i_input_data[116 % IN_WIDTH];
                505 / IN_WIDTH: ping_storage_data_143 <= (fillup_transition == 1'b1) ? i_input_data[505 % IN_WIDTH] : ping_storage_data_143 ^ i_input_data[505 % IN_WIDTH];
                640 / IN_WIDTH: ping_storage_data_143 <= (fillup_transition == 1'b1) ? i_input_data[640 % IN_WIDTH] : ping_storage_data_143 ^ i_input_data[640 % IN_WIDTH];
                710 / IN_WIDTH: ping_storage_data_143 <= (fillup_transition == 1'b1) ? i_input_data[710 % IN_WIDTH] : ping_storage_data_143 ^ i_input_data[710 % IN_WIDTH];
                1091 / IN_WIDTH: ping_storage_data_143 <= (fillup_transition == 1'b1) ? i_input_data[1091 % IN_WIDTH] : ping_storage_data_143 ^ i_input_data[1091 % IN_WIDTH];
                default: ping_storage_data_143 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_143;
                endcase
            end else begin
                case (input_count)
                116 / IN_WIDTH: pong_storage_data_143 <= (fillup_transition == 1'b1) ? i_input_data[116 % IN_WIDTH] : pong_storage_data_143 ^ i_input_data[116 % IN_WIDTH];
                505 / IN_WIDTH: pong_storage_data_143 <= (fillup_transition == 1'b1) ? i_input_data[505 % IN_WIDTH] : pong_storage_data_143 ^ i_input_data[505 % IN_WIDTH];
                640 / IN_WIDTH: pong_storage_data_143 <= (fillup_transition == 1'b1) ? i_input_data[640 % IN_WIDTH] : pong_storage_data_143 ^ i_input_data[640 % IN_WIDTH];
                710 / IN_WIDTH: pong_storage_data_143 <= (fillup_transition == 1'b1) ? i_input_data[710 % IN_WIDTH] : pong_storage_data_143 ^ i_input_data[710 % IN_WIDTH];
                1091 / IN_WIDTH: pong_storage_data_143 <= (fillup_transition == 1'b1) ? i_input_data[1091 % IN_WIDTH] : pong_storage_data_143 ^ i_input_data[1091 % IN_WIDTH];
                default: pong_storage_data_143 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_143;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_143 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_143;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_143 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_143;
            end
        end
    end
end

logic ping_storage_data_144;
logic pong_storage_data_144;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_144 <= 1'b0;
        pong_storage_data_144 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                117 / IN_WIDTH: ping_storage_data_144 <= (fillup_transition == 1'b1) ? i_input_data[117 % IN_WIDTH] : ping_storage_data_144 ^ i_input_data[117 % IN_WIDTH];
                506 / IN_WIDTH: ping_storage_data_144 <= (fillup_transition == 1'b1) ? i_input_data[506 % IN_WIDTH] : ping_storage_data_144 ^ i_input_data[506 % IN_WIDTH];
                641 / IN_WIDTH: ping_storage_data_144 <= (fillup_transition == 1'b1) ? i_input_data[641 % IN_WIDTH] : ping_storage_data_144 ^ i_input_data[641 % IN_WIDTH];
                711 / IN_WIDTH: ping_storage_data_144 <= (fillup_transition == 1'b1) ? i_input_data[711 % IN_WIDTH] : ping_storage_data_144 ^ i_input_data[711 % IN_WIDTH];
                1092 / IN_WIDTH: ping_storage_data_144 <= (fillup_transition == 1'b1) ? i_input_data[1092 % IN_WIDTH] : ping_storage_data_144 ^ i_input_data[1092 % IN_WIDTH];
                default: ping_storage_data_144 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_144;
                endcase
            end else begin
                case (input_count)
                117 / IN_WIDTH: pong_storage_data_144 <= (fillup_transition == 1'b1) ? i_input_data[117 % IN_WIDTH] : pong_storage_data_144 ^ i_input_data[117 % IN_WIDTH];
                506 / IN_WIDTH: pong_storage_data_144 <= (fillup_transition == 1'b1) ? i_input_data[506 % IN_WIDTH] : pong_storage_data_144 ^ i_input_data[506 % IN_WIDTH];
                641 / IN_WIDTH: pong_storage_data_144 <= (fillup_transition == 1'b1) ? i_input_data[641 % IN_WIDTH] : pong_storage_data_144 ^ i_input_data[641 % IN_WIDTH];
                711 / IN_WIDTH: pong_storage_data_144 <= (fillup_transition == 1'b1) ? i_input_data[711 % IN_WIDTH] : pong_storage_data_144 ^ i_input_data[711 % IN_WIDTH];
                1092 / IN_WIDTH: pong_storage_data_144 <= (fillup_transition == 1'b1) ? i_input_data[1092 % IN_WIDTH] : pong_storage_data_144 ^ i_input_data[1092 % IN_WIDTH];
                default: pong_storage_data_144 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_144;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_144 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_144;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_144 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_144;
            end
        end
    end
end

logic ping_storage_data_145;
logic pong_storage_data_145;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_145 <= 1'b0;
        pong_storage_data_145 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                118 / IN_WIDTH: ping_storage_data_145 <= (fillup_transition == 1'b1) ? i_input_data[118 % IN_WIDTH] : ping_storage_data_145 ^ i_input_data[118 % IN_WIDTH];
                507 / IN_WIDTH: ping_storage_data_145 <= (fillup_transition == 1'b1) ? i_input_data[507 % IN_WIDTH] : ping_storage_data_145 ^ i_input_data[507 % IN_WIDTH];
                642 / IN_WIDTH: ping_storage_data_145 <= (fillup_transition == 1'b1) ? i_input_data[642 % IN_WIDTH] : ping_storage_data_145 ^ i_input_data[642 % IN_WIDTH];
                712 / IN_WIDTH: ping_storage_data_145 <= (fillup_transition == 1'b1) ? i_input_data[712 % IN_WIDTH] : ping_storage_data_145 ^ i_input_data[712 % IN_WIDTH];
                1093 / IN_WIDTH: ping_storage_data_145 <= (fillup_transition == 1'b1) ? i_input_data[1093 % IN_WIDTH] : ping_storage_data_145 ^ i_input_data[1093 % IN_WIDTH];
                default: ping_storage_data_145 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_145;
                endcase
            end else begin
                case (input_count)
                118 / IN_WIDTH: pong_storage_data_145 <= (fillup_transition == 1'b1) ? i_input_data[118 % IN_WIDTH] : pong_storage_data_145 ^ i_input_data[118 % IN_WIDTH];
                507 / IN_WIDTH: pong_storage_data_145 <= (fillup_transition == 1'b1) ? i_input_data[507 % IN_WIDTH] : pong_storage_data_145 ^ i_input_data[507 % IN_WIDTH];
                642 / IN_WIDTH: pong_storage_data_145 <= (fillup_transition == 1'b1) ? i_input_data[642 % IN_WIDTH] : pong_storage_data_145 ^ i_input_data[642 % IN_WIDTH];
                712 / IN_WIDTH: pong_storage_data_145 <= (fillup_transition == 1'b1) ? i_input_data[712 % IN_WIDTH] : pong_storage_data_145 ^ i_input_data[712 % IN_WIDTH];
                1093 / IN_WIDTH: pong_storage_data_145 <= (fillup_transition == 1'b1) ? i_input_data[1093 % IN_WIDTH] : pong_storage_data_145 ^ i_input_data[1093 % IN_WIDTH];
                default: pong_storage_data_145 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_145;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_145 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_145;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_145 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_145;
            end
        end
    end
end

logic ping_storage_data_146;
logic pong_storage_data_146;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_146 <= 1'b0;
        pong_storage_data_146 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                119 / IN_WIDTH: ping_storage_data_146 <= (fillup_transition == 1'b1) ? i_input_data[119 % IN_WIDTH] : ping_storage_data_146 ^ i_input_data[119 % IN_WIDTH];
                508 / IN_WIDTH: ping_storage_data_146 <= (fillup_transition == 1'b1) ? i_input_data[508 % IN_WIDTH] : ping_storage_data_146 ^ i_input_data[508 % IN_WIDTH];
                643 / IN_WIDTH: ping_storage_data_146 <= (fillup_transition == 1'b1) ? i_input_data[643 % IN_WIDTH] : ping_storage_data_146 ^ i_input_data[643 % IN_WIDTH];
                713 / IN_WIDTH: ping_storage_data_146 <= (fillup_transition == 1'b1) ? i_input_data[713 % IN_WIDTH] : ping_storage_data_146 ^ i_input_data[713 % IN_WIDTH];
                1094 / IN_WIDTH: ping_storage_data_146 <= (fillup_transition == 1'b1) ? i_input_data[1094 % IN_WIDTH] : ping_storage_data_146 ^ i_input_data[1094 % IN_WIDTH];
                default: ping_storage_data_146 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_146;
                endcase
            end else begin
                case (input_count)
                119 / IN_WIDTH: pong_storage_data_146 <= (fillup_transition == 1'b1) ? i_input_data[119 % IN_WIDTH] : pong_storage_data_146 ^ i_input_data[119 % IN_WIDTH];
                508 / IN_WIDTH: pong_storage_data_146 <= (fillup_transition == 1'b1) ? i_input_data[508 % IN_WIDTH] : pong_storage_data_146 ^ i_input_data[508 % IN_WIDTH];
                643 / IN_WIDTH: pong_storage_data_146 <= (fillup_transition == 1'b1) ? i_input_data[643 % IN_WIDTH] : pong_storage_data_146 ^ i_input_data[643 % IN_WIDTH];
                713 / IN_WIDTH: pong_storage_data_146 <= (fillup_transition == 1'b1) ? i_input_data[713 % IN_WIDTH] : pong_storage_data_146 ^ i_input_data[713 % IN_WIDTH];
                1094 / IN_WIDTH: pong_storage_data_146 <= (fillup_transition == 1'b1) ? i_input_data[1094 % IN_WIDTH] : pong_storage_data_146 ^ i_input_data[1094 % IN_WIDTH];
                default: pong_storage_data_146 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_146;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_146 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_146;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_146 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_146;
            end
        end
    end
end

logic ping_storage_data_147;
logic pong_storage_data_147;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_147 <= 1'b0;
        pong_storage_data_147 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                120 / IN_WIDTH: ping_storage_data_147 <= (fillup_transition == 1'b1) ? i_input_data[120 % IN_WIDTH] : ping_storage_data_147 ^ i_input_data[120 % IN_WIDTH];
                509 / IN_WIDTH: ping_storage_data_147 <= (fillup_transition == 1'b1) ? i_input_data[509 % IN_WIDTH] : ping_storage_data_147 ^ i_input_data[509 % IN_WIDTH];
                644 / IN_WIDTH: ping_storage_data_147 <= (fillup_transition == 1'b1) ? i_input_data[644 % IN_WIDTH] : ping_storage_data_147 ^ i_input_data[644 % IN_WIDTH];
                714 / IN_WIDTH: ping_storage_data_147 <= (fillup_transition == 1'b1) ? i_input_data[714 % IN_WIDTH] : ping_storage_data_147 ^ i_input_data[714 % IN_WIDTH];
                1095 / IN_WIDTH: ping_storage_data_147 <= (fillup_transition == 1'b1) ? i_input_data[1095 % IN_WIDTH] : ping_storage_data_147 ^ i_input_data[1095 % IN_WIDTH];
                default: ping_storage_data_147 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_147;
                endcase
            end else begin
                case (input_count)
                120 / IN_WIDTH: pong_storage_data_147 <= (fillup_transition == 1'b1) ? i_input_data[120 % IN_WIDTH] : pong_storage_data_147 ^ i_input_data[120 % IN_WIDTH];
                509 / IN_WIDTH: pong_storage_data_147 <= (fillup_transition == 1'b1) ? i_input_data[509 % IN_WIDTH] : pong_storage_data_147 ^ i_input_data[509 % IN_WIDTH];
                644 / IN_WIDTH: pong_storage_data_147 <= (fillup_transition == 1'b1) ? i_input_data[644 % IN_WIDTH] : pong_storage_data_147 ^ i_input_data[644 % IN_WIDTH];
                714 / IN_WIDTH: pong_storage_data_147 <= (fillup_transition == 1'b1) ? i_input_data[714 % IN_WIDTH] : pong_storage_data_147 ^ i_input_data[714 % IN_WIDTH];
                1095 / IN_WIDTH: pong_storage_data_147 <= (fillup_transition == 1'b1) ? i_input_data[1095 % IN_WIDTH] : pong_storage_data_147 ^ i_input_data[1095 % IN_WIDTH];
                default: pong_storage_data_147 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_147;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_147 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_147;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_147 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_147;
            end
        end
    end
end

logic ping_storage_data_148;
logic pong_storage_data_148;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_148 <= 1'b0;
        pong_storage_data_148 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                121 / IN_WIDTH: ping_storage_data_148 <= (fillup_transition == 1'b1) ? i_input_data[121 % IN_WIDTH] : ping_storage_data_148 ^ i_input_data[121 % IN_WIDTH];
                510 / IN_WIDTH: ping_storage_data_148 <= (fillup_transition == 1'b1) ? i_input_data[510 % IN_WIDTH] : ping_storage_data_148 ^ i_input_data[510 % IN_WIDTH];
                645 / IN_WIDTH: ping_storage_data_148 <= (fillup_transition == 1'b1) ? i_input_data[645 % IN_WIDTH] : ping_storage_data_148 ^ i_input_data[645 % IN_WIDTH];
                715 / IN_WIDTH: ping_storage_data_148 <= (fillup_transition == 1'b1) ? i_input_data[715 % IN_WIDTH] : ping_storage_data_148 ^ i_input_data[715 % IN_WIDTH];
                1096 / IN_WIDTH: ping_storage_data_148 <= (fillup_transition == 1'b1) ? i_input_data[1096 % IN_WIDTH] : ping_storage_data_148 ^ i_input_data[1096 % IN_WIDTH];
                default: ping_storage_data_148 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_148;
                endcase
            end else begin
                case (input_count)
                121 / IN_WIDTH: pong_storage_data_148 <= (fillup_transition == 1'b1) ? i_input_data[121 % IN_WIDTH] : pong_storage_data_148 ^ i_input_data[121 % IN_WIDTH];
                510 / IN_WIDTH: pong_storage_data_148 <= (fillup_transition == 1'b1) ? i_input_data[510 % IN_WIDTH] : pong_storage_data_148 ^ i_input_data[510 % IN_WIDTH];
                645 / IN_WIDTH: pong_storage_data_148 <= (fillup_transition == 1'b1) ? i_input_data[645 % IN_WIDTH] : pong_storage_data_148 ^ i_input_data[645 % IN_WIDTH];
                715 / IN_WIDTH: pong_storage_data_148 <= (fillup_transition == 1'b1) ? i_input_data[715 % IN_WIDTH] : pong_storage_data_148 ^ i_input_data[715 % IN_WIDTH];
                1096 / IN_WIDTH: pong_storage_data_148 <= (fillup_transition == 1'b1) ? i_input_data[1096 % IN_WIDTH] : pong_storage_data_148 ^ i_input_data[1096 % IN_WIDTH];
                default: pong_storage_data_148 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_148;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_148 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_148;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_148 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_148;
            end
        end
    end
end

logic ping_storage_data_149;
logic pong_storage_data_149;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_149 <= 1'b0;
        pong_storage_data_149 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                122 / IN_WIDTH: ping_storage_data_149 <= (fillup_transition == 1'b1) ? i_input_data[122 % IN_WIDTH] : ping_storage_data_149 ^ i_input_data[122 % IN_WIDTH];
                511 / IN_WIDTH: ping_storage_data_149 <= (fillup_transition == 1'b1) ? i_input_data[511 % IN_WIDTH] : ping_storage_data_149 ^ i_input_data[511 % IN_WIDTH];
                646 / IN_WIDTH: ping_storage_data_149 <= (fillup_transition == 1'b1) ? i_input_data[646 % IN_WIDTH] : ping_storage_data_149 ^ i_input_data[646 % IN_WIDTH];
                716 / IN_WIDTH: ping_storage_data_149 <= (fillup_transition == 1'b1) ? i_input_data[716 % IN_WIDTH] : ping_storage_data_149 ^ i_input_data[716 % IN_WIDTH];
                1097 / IN_WIDTH: ping_storage_data_149 <= (fillup_transition == 1'b1) ? i_input_data[1097 % IN_WIDTH] : ping_storage_data_149 ^ i_input_data[1097 % IN_WIDTH];
                default: ping_storage_data_149 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_149;
                endcase
            end else begin
                case (input_count)
                122 / IN_WIDTH: pong_storage_data_149 <= (fillup_transition == 1'b1) ? i_input_data[122 % IN_WIDTH] : pong_storage_data_149 ^ i_input_data[122 % IN_WIDTH];
                511 / IN_WIDTH: pong_storage_data_149 <= (fillup_transition == 1'b1) ? i_input_data[511 % IN_WIDTH] : pong_storage_data_149 ^ i_input_data[511 % IN_WIDTH];
                646 / IN_WIDTH: pong_storage_data_149 <= (fillup_transition == 1'b1) ? i_input_data[646 % IN_WIDTH] : pong_storage_data_149 ^ i_input_data[646 % IN_WIDTH];
                716 / IN_WIDTH: pong_storage_data_149 <= (fillup_transition == 1'b1) ? i_input_data[716 % IN_WIDTH] : pong_storage_data_149 ^ i_input_data[716 % IN_WIDTH];
                1097 / IN_WIDTH: pong_storage_data_149 <= (fillup_transition == 1'b1) ? i_input_data[1097 % IN_WIDTH] : pong_storage_data_149 ^ i_input_data[1097 % IN_WIDTH];
                default: pong_storage_data_149 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_149;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_149 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_149;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_149 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_149;
            end
        end
    end
end

logic ping_storage_data_150;
logic pong_storage_data_150;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_150 <= 1'b0;
        pong_storage_data_150 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                123 / IN_WIDTH: ping_storage_data_150 <= (fillup_transition == 1'b1) ? i_input_data[123 % IN_WIDTH] : ping_storage_data_150 ^ i_input_data[123 % IN_WIDTH];
                512 / IN_WIDTH: ping_storage_data_150 <= (fillup_transition == 1'b1) ? i_input_data[512 % IN_WIDTH] : ping_storage_data_150 ^ i_input_data[512 % IN_WIDTH];
                647 / IN_WIDTH: ping_storage_data_150 <= (fillup_transition == 1'b1) ? i_input_data[647 % IN_WIDTH] : ping_storage_data_150 ^ i_input_data[647 % IN_WIDTH];
                717 / IN_WIDTH: ping_storage_data_150 <= (fillup_transition == 1'b1) ? i_input_data[717 % IN_WIDTH] : ping_storage_data_150 ^ i_input_data[717 % IN_WIDTH];
                1098 / IN_WIDTH: ping_storage_data_150 <= (fillup_transition == 1'b1) ? i_input_data[1098 % IN_WIDTH] : ping_storage_data_150 ^ i_input_data[1098 % IN_WIDTH];
                default: ping_storage_data_150 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_150;
                endcase
            end else begin
                case (input_count)
                123 / IN_WIDTH: pong_storage_data_150 <= (fillup_transition == 1'b1) ? i_input_data[123 % IN_WIDTH] : pong_storage_data_150 ^ i_input_data[123 % IN_WIDTH];
                512 / IN_WIDTH: pong_storage_data_150 <= (fillup_transition == 1'b1) ? i_input_data[512 % IN_WIDTH] : pong_storage_data_150 ^ i_input_data[512 % IN_WIDTH];
                647 / IN_WIDTH: pong_storage_data_150 <= (fillup_transition == 1'b1) ? i_input_data[647 % IN_WIDTH] : pong_storage_data_150 ^ i_input_data[647 % IN_WIDTH];
                717 / IN_WIDTH: pong_storage_data_150 <= (fillup_transition == 1'b1) ? i_input_data[717 % IN_WIDTH] : pong_storage_data_150 ^ i_input_data[717 % IN_WIDTH];
                1098 / IN_WIDTH: pong_storage_data_150 <= (fillup_transition == 1'b1) ? i_input_data[1098 % IN_WIDTH] : pong_storage_data_150 ^ i_input_data[1098 % IN_WIDTH];
                default: pong_storage_data_150 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_150;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_150 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_150;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_150 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_150;
            end
        end
    end
end

logic ping_storage_data_151;
logic pong_storage_data_151;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_151 <= 1'b0;
        pong_storage_data_151 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                124 / IN_WIDTH: ping_storage_data_151 <= (fillup_transition == 1'b1) ? i_input_data[124 % IN_WIDTH] : ping_storage_data_151 ^ i_input_data[124 % IN_WIDTH];
                513 / IN_WIDTH: ping_storage_data_151 <= (fillup_transition == 1'b1) ? i_input_data[513 % IN_WIDTH] : ping_storage_data_151 ^ i_input_data[513 % IN_WIDTH];
                648 / IN_WIDTH: ping_storage_data_151 <= (fillup_transition == 1'b1) ? i_input_data[648 % IN_WIDTH] : ping_storage_data_151 ^ i_input_data[648 % IN_WIDTH];
                718 / IN_WIDTH: ping_storage_data_151 <= (fillup_transition == 1'b1) ? i_input_data[718 % IN_WIDTH] : ping_storage_data_151 ^ i_input_data[718 % IN_WIDTH];
                1099 / IN_WIDTH: ping_storage_data_151 <= (fillup_transition == 1'b1) ? i_input_data[1099 % IN_WIDTH] : ping_storage_data_151 ^ i_input_data[1099 % IN_WIDTH];
                default: ping_storage_data_151 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_151;
                endcase
            end else begin
                case (input_count)
                124 / IN_WIDTH: pong_storage_data_151 <= (fillup_transition == 1'b1) ? i_input_data[124 % IN_WIDTH] : pong_storage_data_151 ^ i_input_data[124 % IN_WIDTH];
                513 / IN_WIDTH: pong_storage_data_151 <= (fillup_transition == 1'b1) ? i_input_data[513 % IN_WIDTH] : pong_storage_data_151 ^ i_input_data[513 % IN_WIDTH];
                648 / IN_WIDTH: pong_storage_data_151 <= (fillup_transition == 1'b1) ? i_input_data[648 % IN_WIDTH] : pong_storage_data_151 ^ i_input_data[648 % IN_WIDTH];
                718 / IN_WIDTH: pong_storage_data_151 <= (fillup_transition == 1'b1) ? i_input_data[718 % IN_WIDTH] : pong_storage_data_151 ^ i_input_data[718 % IN_WIDTH];
                1099 / IN_WIDTH: pong_storage_data_151 <= (fillup_transition == 1'b1) ? i_input_data[1099 % IN_WIDTH] : pong_storage_data_151 ^ i_input_data[1099 % IN_WIDTH];
                default: pong_storage_data_151 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_151;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_151 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_151;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_151 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_151;
            end
        end
    end
end

logic ping_storage_data_152;
logic pong_storage_data_152;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_152 <= 1'b0;
        pong_storage_data_152 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                125 / IN_WIDTH: ping_storage_data_152 <= (fillup_transition == 1'b1) ? i_input_data[125 % IN_WIDTH] : ping_storage_data_152 ^ i_input_data[125 % IN_WIDTH];
                514 / IN_WIDTH: ping_storage_data_152 <= (fillup_transition == 1'b1) ? i_input_data[514 % IN_WIDTH] : ping_storage_data_152 ^ i_input_data[514 % IN_WIDTH];
                649 / IN_WIDTH: ping_storage_data_152 <= (fillup_transition == 1'b1) ? i_input_data[649 % IN_WIDTH] : ping_storage_data_152 ^ i_input_data[649 % IN_WIDTH];
                719 / IN_WIDTH: ping_storage_data_152 <= (fillup_transition == 1'b1) ? i_input_data[719 % IN_WIDTH] : ping_storage_data_152 ^ i_input_data[719 % IN_WIDTH];
                1100 / IN_WIDTH: ping_storage_data_152 <= (fillup_transition == 1'b1) ? i_input_data[1100 % IN_WIDTH] : ping_storage_data_152 ^ i_input_data[1100 % IN_WIDTH];
                default: ping_storage_data_152 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_152;
                endcase
            end else begin
                case (input_count)
                125 / IN_WIDTH: pong_storage_data_152 <= (fillup_transition == 1'b1) ? i_input_data[125 % IN_WIDTH] : pong_storage_data_152 ^ i_input_data[125 % IN_WIDTH];
                514 / IN_WIDTH: pong_storage_data_152 <= (fillup_transition == 1'b1) ? i_input_data[514 % IN_WIDTH] : pong_storage_data_152 ^ i_input_data[514 % IN_WIDTH];
                649 / IN_WIDTH: pong_storage_data_152 <= (fillup_transition == 1'b1) ? i_input_data[649 % IN_WIDTH] : pong_storage_data_152 ^ i_input_data[649 % IN_WIDTH];
                719 / IN_WIDTH: pong_storage_data_152 <= (fillup_transition == 1'b1) ? i_input_data[719 % IN_WIDTH] : pong_storage_data_152 ^ i_input_data[719 % IN_WIDTH];
                1100 / IN_WIDTH: pong_storage_data_152 <= (fillup_transition == 1'b1) ? i_input_data[1100 % IN_WIDTH] : pong_storage_data_152 ^ i_input_data[1100 % IN_WIDTH];
                default: pong_storage_data_152 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_152;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_152 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_152;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_152 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_152;
            end
        end
    end
end

logic ping_storage_data_153;
logic pong_storage_data_153;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_153 <= 1'b0;
        pong_storage_data_153 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                126 / IN_WIDTH: ping_storage_data_153 <= (fillup_transition == 1'b1) ? i_input_data[126 % IN_WIDTH] : ping_storage_data_153 ^ i_input_data[126 % IN_WIDTH];
                515 / IN_WIDTH: ping_storage_data_153 <= (fillup_transition == 1'b1) ? i_input_data[515 % IN_WIDTH] : ping_storage_data_153 ^ i_input_data[515 % IN_WIDTH];
                650 / IN_WIDTH: ping_storage_data_153 <= (fillup_transition == 1'b1) ? i_input_data[650 % IN_WIDTH] : ping_storage_data_153 ^ i_input_data[650 % IN_WIDTH];
                720 / IN_WIDTH: ping_storage_data_153 <= (fillup_transition == 1'b1) ? i_input_data[720 % IN_WIDTH] : ping_storage_data_153 ^ i_input_data[720 % IN_WIDTH];
                1101 / IN_WIDTH: ping_storage_data_153 <= (fillup_transition == 1'b1) ? i_input_data[1101 % IN_WIDTH] : ping_storage_data_153 ^ i_input_data[1101 % IN_WIDTH];
                default: ping_storage_data_153 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_153;
                endcase
            end else begin
                case (input_count)
                126 / IN_WIDTH: pong_storage_data_153 <= (fillup_transition == 1'b1) ? i_input_data[126 % IN_WIDTH] : pong_storage_data_153 ^ i_input_data[126 % IN_WIDTH];
                515 / IN_WIDTH: pong_storage_data_153 <= (fillup_transition == 1'b1) ? i_input_data[515 % IN_WIDTH] : pong_storage_data_153 ^ i_input_data[515 % IN_WIDTH];
                650 / IN_WIDTH: pong_storage_data_153 <= (fillup_transition == 1'b1) ? i_input_data[650 % IN_WIDTH] : pong_storage_data_153 ^ i_input_data[650 % IN_WIDTH];
                720 / IN_WIDTH: pong_storage_data_153 <= (fillup_transition == 1'b1) ? i_input_data[720 % IN_WIDTH] : pong_storage_data_153 ^ i_input_data[720 % IN_WIDTH];
                1101 / IN_WIDTH: pong_storage_data_153 <= (fillup_transition == 1'b1) ? i_input_data[1101 % IN_WIDTH] : pong_storage_data_153 ^ i_input_data[1101 % IN_WIDTH];
                default: pong_storage_data_153 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_153;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_153 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_153;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_153 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_153;
            end
        end
    end
end

logic ping_storage_data_154;
logic pong_storage_data_154;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_154 <= 1'b0;
        pong_storage_data_154 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                127 / IN_WIDTH: ping_storage_data_154 <= (fillup_transition == 1'b1) ? i_input_data[127 % IN_WIDTH] : ping_storage_data_154 ^ i_input_data[127 % IN_WIDTH];
                516 / IN_WIDTH: ping_storage_data_154 <= (fillup_transition == 1'b1) ? i_input_data[516 % IN_WIDTH] : ping_storage_data_154 ^ i_input_data[516 % IN_WIDTH];
                651 / IN_WIDTH: ping_storage_data_154 <= (fillup_transition == 1'b1) ? i_input_data[651 % IN_WIDTH] : ping_storage_data_154 ^ i_input_data[651 % IN_WIDTH];
                721 / IN_WIDTH: ping_storage_data_154 <= (fillup_transition == 1'b1) ? i_input_data[721 % IN_WIDTH] : ping_storage_data_154 ^ i_input_data[721 % IN_WIDTH];
                1102 / IN_WIDTH: ping_storage_data_154 <= (fillup_transition == 1'b1) ? i_input_data[1102 % IN_WIDTH] : ping_storage_data_154 ^ i_input_data[1102 % IN_WIDTH];
                default: ping_storage_data_154 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_154;
                endcase
            end else begin
                case (input_count)
                127 / IN_WIDTH: pong_storage_data_154 <= (fillup_transition == 1'b1) ? i_input_data[127 % IN_WIDTH] : pong_storage_data_154 ^ i_input_data[127 % IN_WIDTH];
                516 / IN_WIDTH: pong_storage_data_154 <= (fillup_transition == 1'b1) ? i_input_data[516 % IN_WIDTH] : pong_storage_data_154 ^ i_input_data[516 % IN_WIDTH];
                651 / IN_WIDTH: pong_storage_data_154 <= (fillup_transition == 1'b1) ? i_input_data[651 % IN_WIDTH] : pong_storage_data_154 ^ i_input_data[651 % IN_WIDTH];
                721 / IN_WIDTH: pong_storage_data_154 <= (fillup_transition == 1'b1) ? i_input_data[721 % IN_WIDTH] : pong_storage_data_154 ^ i_input_data[721 % IN_WIDTH];
                1102 / IN_WIDTH: pong_storage_data_154 <= (fillup_transition == 1'b1) ? i_input_data[1102 % IN_WIDTH] : pong_storage_data_154 ^ i_input_data[1102 % IN_WIDTH];
                default: pong_storage_data_154 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_154;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_154 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_154;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_154 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_154;
            end
        end
    end
end

logic ping_storage_data_155;
logic pong_storage_data_155;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_155 <= 1'b0;
        pong_storage_data_155 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                128 / IN_WIDTH: ping_storage_data_155 <= (fillup_transition == 1'b1) ? i_input_data[128 % IN_WIDTH] : ping_storage_data_155 ^ i_input_data[128 % IN_WIDTH];
                517 / IN_WIDTH: ping_storage_data_155 <= (fillup_transition == 1'b1) ? i_input_data[517 % IN_WIDTH] : ping_storage_data_155 ^ i_input_data[517 % IN_WIDTH];
                652 / IN_WIDTH: ping_storage_data_155 <= (fillup_transition == 1'b1) ? i_input_data[652 % IN_WIDTH] : ping_storage_data_155 ^ i_input_data[652 % IN_WIDTH];
                722 / IN_WIDTH: ping_storage_data_155 <= (fillup_transition == 1'b1) ? i_input_data[722 % IN_WIDTH] : ping_storage_data_155 ^ i_input_data[722 % IN_WIDTH];
                1103 / IN_WIDTH: ping_storage_data_155 <= (fillup_transition == 1'b1) ? i_input_data[1103 % IN_WIDTH] : ping_storage_data_155 ^ i_input_data[1103 % IN_WIDTH];
                default: ping_storage_data_155 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_155;
                endcase
            end else begin
                case (input_count)
                128 / IN_WIDTH: pong_storage_data_155 <= (fillup_transition == 1'b1) ? i_input_data[128 % IN_WIDTH] : pong_storage_data_155 ^ i_input_data[128 % IN_WIDTH];
                517 / IN_WIDTH: pong_storage_data_155 <= (fillup_transition == 1'b1) ? i_input_data[517 % IN_WIDTH] : pong_storage_data_155 ^ i_input_data[517 % IN_WIDTH];
                652 / IN_WIDTH: pong_storage_data_155 <= (fillup_transition == 1'b1) ? i_input_data[652 % IN_WIDTH] : pong_storage_data_155 ^ i_input_data[652 % IN_WIDTH];
                722 / IN_WIDTH: pong_storage_data_155 <= (fillup_transition == 1'b1) ? i_input_data[722 % IN_WIDTH] : pong_storage_data_155 ^ i_input_data[722 % IN_WIDTH];
                1103 / IN_WIDTH: pong_storage_data_155 <= (fillup_transition == 1'b1) ? i_input_data[1103 % IN_WIDTH] : pong_storage_data_155 ^ i_input_data[1103 % IN_WIDTH];
                default: pong_storage_data_155 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_155;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_155 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_155;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_155 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_155;
            end
        end
    end
end

logic ping_storage_data_156;
logic pong_storage_data_156;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_156 <= 1'b0;
        pong_storage_data_156 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                129 / IN_WIDTH: ping_storage_data_156 <= (fillup_transition == 1'b1) ? i_input_data[129 % IN_WIDTH] : ping_storage_data_156 ^ i_input_data[129 % IN_WIDTH];
                518 / IN_WIDTH: ping_storage_data_156 <= (fillup_transition == 1'b1) ? i_input_data[518 % IN_WIDTH] : ping_storage_data_156 ^ i_input_data[518 % IN_WIDTH];
                653 / IN_WIDTH: ping_storage_data_156 <= (fillup_transition == 1'b1) ? i_input_data[653 % IN_WIDTH] : ping_storage_data_156 ^ i_input_data[653 % IN_WIDTH];
                723 / IN_WIDTH: ping_storage_data_156 <= (fillup_transition == 1'b1) ? i_input_data[723 % IN_WIDTH] : ping_storage_data_156 ^ i_input_data[723 % IN_WIDTH];
                1104 / IN_WIDTH: ping_storage_data_156 <= (fillup_transition == 1'b1) ? i_input_data[1104 % IN_WIDTH] : ping_storage_data_156 ^ i_input_data[1104 % IN_WIDTH];
                default: ping_storage_data_156 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_156;
                endcase
            end else begin
                case (input_count)
                129 / IN_WIDTH: pong_storage_data_156 <= (fillup_transition == 1'b1) ? i_input_data[129 % IN_WIDTH] : pong_storage_data_156 ^ i_input_data[129 % IN_WIDTH];
                518 / IN_WIDTH: pong_storage_data_156 <= (fillup_transition == 1'b1) ? i_input_data[518 % IN_WIDTH] : pong_storage_data_156 ^ i_input_data[518 % IN_WIDTH];
                653 / IN_WIDTH: pong_storage_data_156 <= (fillup_transition == 1'b1) ? i_input_data[653 % IN_WIDTH] : pong_storage_data_156 ^ i_input_data[653 % IN_WIDTH];
                723 / IN_WIDTH: pong_storage_data_156 <= (fillup_transition == 1'b1) ? i_input_data[723 % IN_WIDTH] : pong_storage_data_156 ^ i_input_data[723 % IN_WIDTH];
                1104 / IN_WIDTH: pong_storage_data_156 <= (fillup_transition == 1'b1) ? i_input_data[1104 % IN_WIDTH] : pong_storage_data_156 ^ i_input_data[1104 % IN_WIDTH];
                default: pong_storage_data_156 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_156;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_156 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_156;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_156 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_156;
            end
        end
    end
end

logic ping_storage_data_157;
logic pong_storage_data_157;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_157 <= 1'b0;
        pong_storage_data_157 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                130 / IN_WIDTH: ping_storage_data_157 <= (fillup_transition == 1'b1) ? i_input_data[130 % IN_WIDTH] : ping_storage_data_157 ^ i_input_data[130 % IN_WIDTH];
                519 / IN_WIDTH: ping_storage_data_157 <= (fillup_transition == 1'b1) ? i_input_data[519 % IN_WIDTH] : ping_storage_data_157 ^ i_input_data[519 % IN_WIDTH];
                654 / IN_WIDTH: ping_storage_data_157 <= (fillup_transition == 1'b1) ? i_input_data[654 % IN_WIDTH] : ping_storage_data_157 ^ i_input_data[654 % IN_WIDTH];
                724 / IN_WIDTH: ping_storage_data_157 <= (fillup_transition == 1'b1) ? i_input_data[724 % IN_WIDTH] : ping_storage_data_157 ^ i_input_data[724 % IN_WIDTH];
                1105 / IN_WIDTH: ping_storage_data_157 <= (fillup_transition == 1'b1) ? i_input_data[1105 % IN_WIDTH] : ping_storage_data_157 ^ i_input_data[1105 % IN_WIDTH];
                default: ping_storage_data_157 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_157;
                endcase
            end else begin
                case (input_count)
                130 / IN_WIDTH: pong_storage_data_157 <= (fillup_transition == 1'b1) ? i_input_data[130 % IN_WIDTH] : pong_storage_data_157 ^ i_input_data[130 % IN_WIDTH];
                519 / IN_WIDTH: pong_storage_data_157 <= (fillup_transition == 1'b1) ? i_input_data[519 % IN_WIDTH] : pong_storage_data_157 ^ i_input_data[519 % IN_WIDTH];
                654 / IN_WIDTH: pong_storage_data_157 <= (fillup_transition == 1'b1) ? i_input_data[654 % IN_WIDTH] : pong_storage_data_157 ^ i_input_data[654 % IN_WIDTH];
                724 / IN_WIDTH: pong_storage_data_157 <= (fillup_transition == 1'b1) ? i_input_data[724 % IN_WIDTH] : pong_storage_data_157 ^ i_input_data[724 % IN_WIDTH];
                1105 / IN_WIDTH: pong_storage_data_157 <= (fillup_transition == 1'b1) ? i_input_data[1105 % IN_WIDTH] : pong_storage_data_157 ^ i_input_data[1105 % IN_WIDTH];
                default: pong_storage_data_157 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_157;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_157 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_157;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_157 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_157;
            end
        end
    end
end

logic ping_storage_data_158;
logic pong_storage_data_158;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_158 <= 1'b0;
        pong_storage_data_158 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                131 / IN_WIDTH: ping_storage_data_158 <= (fillup_transition == 1'b1) ? i_input_data[131 % IN_WIDTH] : ping_storage_data_158 ^ i_input_data[131 % IN_WIDTH];
                520 / IN_WIDTH: ping_storage_data_158 <= (fillup_transition == 1'b1) ? i_input_data[520 % IN_WIDTH] : ping_storage_data_158 ^ i_input_data[520 % IN_WIDTH];
                655 / IN_WIDTH: ping_storage_data_158 <= (fillup_transition == 1'b1) ? i_input_data[655 % IN_WIDTH] : ping_storage_data_158 ^ i_input_data[655 % IN_WIDTH];
                725 / IN_WIDTH: ping_storage_data_158 <= (fillup_transition == 1'b1) ? i_input_data[725 % IN_WIDTH] : ping_storage_data_158 ^ i_input_data[725 % IN_WIDTH];
                1106 / IN_WIDTH: ping_storage_data_158 <= (fillup_transition == 1'b1) ? i_input_data[1106 % IN_WIDTH] : ping_storage_data_158 ^ i_input_data[1106 % IN_WIDTH];
                default: ping_storage_data_158 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_158;
                endcase
            end else begin
                case (input_count)
                131 / IN_WIDTH: pong_storage_data_158 <= (fillup_transition == 1'b1) ? i_input_data[131 % IN_WIDTH] : pong_storage_data_158 ^ i_input_data[131 % IN_WIDTH];
                520 / IN_WIDTH: pong_storage_data_158 <= (fillup_transition == 1'b1) ? i_input_data[520 % IN_WIDTH] : pong_storage_data_158 ^ i_input_data[520 % IN_WIDTH];
                655 / IN_WIDTH: pong_storage_data_158 <= (fillup_transition == 1'b1) ? i_input_data[655 % IN_WIDTH] : pong_storage_data_158 ^ i_input_data[655 % IN_WIDTH];
                725 / IN_WIDTH: pong_storage_data_158 <= (fillup_transition == 1'b1) ? i_input_data[725 % IN_WIDTH] : pong_storage_data_158 ^ i_input_data[725 % IN_WIDTH];
                1106 / IN_WIDTH: pong_storage_data_158 <= (fillup_transition == 1'b1) ? i_input_data[1106 % IN_WIDTH] : pong_storage_data_158 ^ i_input_data[1106 % IN_WIDTH];
                default: pong_storage_data_158 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_158;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_158 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_158;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_158 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_158;
            end
        end
    end
end

logic ping_storage_data_159;
logic pong_storage_data_159;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_159 <= 1'b0;
        pong_storage_data_159 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                132 / IN_WIDTH: ping_storage_data_159 <= (fillup_transition == 1'b1) ? i_input_data[132 % IN_WIDTH] : ping_storage_data_159 ^ i_input_data[132 % IN_WIDTH];
                521 / IN_WIDTH: ping_storage_data_159 <= (fillup_transition == 1'b1) ? i_input_data[521 % IN_WIDTH] : ping_storage_data_159 ^ i_input_data[521 % IN_WIDTH];
                656 / IN_WIDTH: ping_storage_data_159 <= (fillup_transition == 1'b1) ? i_input_data[656 % IN_WIDTH] : ping_storage_data_159 ^ i_input_data[656 % IN_WIDTH];
                726 / IN_WIDTH: ping_storage_data_159 <= (fillup_transition == 1'b1) ? i_input_data[726 % IN_WIDTH] : ping_storage_data_159 ^ i_input_data[726 % IN_WIDTH];
                1107 / IN_WIDTH: ping_storage_data_159 <= (fillup_transition == 1'b1) ? i_input_data[1107 % IN_WIDTH] : ping_storage_data_159 ^ i_input_data[1107 % IN_WIDTH];
                default: ping_storage_data_159 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_159;
                endcase
            end else begin
                case (input_count)
                132 / IN_WIDTH: pong_storage_data_159 <= (fillup_transition == 1'b1) ? i_input_data[132 % IN_WIDTH] : pong_storage_data_159 ^ i_input_data[132 % IN_WIDTH];
                521 / IN_WIDTH: pong_storage_data_159 <= (fillup_transition == 1'b1) ? i_input_data[521 % IN_WIDTH] : pong_storage_data_159 ^ i_input_data[521 % IN_WIDTH];
                656 / IN_WIDTH: pong_storage_data_159 <= (fillup_transition == 1'b1) ? i_input_data[656 % IN_WIDTH] : pong_storage_data_159 ^ i_input_data[656 % IN_WIDTH];
                726 / IN_WIDTH: pong_storage_data_159 <= (fillup_transition == 1'b1) ? i_input_data[726 % IN_WIDTH] : pong_storage_data_159 ^ i_input_data[726 % IN_WIDTH];
                1107 / IN_WIDTH: pong_storage_data_159 <= (fillup_transition == 1'b1) ? i_input_data[1107 % IN_WIDTH] : pong_storage_data_159 ^ i_input_data[1107 % IN_WIDTH];
                default: pong_storage_data_159 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_159;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_159 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_159;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_159 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_159;
            end
        end
    end
end

logic ping_storage_data_160;
logic pong_storage_data_160;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_160 <= 1'b0;
        pong_storage_data_160 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                133 / IN_WIDTH: ping_storage_data_160 <= (fillup_transition == 1'b1) ? i_input_data[133 % IN_WIDTH] : ping_storage_data_160 ^ i_input_data[133 % IN_WIDTH];
                522 / IN_WIDTH: ping_storage_data_160 <= (fillup_transition == 1'b1) ? i_input_data[522 % IN_WIDTH] : ping_storage_data_160 ^ i_input_data[522 % IN_WIDTH];
                657 / IN_WIDTH: ping_storage_data_160 <= (fillup_transition == 1'b1) ? i_input_data[657 % IN_WIDTH] : ping_storage_data_160 ^ i_input_data[657 % IN_WIDTH];
                727 / IN_WIDTH: ping_storage_data_160 <= (fillup_transition == 1'b1) ? i_input_data[727 % IN_WIDTH] : ping_storage_data_160 ^ i_input_data[727 % IN_WIDTH];
                1108 / IN_WIDTH: ping_storage_data_160 <= (fillup_transition == 1'b1) ? i_input_data[1108 % IN_WIDTH] : ping_storage_data_160 ^ i_input_data[1108 % IN_WIDTH];
                default: ping_storage_data_160 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_160;
                endcase
            end else begin
                case (input_count)
                133 / IN_WIDTH: pong_storage_data_160 <= (fillup_transition == 1'b1) ? i_input_data[133 % IN_WIDTH] : pong_storage_data_160 ^ i_input_data[133 % IN_WIDTH];
                522 / IN_WIDTH: pong_storage_data_160 <= (fillup_transition == 1'b1) ? i_input_data[522 % IN_WIDTH] : pong_storage_data_160 ^ i_input_data[522 % IN_WIDTH];
                657 / IN_WIDTH: pong_storage_data_160 <= (fillup_transition == 1'b1) ? i_input_data[657 % IN_WIDTH] : pong_storage_data_160 ^ i_input_data[657 % IN_WIDTH];
                727 / IN_WIDTH: pong_storage_data_160 <= (fillup_transition == 1'b1) ? i_input_data[727 % IN_WIDTH] : pong_storage_data_160 ^ i_input_data[727 % IN_WIDTH];
                1108 / IN_WIDTH: pong_storage_data_160 <= (fillup_transition == 1'b1) ? i_input_data[1108 % IN_WIDTH] : pong_storage_data_160 ^ i_input_data[1108 % IN_WIDTH];
                default: pong_storage_data_160 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_160;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_160 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_160;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_160 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_160;
            end
        end
    end
end

logic ping_storage_data_161;
logic pong_storage_data_161;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_161 <= 1'b0;
        pong_storage_data_161 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                134 / IN_WIDTH: ping_storage_data_161 <= (fillup_transition == 1'b1) ? i_input_data[134 % IN_WIDTH] : ping_storage_data_161 ^ i_input_data[134 % IN_WIDTH];
                523 / IN_WIDTH: ping_storage_data_161 <= (fillup_transition == 1'b1) ? i_input_data[523 % IN_WIDTH] : ping_storage_data_161 ^ i_input_data[523 % IN_WIDTH];
                658 / IN_WIDTH: ping_storage_data_161 <= (fillup_transition == 1'b1) ? i_input_data[658 % IN_WIDTH] : ping_storage_data_161 ^ i_input_data[658 % IN_WIDTH];
                728 / IN_WIDTH: ping_storage_data_161 <= (fillup_transition == 1'b1) ? i_input_data[728 % IN_WIDTH] : ping_storage_data_161 ^ i_input_data[728 % IN_WIDTH];
                1109 / IN_WIDTH: ping_storage_data_161 <= (fillup_transition == 1'b1) ? i_input_data[1109 % IN_WIDTH] : ping_storage_data_161 ^ i_input_data[1109 % IN_WIDTH];
                default: ping_storage_data_161 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_161;
                endcase
            end else begin
                case (input_count)
                134 / IN_WIDTH: pong_storage_data_161 <= (fillup_transition == 1'b1) ? i_input_data[134 % IN_WIDTH] : pong_storage_data_161 ^ i_input_data[134 % IN_WIDTH];
                523 / IN_WIDTH: pong_storage_data_161 <= (fillup_transition == 1'b1) ? i_input_data[523 % IN_WIDTH] : pong_storage_data_161 ^ i_input_data[523 % IN_WIDTH];
                658 / IN_WIDTH: pong_storage_data_161 <= (fillup_transition == 1'b1) ? i_input_data[658 % IN_WIDTH] : pong_storage_data_161 ^ i_input_data[658 % IN_WIDTH];
                728 / IN_WIDTH: pong_storage_data_161 <= (fillup_transition == 1'b1) ? i_input_data[728 % IN_WIDTH] : pong_storage_data_161 ^ i_input_data[728 % IN_WIDTH];
                1109 / IN_WIDTH: pong_storage_data_161 <= (fillup_transition == 1'b1) ? i_input_data[1109 % IN_WIDTH] : pong_storage_data_161 ^ i_input_data[1109 % IN_WIDTH];
                default: pong_storage_data_161 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_161;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_161 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_161;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_161 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_161;
            end
        end
    end
end

logic ping_storage_data_162;
logic pong_storage_data_162;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_162 <= 1'b0;
        pong_storage_data_162 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                135 / IN_WIDTH: ping_storage_data_162 <= (fillup_transition == 1'b1) ? i_input_data[135 % IN_WIDTH] : ping_storage_data_162 ^ i_input_data[135 % IN_WIDTH];
                524 / IN_WIDTH: ping_storage_data_162 <= (fillup_transition == 1'b1) ? i_input_data[524 % IN_WIDTH] : ping_storage_data_162 ^ i_input_data[524 % IN_WIDTH];
                659 / IN_WIDTH: ping_storage_data_162 <= (fillup_transition == 1'b1) ? i_input_data[659 % IN_WIDTH] : ping_storage_data_162 ^ i_input_data[659 % IN_WIDTH];
                729 / IN_WIDTH: ping_storage_data_162 <= (fillup_transition == 1'b1) ? i_input_data[729 % IN_WIDTH] : ping_storage_data_162 ^ i_input_data[729 % IN_WIDTH];
                1110 / IN_WIDTH: ping_storage_data_162 <= (fillup_transition == 1'b1) ? i_input_data[1110 % IN_WIDTH] : ping_storage_data_162 ^ i_input_data[1110 % IN_WIDTH];
                default: ping_storage_data_162 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_162;
                endcase
            end else begin
                case (input_count)
                135 / IN_WIDTH: pong_storage_data_162 <= (fillup_transition == 1'b1) ? i_input_data[135 % IN_WIDTH] : pong_storage_data_162 ^ i_input_data[135 % IN_WIDTH];
                524 / IN_WIDTH: pong_storage_data_162 <= (fillup_transition == 1'b1) ? i_input_data[524 % IN_WIDTH] : pong_storage_data_162 ^ i_input_data[524 % IN_WIDTH];
                659 / IN_WIDTH: pong_storage_data_162 <= (fillup_transition == 1'b1) ? i_input_data[659 % IN_WIDTH] : pong_storage_data_162 ^ i_input_data[659 % IN_WIDTH];
                729 / IN_WIDTH: pong_storage_data_162 <= (fillup_transition == 1'b1) ? i_input_data[729 % IN_WIDTH] : pong_storage_data_162 ^ i_input_data[729 % IN_WIDTH];
                1110 / IN_WIDTH: pong_storage_data_162 <= (fillup_transition == 1'b1) ? i_input_data[1110 % IN_WIDTH] : pong_storage_data_162 ^ i_input_data[1110 % IN_WIDTH];
                default: pong_storage_data_162 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_162;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_162 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_162;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_162 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_162;
            end
        end
    end
end

logic ping_storage_data_163;
logic pong_storage_data_163;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_163 <= 1'b0;
        pong_storage_data_163 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                136 / IN_WIDTH: ping_storage_data_163 <= (fillup_transition == 1'b1) ? i_input_data[136 % IN_WIDTH] : ping_storage_data_163 ^ i_input_data[136 % IN_WIDTH];
                525 / IN_WIDTH: ping_storage_data_163 <= (fillup_transition == 1'b1) ? i_input_data[525 % IN_WIDTH] : ping_storage_data_163 ^ i_input_data[525 % IN_WIDTH];
                660 / IN_WIDTH: ping_storage_data_163 <= (fillup_transition == 1'b1) ? i_input_data[660 % IN_WIDTH] : ping_storage_data_163 ^ i_input_data[660 % IN_WIDTH];
                730 / IN_WIDTH: ping_storage_data_163 <= (fillup_transition == 1'b1) ? i_input_data[730 % IN_WIDTH] : ping_storage_data_163 ^ i_input_data[730 % IN_WIDTH];
                1111 / IN_WIDTH: ping_storage_data_163 <= (fillup_transition == 1'b1) ? i_input_data[1111 % IN_WIDTH] : ping_storage_data_163 ^ i_input_data[1111 % IN_WIDTH];
                default: ping_storage_data_163 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_163;
                endcase
            end else begin
                case (input_count)
                136 / IN_WIDTH: pong_storage_data_163 <= (fillup_transition == 1'b1) ? i_input_data[136 % IN_WIDTH] : pong_storage_data_163 ^ i_input_data[136 % IN_WIDTH];
                525 / IN_WIDTH: pong_storage_data_163 <= (fillup_transition == 1'b1) ? i_input_data[525 % IN_WIDTH] : pong_storage_data_163 ^ i_input_data[525 % IN_WIDTH];
                660 / IN_WIDTH: pong_storage_data_163 <= (fillup_transition == 1'b1) ? i_input_data[660 % IN_WIDTH] : pong_storage_data_163 ^ i_input_data[660 % IN_WIDTH];
                730 / IN_WIDTH: pong_storage_data_163 <= (fillup_transition == 1'b1) ? i_input_data[730 % IN_WIDTH] : pong_storage_data_163 ^ i_input_data[730 % IN_WIDTH];
                1111 / IN_WIDTH: pong_storage_data_163 <= (fillup_transition == 1'b1) ? i_input_data[1111 % IN_WIDTH] : pong_storage_data_163 ^ i_input_data[1111 % IN_WIDTH];
                default: pong_storage_data_163 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_163;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_163 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_163;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_163 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_163;
            end
        end
    end
end

logic ping_storage_data_164;
logic pong_storage_data_164;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_164 <= 1'b0;
        pong_storage_data_164 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                137 / IN_WIDTH: ping_storage_data_164 <= (fillup_transition == 1'b1) ? i_input_data[137 % IN_WIDTH] : ping_storage_data_164 ^ i_input_data[137 % IN_WIDTH];
                526 / IN_WIDTH: ping_storage_data_164 <= (fillup_transition == 1'b1) ? i_input_data[526 % IN_WIDTH] : ping_storage_data_164 ^ i_input_data[526 % IN_WIDTH];
                661 / IN_WIDTH: ping_storage_data_164 <= (fillup_transition == 1'b1) ? i_input_data[661 % IN_WIDTH] : ping_storage_data_164 ^ i_input_data[661 % IN_WIDTH];
                731 / IN_WIDTH: ping_storage_data_164 <= (fillup_transition == 1'b1) ? i_input_data[731 % IN_WIDTH] : ping_storage_data_164 ^ i_input_data[731 % IN_WIDTH];
                1112 / IN_WIDTH: ping_storage_data_164 <= (fillup_transition == 1'b1) ? i_input_data[1112 % IN_WIDTH] : ping_storage_data_164 ^ i_input_data[1112 % IN_WIDTH];
                default: ping_storage_data_164 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_164;
                endcase
            end else begin
                case (input_count)
                137 / IN_WIDTH: pong_storage_data_164 <= (fillup_transition == 1'b1) ? i_input_data[137 % IN_WIDTH] : pong_storage_data_164 ^ i_input_data[137 % IN_WIDTH];
                526 / IN_WIDTH: pong_storage_data_164 <= (fillup_transition == 1'b1) ? i_input_data[526 % IN_WIDTH] : pong_storage_data_164 ^ i_input_data[526 % IN_WIDTH];
                661 / IN_WIDTH: pong_storage_data_164 <= (fillup_transition == 1'b1) ? i_input_data[661 % IN_WIDTH] : pong_storage_data_164 ^ i_input_data[661 % IN_WIDTH];
                731 / IN_WIDTH: pong_storage_data_164 <= (fillup_transition == 1'b1) ? i_input_data[731 % IN_WIDTH] : pong_storage_data_164 ^ i_input_data[731 % IN_WIDTH];
                1112 / IN_WIDTH: pong_storage_data_164 <= (fillup_transition == 1'b1) ? i_input_data[1112 % IN_WIDTH] : pong_storage_data_164 ^ i_input_data[1112 % IN_WIDTH];
                default: pong_storage_data_164 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_164;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_164 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_164;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_164 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_164;
            end
        end
    end
end

logic ping_storage_data_165;
logic pong_storage_data_165;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_165 <= 1'b0;
        pong_storage_data_165 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                138 / IN_WIDTH: ping_storage_data_165 <= (fillup_transition == 1'b1) ? i_input_data[138 % IN_WIDTH] : ping_storage_data_165 ^ i_input_data[138 % IN_WIDTH];
                527 / IN_WIDTH: ping_storage_data_165 <= (fillup_transition == 1'b1) ? i_input_data[527 % IN_WIDTH] : ping_storage_data_165 ^ i_input_data[527 % IN_WIDTH];
                662 / IN_WIDTH: ping_storage_data_165 <= (fillup_transition == 1'b1) ? i_input_data[662 % IN_WIDTH] : ping_storage_data_165 ^ i_input_data[662 % IN_WIDTH];
                732 / IN_WIDTH: ping_storage_data_165 <= (fillup_transition == 1'b1) ? i_input_data[732 % IN_WIDTH] : ping_storage_data_165 ^ i_input_data[732 % IN_WIDTH];
                1113 / IN_WIDTH: ping_storage_data_165 <= (fillup_transition == 1'b1) ? i_input_data[1113 % IN_WIDTH] : ping_storage_data_165 ^ i_input_data[1113 % IN_WIDTH];
                default: ping_storage_data_165 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_165;
                endcase
            end else begin
                case (input_count)
                138 / IN_WIDTH: pong_storage_data_165 <= (fillup_transition == 1'b1) ? i_input_data[138 % IN_WIDTH] : pong_storage_data_165 ^ i_input_data[138 % IN_WIDTH];
                527 / IN_WIDTH: pong_storage_data_165 <= (fillup_transition == 1'b1) ? i_input_data[527 % IN_WIDTH] : pong_storage_data_165 ^ i_input_data[527 % IN_WIDTH];
                662 / IN_WIDTH: pong_storage_data_165 <= (fillup_transition == 1'b1) ? i_input_data[662 % IN_WIDTH] : pong_storage_data_165 ^ i_input_data[662 % IN_WIDTH];
                732 / IN_WIDTH: pong_storage_data_165 <= (fillup_transition == 1'b1) ? i_input_data[732 % IN_WIDTH] : pong_storage_data_165 ^ i_input_data[732 % IN_WIDTH];
                1113 / IN_WIDTH: pong_storage_data_165 <= (fillup_transition == 1'b1) ? i_input_data[1113 % IN_WIDTH] : pong_storage_data_165 ^ i_input_data[1113 % IN_WIDTH];
                default: pong_storage_data_165 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_165;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_165 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_165;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_165 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_165;
            end
        end
    end
end

logic ping_storage_data_166;
logic pong_storage_data_166;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_166 <= 1'b0;
        pong_storage_data_166 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                139 / IN_WIDTH: ping_storage_data_166 <= (fillup_transition == 1'b1) ? i_input_data[139 % IN_WIDTH] : ping_storage_data_166 ^ i_input_data[139 % IN_WIDTH];
                528 / IN_WIDTH: ping_storage_data_166 <= (fillup_transition == 1'b1) ? i_input_data[528 % IN_WIDTH] : ping_storage_data_166 ^ i_input_data[528 % IN_WIDTH];
                663 / IN_WIDTH: ping_storage_data_166 <= (fillup_transition == 1'b1) ? i_input_data[663 % IN_WIDTH] : ping_storage_data_166 ^ i_input_data[663 % IN_WIDTH];
                733 / IN_WIDTH: ping_storage_data_166 <= (fillup_transition == 1'b1) ? i_input_data[733 % IN_WIDTH] : ping_storage_data_166 ^ i_input_data[733 % IN_WIDTH];
                1114 / IN_WIDTH: ping_storage_data_166 <= (fillup_transition == 1'b1) ? i_input_data[1114 % IN_WIDTH] : ping_storage_data_166 ^ i_input_data[1114 % IN_WIDTH];
                default: ping_storage_data_166 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_166;
                endcase
            end else begin
                case (input_count)
                139 / IN_WIDTH: pong_storage_data_166 <= (fillup_transition == 1'b1) ? i_input_data[139 % IN_WIDTH] : pong_storage_data_166 ^ i_input_data[139 % IN_WIDTH];
                528 / IN_WIDTH: pong_storage_data_166 <= (fillup_transition == 1'b1) ? i_input_data[528 % IN_WIDTH] : pong_storage_data_166 ^ i_input_data[528 % IN_WIDTH];
                663 / IN_WIDTH: pong_storage_data_166 <= (fillup_transition == 1'b1) ? i_input_data[663 % IN_WIDTH] : pong_storage_data_166 ^ i_input_data[663 % IN_WIDTH];
                733 / IN_WIDTH: pong_storage_data_166 <= (fillup_transition == 1'b1) ? i_input_data[733 % IN_WIDTH] : pong_storage_data_166 ^ i_input_data[733 % IN_WIDTH];
                1114 / IN_WIDTH: pong_storage_data_166 <= (fillup_transition == 1'b1) ? i_input_data[1114 % IN_WIDTH] : pong_storage_data_166 ^ i_input_data[1114 % IN_WIDTH];
                default: pong_storage_data_166 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_166;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_166 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_166;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_166 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_166;
            end
        end
    end
end

logic ping_storage_data_167;
logic pong_storage_data_167;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_167 <= 1'b0;
        pong_storage_data_167 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                140 / IN_WIDTH: ping_storage_data_167 <= (fillup_transition == 1'b1) ? i_input_data[140 % IN_WIDTH] : ping_storage_data_167 ^ i_input_data[140 % IN_WIDTH];
                529 / IN_WIDTH: ping_storage_data_167 <= (fillup_transition == 1'b1) ? i_input_data[529 % IN_WIDTH] : ping_storage_data_167 ^ i_input_data[529 % IN_WIDTH];
                664 / IN_WIDTH: ping_storage_data_167 <= (fillup_transition == 1'b1) ? i_input_data[664 % IN_WIDTH] : ping_storage_data_167 ^ i_input_data[664 % IN_WIDTH];
                734 / IN_WIDTH: ping_storage_data_167 <= (fillup_transition == 1'b1) ? i_input_data[734 % IN_WIDTH] : ping_storage_data_167 ^ i_input_data[734 % IN_WIDTH];
                1115 / IN_WIDTH: ping_storage_data_167 <= (fillup_transition == 1'b1) ? i_input_data[1115 % IN_WIDTH] : ping_storage_data_167 ^ i_input_data[1115 % IN_WIDTH];
                default: ping_storage_data_167 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_167;
                endcase
            end else begin
                case (input_count)
                140 / IN_WIDTH: pong_storage_data_167 <= (fillup_transition == 1'b1) ? i_input_data[140 % IN_WIDTH] : pong_storage_data_167 ^ i_input_data[140 % IN_WIDTH];
                529 / IN_WIDTH: pong_storage_data_167 <= (fillup_transition == 1'b1) ? i_input_data[529 % IN_WIDTH] : pong_storage_data_167 ^ i_input_data[529 % IN_WIDTH];
                664 / IN_WIDTH: pong_storage_data_167 <= (fillup_transition == 1'b1) ? i_input_data[664 % IN_WIDTH] : pong_storage_data_167 ^ i_input_data[664 % IN_WIDTH];
                734 / IN_WIDTH: pong_storage_data_167 <= (fillup_transition == 1'b1) ? i_input_data[734 % IN_WIDTH] : pong_storage_data_167 ^ i_input_data[734 % IN_WIDTH];
                1115 / IN_WIDTH: pong_storage_data_167 <= (fillup_transition == 1'b1) ? i_input_data[1115 % IN_WIDTH] : pong_storage_data_167 ^ i_input_data[1115 % IN_WIDTH];
                default: pong_storage_data_167 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_167;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_167 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_167;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_167 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_167;
            end
        end
    end
end

logic ping_storage_data_168;
logic pong_storage_data_168;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_168 <= 1'b0;
        pong_storage_data_168 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                141 / IN_WIDTH: ping_storage_data_168 <= (fillup_transition == 1'b1) ? i_input_data[141 % IN_WIDTH] : ping_storage_data_168 ^ i_input_data[141 % IN_WIDTH];
                530 / IN_WIDTH: ping_storage_data_168 <= (fillup_transition == 1'b1) ? i_input_data[530 % IN_WIDTH] : ping_storage_data_168 ^ i_input_data[530 % IN_WIDTH];
                665 / IN_WIDTH: ping_storage_data_168 <= (fillup_transition == 1'b1) ? i_input_data[665 % IN_WIDTH] : ping_storage_data_168 ^ i_input_data[665 % IN_WIDTH];
                735 / IN_WIDTH: ping_storage_data_168 <= (fillup_transition == 1'b1) ? i_input_data[735 % IN_WIDTH] : ping_storage_data_168 ^ i_input_data[735 % IN_WIDTH];
                1116 / IN_WIDTH: ping_storage_data_168 <= (fillup_transition == 1'b1) ? i_input_data[1116 % IN_WIDTH] : ping_storage_data_168 ^ i_input_data[1116 % IN_WIDTH];
                default: ping_storage_data_168 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_168;
                endcase
            end else begin
                case (input_count)
                141 / IN_WIDTH: pong_storage_data_168 <= (fillup_transition == 1'b1) ? i_input_data[141 % IN_WIDTH] : pong_storage_data_168 ^ i_input_data[141 % IN_WIDTH];
                530 / IN_WIDTH: pong_storage_data_168 <= (fillup_transition == 1'b1) ? i_input_data[530 % IN_WIDTH] : pong_storage_data_168 ^ i_input_data[530 % IN_WIDTH];
                665 / IN_WIDTH: pong_storage_data_168 <= (fillup_transition == 1'b1) ? i_input_data[665 % IN_WIDTH] : pong_storage_data_168 ^ i_input_data[665 % IN_WIDTH];
                735 / IN_WIDTH: pong_storage_data_168 <= (fillup_transition == 1'b1) ? i_input_data[735 % IN_WIDTH] : pong_storage_data_168 ^ i_input_data[735 % IN_WIDTH];
                1116 / IN_WIDTH: pong_storage_data_168 <= (fillup_transition == 1'b1) ? i_input_data[1116 % IN_WIDTH] : pong_storage_data_168 ^ i_input_data[1116 % IN_WIDTH];
                default: pong_storage_data_168 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_168;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_168 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_168;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_168 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_168;
            end
        end
    end
end

logic ping_storage_data_169;
logic pong_storage_data_169;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_169 <= 1'b0;
        pong_storage_data_169 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                142 / IN_WIDTH: ping_storage_data_169 <= (fillup_transition == 1'b1) ? i_input_data[142 % IN_WIDTH] : ping_storage_data_169 ^ i_input_data[142 % IN_WIDTH];
                531 / IN_WIDTH: ping_storage_data_169 <= (fillup_transition == 1'b1) ? i_input_data[531 % IN_WIDTH] : ping_storage_data_169 ^ i_input_data[531 % IN_WIDTH];
                666 / IN_WIDTH: ping_storage_data_169 <= (fillup_transition == 1'b1) ? i_input_data[666 % IN_WIDTH] : ping_storage_data_169 ^ i_input_data[666 % IN_WIDTH];
                736 / IN_WIDTH: ping_storage_data_169 <= (fillup_transition == 1'b1) ? i_input_data[736 % IN_WIDTH] : ping_storage_data_169 ^ i_input_data[736 % IN_WIDTH];
                1117 / IN_WIDTH: ping_storage_data_169 <= (fillup_transition == 1'b1) ? i_input_data[1117 % IN_WIDTH] : ping_storage_data_169 ^ i_input_data[1117 % IN_WIDTH];
                default: ping_storage_data_169 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_169;
                endcase
            end else begin
                case (input_count)
                142 / IN_WIDTH: pong_storage_data_169 <= (fillup_transition == 1'b1) ? i_input_data[142 % IN_WIDTH] : pong_storage_data_169 ^ i_input_data[142 % IN_WIDTH];
                531 / IN_WIDTH: pong_storage_data_169 <= (fillup_transition == 1'b1) ? i_input_data[531 % IN_WIDTH] : pong_storage_data_169 ^ i_input_data[531 % IN_WIDTH];
                666 / IN_WIDTH: pong_storage_data_169 <= (fillup_transition == 1'b1) ? i_input_data[666 % IN_WIDTH] : pong_storage_data_169 ^ i_input_data[666 % IN_WIDTH];
                736 / IN_WIDTH: pong_storage_data_169 <= (fillup_transition == 1'b1) ? i_input_data[736 % IN_WIDTH] : pong_storage_data_169 ^ i_input_data[736 % IN_WIDTH];
                1117 / IN_WIDTH: pong_storage_data_169 <= (fillup_transition == 1'b1) ? i_input_data[1117 % IN_WIDTH] : pong_storage_data_169 ^ i_input_data[1117 % IN_WIDTH];
                default: pong_storage_data_169 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_169;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_169 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_169;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_169 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_169;
            end
        end
    end
end

logic ping_storage_data_170;
logic pong_storage_data_170;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_170 <= 1'b0;
        pong_storage_data_170 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                143 / IN_WIDTH: ping_storage_data_170 <= (fillup_transition == 1'b1) ? i_input_data[143 % IN_WIDTH] : ping_storage_data_170 ^ i_input_data[143 % IN_WIDTH];
                532 / IN_WIDTH: ping_storage_data_170 <= (fillup_transition == 1'b1) ? i_input_data[532 % IN_WIDTH] : ping_storage_data_170 ^ i_input_data[532 % IN_WIDTH];
                667 / IN_WIDTH: ping_storage_data_170 <= (fillup_transition == 1'b1) ? i_input_data[667 % IN_WIDTH] : ping_storage_data_170 ^ i_input_data[667 % IN_WIDTH];
                737 / IN_WIDTH: ping_storage_data_170 <= (fillup_transition == 1'b1) ? i_input_data[737 % IN_WIDTH] : ping_storage_data_170 ^ i_input_data[737 % IN_WIDTH];
                1118 / IN_WIDTH: ping_storage_data_170 <= (fillup_transition == 1'b1) ? i_input_data[1118 % IN_WIDTH] : ping_storage_data_170 ^ i_input_data[1118 % IN_WIDTH];
                default: ping_storage_data_170 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_170;
                endcase
            end else begin
                case (input_count)
                143 / IN_WIDTH: pong_storage_data_170 <= (fillup_transition == 1'b1) ? i_input_data[143 % IN_WIDTH] : pong_storage_data_170 ^ i_input_data[143 % IN_WIDTH];
                532 / IN_WIDTH: pong_storage_data_170 <= (fillup_transition == 1'b1) ? i_input_data[532 % IN_WIDTH] : pong_storage_data_170 ^ i_input_data[532 % IN_WIDTH];
                667 / IN_WIDTH: pong_storage_data_170 <= (fillup_transition == 1'b1) ? i_input_data[667 % IN_WIDTH] : pong_storage_data_170 ^ i_input_data[667 % IN_WIDTH];
                737 / IN_WIDTH: pong_storage_data_170 <= (fillup_transition == 1'b1) ? i_input_data[737 % IN_WIDTH] : pong_storage_data_170 ^ i_input_data[737 % IN_WIDTH];
                1118 / IN_WIDTH: pong_storage_data_170 <= (fillup_transition == 1'b1) ? i_input_data[1118 % IN_WIDTH] : pong_storage_data_170 ^ i_input_data[1118 % IN_WIDTH];
                default: pong_storage_data_170 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_170;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_170 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_170;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_170 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_170;
            end
        end
    end
end

logic ping_storage_data_171;
logic pong_storage_data_171;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_171 <= 1'b0;
        pong_storage_data_171 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                144 / IN_WIDTH: ping_storage_data_171 <= (fillup_transition == 1'b1) ? i_input_data[144 % IN_WIDTH] : ping_storage_data_171 ^ i_input_data[144 % IN_WIDTH];
                533 / IN_WIDTH: ping_storage_data_171 <= (fillup_transition == 1'b1) ? i_input_data[533 % IN_WIDTH] : ping_storage_data_171 ^ i_input_data[533 % IN_WIDTH];
                668 / IN_WIDTH: ping_storage_data_171 <= (fillup_transition == 1'b1) ? i_input_data[668 % IN_WIDTH] : ping_storage_data_171 ^ i_input_data[668 % IN_WIDTH];
                738 / IN_WIDTH: ping_storage_data_171 <= (fillup_transition == 1'b1) ? i_input_data[738 % IN_WIDTH] : ping_storage_data_171 ^ i_input_data[738 % IN_WIDTH];
                1119 / IN_WIDTH: ping_storage_data_171 <= (fillup_transition == 1'b1) ? i_input_data[1119 % IN_WIDTH] : ping_storage_data_171 ^ i_input_data[1119 % IN_WIDTH];
                default: ping_storage_data_171 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_171;
                endcase
            end else begin
                case (input_count)
                144 / IN_WIDTH: pong_storage_data_171 <= (fillup_transition == 1'b1) ? i_input_data[144 % IN_WIDTH] : pong_storage_data_171 ^ i_input_data[144 % IN_WIDTH];
                533 / IN_WIDTH: pong_storage_data_171 <= (fillup_transition == 1'b1) ? i_input_data[533 % IN_WIDTH] : pong_storage_data_171 ^ i_input_data[533 % IN_WIDTH];
                668 / IN_WIDTH: pong_storage_data_171 <= (fillup_transition == 1'b1) ? i_input_data[668 % IN_WIDTH] : pong_storage_data_171 ^ i_input_data[668 % IN_WIDTH];
                738 / IN_WIDTH: pong_storage_data_171 <= (fillup_transition == 1'b1) ? i_input_data[738 % IN_WIDTH] : pong_storage_data_171 ^ i_input_data[738 % IN_WIDTH];
                1119 / IN_WIDTH: pong_storage_data_171 <= (fillup_transition == 1'b1) ? i_input_data[1119 % IN_WIDTH] : pong_storage_data_171 ^ i_input_data[1119 % IN_WIDTH];
                default: pong_storage_data_171 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_171;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_171 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_171;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_171 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_171;
            end
        end
    end
end

logic ping_storage_data_172;
logic pong_storage_data_172;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_172 <= 1'b0;
        pong_storage_data_172 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                145 / IN_WIDTH: ping_storage_data_172 <= (fillup_transition == 1'b1) ? i_input_data[145 % IN_WIDTH] : ping_storage_data_172 ^ i_input_data[145 % IN_WIDTH];
                534 / IN_WIDTH: ping_storage_data_172 <= (fillup_transition == 1'b1) ? i_input_data[534 % IN_WIDTH] : ping_storage_data_172 ^ i_input_data[534 % IN_WIDTH];
                669 / IN_WIDTH: ping_storage_data_172 <= (fillup_transition == 1'b1) ? i_input_data[669 % IN_WIDTH] : ping_storage_data_172 ^ i_input_data[669 % IN_WIDTH];
                739 / IN_WIDTH: ping_storage_data_172 <= (fillup_transition == 1'b1) ? i_input_data[739 % IN_WIDTH] : ping_storage_data_172 ^ i_input_data[739 % IN_WIDTH];
                1120 / IN_WIDTH: ping_storage_data_172 <= (fillup_transition == 1'b1) ? i_input_data[1120 % IN_WIDTH] : ping_storage_data_172 ^ i_input_data[1120 % IN_WIDTH];
                default: ping_storage_data_172 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_172;
                endcase
            end else begin
                case (input_count)
                145 / IN_WIDTH: pong_storage_data_172 <= (fillup_transition == 1'b1) ? i_input_data[145 % IN_WIDTH] : pong_storage_data_172 ^ i_input_data[145 % IN_WIDTH];
                534 / IN_WIDTH: pong_storage_data_172 <= (fillup_transition == 1'b1) ? i_input_data[534 % IN_WIDTH] : pong_storage_data_172 ^ i_input_data[534 % IN_WIDTH];
                669 / IN_WIDTH: pong_storage_data_172 <= (fillup_transition == 1'b1) ? i_input_data[669 % IN_WIDTH] : pong_storage_data_172 ^ i_input_data[669 % IN_WIDTH];
                739 / IN_WIDTH: pong_storage_data_172 <= (fillup_transition == 1'b1) ? i_input_data[739 % IN_WIDTH] : pong_storage_data_172 ^ i_input_data[739 % IN_WIDTH];
                1120 / IN_WIDTH: pong_storage_data_172 <= (fillup_transition == 1'b1) ? i_input_data[1120 % IN_WIDTH] : pong_storage_data_172 ^ i_input_data[1120 % IN_WIDTH];
                default: pong_storage_data_172 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_172;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_172 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_172;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_172 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_172;
            end
        end
    end
end

logic ping_storage_data_173;
logic pong_storage_data_173;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_173 <= 1'b0;
        pong_storage_data_173 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                146 / IN_WIDTH: ping_storage_data_173 <= (fillup_transition == 1'b1) ? i_input_data[146 % IN_WIDTH] : ping_storage_data_173 ^ i_input_data[146 % IN_WIDTH];
                535 / IN_WIDTH: ping_storage_data_173 <= (fillup_transition == 1'b1) ? i_input_data[535 % IN_WIDTH] : ping_storage_data_173 ^ i_input_data[535 % IN_WIDTH];
                670 / IN_WIDTH: ping_storage_data_173 <= (fillup_transition == 1'b1) ? i_input_data[670 % IN_WIDTH] : ping_storage_data_173 ^ i_input_data[670 % IN_WIDTH];
                740 / IN_WIDTH: ping_storage_data_173 <= (fillup_transition == 1'b1) ? i_input_data[740 % IN_WIDTH] : ping_storage_data_173 ^ i_input_data[740 % IN_WIDTH];
                1121 / IN_WIDTH: ping_storage_data_173 <= (fillup_transition == 1'b1) ? i_input_data[1121 % IN_WIDTH] : ping_storage_data_173 ^ i_input_data[1121 % IN_WIDTH];
                default: ping_storage_data_173 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_173;
                endcase
            end else begin
                case (input_count)
                146 / IN_WIDTH: pong_storage_data_173 <= (fillup_transition == 1'b1) ? i_input_data[146 % IN_WIDTH] : pong_storage_data_173 ^ i_input_data[146 % IN_WIDTH];
                535 / IN_WIDTH: pong_storage_data_173 <= (fillup_transition == 1'b1) ? i_input_data[535 % IN_WIDTH] : pong_storage_data_173 ^ i_input_data[535 % IN_WIDTH];
                670 / IN_WIDTH: pong_storage_data_173 <= (fillup_transition == 1'b1) ? i_input_data[670 % IN_WIDTH] : pong_storage_data_173 ^ i_input_data[670 % IN_WIDTH];
                740 / IN_WIDTH: pong_storage_data_173 <= (fillup_transition == 1'b1) ? i_input_data[740 % IN_WIDTH] : pong_storage_data_173 ^ i_input_data[740 % IN_WIDTH];
                1121 / IN_WIDTH: pong_storage_data_173 <= (fillup_transition == 1'b1) ? i_input_data[1121 % IN_WIDTH] : pong_storage_data_173 ^ i_input_data[1121 % IN_WIDTH];
                default: pong_storage_data_173 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_173;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_173 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_173;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_173 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_173;
            end
        end
    end
end

logic ping_storage_data_174;
logic pong_storage_data_174;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_174 <= 1'b0;
        pong_storage_data_174 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                147 / IN_WIDTH: ping_storage_data_174 <= (fillup_transition == 1'b1) ? i_input_data[147 % IN_WIDTH] : ping_storage_data_174 ^ i_input_data[147 % IN_WIDTH];
                536 / IN_WIDTH: ping_storage_data_174 <= (fillup_transition == 1'b1) ? i_input_data[536 % IN_WIDTH] : ping_storage_data_174 ^ i_input_data[536 % IN_WIDTH];
                671 / IN_WIDTH: ping_storage_data_174 <= (fillup_transition == 1'b1) ? i_input_data[671 % IN_WIDTH] : ping_storage_data_174 ^ i_input_data[671 % IN_WIDTH];
                741 / IN_WIDTH: ping_storage_data_174 <= (fillup_transition == 1'b1) ? i_input_data[741 % IN_WIDTH] : ping_storage_data_174 ^ i_input_data[741 % IN_WIDTH];
                1122 / IN_WIDTH: ping_storage_data_174 <= (fillup_transition == 1'b1) ? i_input_data[1122 % IN_WIDTH] : ping_storage_data_174 ^ i_input_data[1122 % IN_WIDTH];
                default: ping_storage_data_174 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_174;
                endcase
            end else begin
                case (input_count)
                147 / IN_WIDTH: pong_storage_data_174 <= (fillup_transition == 1'b1) ? i_input_data[147 % IN_WIDTH] : pong_storage_data_174 ^ i_input_data[147 % IN_WIDTH];
                536 / IN_WIDTH: pong_storage_data_174 <= (fillup_transition == 1'b1) ? i_input_data[536 % IN_WIDTH] : pong_storage_data_174 ^ i_input_data[536 % IN_WIDTH];
                671 / IN_WIDTH: pong_storage_data_174 <= (fillup_transition == 1'b1) ? i_input_data[671 % IN_WIDTH] : pong_storage_data_174 ^ i_input_data[671 % IN_WIDTH];
                741 / IN_WIDTH: pong_storage_data_174 <= (fillup_transition == 1'b1) ? i_input_data[741 % IN_WIDTH] : pong_storage_data_174 ^ i_input_data[741 % IN_WIDTH];
                1122 / IN_WIDTH: pong_storage_data_174 <= (fillup_transition == 1'b1) ? i_input_data[1122 % IN_WIDTH] : pong_storage_data_174 ^ i_input_data[1122 % IN_WIDTH];
                default: pong_storage_data_174 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_174;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_174 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_174;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_174 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_174;
            end
        end
    end
end

logic ping_storage_data_175;
logic pong_storage_data_175;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_175 <= 1'b0;
        pong_storage_data_175 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                148 / IN_WIDTH: ping_storage_data_175 <= (fillup_transition == 1'b1) ? i_input_data[148 % IN_WIDTH] : ping_storage_data_175 ^ i_input_data[148 % IN_WIDTH];
                537 / IN_WIDTH: ping_storage_data_175 <= (fillup_transition == 1'b1) ? i_input_data[537 % IN_WIDTH] : ping_storage_data_175 ^ i_input_data[537 % IN_WIDTH];
                576 / IN_WIDTH: ping_storage_data_175 <= (fillup_transition == 1'b1) ? i_input_data[576 % IN_WIDTH] : ping_storage_data_175 ^ i_input_data[576 % IN_WIDTH];
                742 / IN_WIDTH: ping_storage_data_175 <= (fillup_transition == 1'b1) ? i_input_data[742 % IN_WIDTH] : ping_storage_data_175 ^ i_input_data[742 % IN_WIDTH];
                1123 / IN_WIDTH: ping_storage_data_175 <= (fillup_transition == 1'b1) ? i_input_data[1123 % IN_WIDTH] : ping_storage_data_175 ^ i_input_data[1123 % IN_WIDTH];
                default: ping_storage_data_175 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_175;
                endcase
            end else begin
                case (input_count)
                148 / IN_WIDTH: pong_storage_data_175 <= (fillup_transition == 1'b1) ? i_input_data[148 % IN_WIDTH] : pong_storage_data_175 ^ i_input_data[148 % IN_WIDTH];
                537 / IN_WIDTH: pong_storage_data_175 <= (fillup_transition == 1'b1) ? i_input_data[537 % IN_WIDTH] : pong_storage_data_175 ^ i_input_data[537 % IN_WIDTH];
                576 / IN_WIDTH: pong_storage_data_175 <= (fillup_transition == 1'b1) ? i_input_data[576 % IN_WIDTH] : pong_storage_data_175 ^ i_input_data[576 % IN_WIDTH];
                742 / IN_WIDTH: pong_storage_data_175 <= (fillup_transition == 1'b1) ? i_input_data[742 % IN_WIDTH] : pong_storage_data_175 ^ i_input_data[742 % IN_WIDTH];
                1123 / IN_WIDTH: pong_storage_data_175 <= (fillup_transition == 1'b1) ? i_input_data[1123 % IN_WIDTH] : pong_storage_data_175 ^ i_input_data[1123 % IN_WIDTH];
                default: pong_storage_data_175 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_175;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_175 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_175;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_175 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_175;
            end
        end
    end
end

logic ping_storage_data_176;
logic pong_storage_data_176;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_176 <= 1'b0;
        pong_storage_data_176 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                149 / IN_WIDTH: ping_storage_data_176 <= (fillup_transition == 1'b1) ? i_input_data[149 % IN_WIDTH] : ping_storage_data_176 ^ i_input_data[149 % IN_WIDTH];
                538 / IN_WIDTH: ping_storage_data_176 <= (fillup_transition == 1'b1) ? i_input_data[538 % IN_WIDTH] : ping_storage_data_176 ^ i_input_data[538 % IN_WIDTH];
                577 / IN_WIDTH: ping_storage_data_176 <= (fillup_transition == 1'b1) ? i_input_data[577 % IN_WIDTH] : ping_storage_data_176 ^ i_input_data[577 % IN_WIDTH];
                743 / IN_WIDTH: ping_storage_data_176 <= (fillup_transition == 1'b1) ? i_input_data[743 % IN_WIDTH] : ping_storage_data_176 ^ i_input_data[743 % IN_WIDTH];
                1124 / IN_WIDTH: ping_storage_data_176 <= (fillup_transition == 1'b1) ? i_input_data[1124 % IN_WIDTH] : ping_storage_data_176 ^ i_input_data[1124 % IN_WIDTH];
                default: ping_storage_data_176 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_176;
                endcase
            end else begin
                case (input_count)
                149 / IN_WIDTH: pong_storage_data_176 <= (fillup_transition == 1'b1) ? i_input_data[149 % IN_WIDTH] : pong_storage_data_176 ^ i_input_data[149 % IN_WIDTH];
                538 / IN_WIDTH: pong_storage_data_176 <= (fillup_transition == 1'b1) ? i_input_data[538 % IN_WIDTH] : pong_storage_data_176 ^ i_input_data[538 % IN_WIDTH];
                577 / IN_WIDTH: pong_storage_data_176 <= (fillup_transition == 1'b1) ? i_input_data[577 % IN_WIDTH] : pong_storage_data_176 ^ i_input_data[577 % IN_WIDTH];
                743 / IN_WIDTH: pong_storage_data_176 <= (fillup_transition == 1'b1) ? i_input_data[743 % IN_WIDTH] : pong_storage_data_176 ^ i_input_data[743 % IN_WIDTH];
                1124 / IN_WIDTH: pong_storage_data_176 <= (fillup_transition == 1'b1) ? i_input_data[1124 % IN_WIDTH] : pong_storage_data_176 ^ i_input_data[1124 % IN_WIDTH];
                default: pong_storage_data_176 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_176;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_176 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_176;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_176 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_176;
            end
        end
    end
end

logic ping_storage_data_177;
logic pong_storage_data_177;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_177 <= 1'b0;
        pong_storage_data_177 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                150 / IN_WIDTH: ping_storage_data_177 <= (fillup_transition == 1'b1) ? i_input_data[150 % IN_WIDTH] : ping_storage_data_177 ^ i_input_data[150 % IN_WIDTH];
                539 / IN_WIDTH: ping_storage_data_177 <= (fillup_transition == 1'b1) ? i_input_data[539 % IN_WIDTH] : ping_storage_data_177 ^ i_input_data[539 % IN_WIDTH];
                578 / IN_WIDTH: ping_storage_data_177 <= (fillup_transition == 1'b1) ? i_input_data[578 % IN_WIDTH] : ping_storage_data_177 ^ i_input_data[578 % IN_WIDTH];
                744 / IN_WIDTH: ping_storage_data_177 <= (fillup_transition == 1'b1) ? i_input_data[744 % IN_WIDTH] : ping_storage_data_177 ^ i_input_data[744 % IN_WIDTH];
                1125 / IN_WIDTH: ping_storage_data_177 <= (fillup_transition == 1'b1) ? i_input_data[1125 % IN_WIDTH] : ping_storage_data_177 ^ i_input_data[1125 % IN_WIDTH];
                default: ping_storage_data_177 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_177;
                endcase
            end else begin
                case (input_count)
                150 / IN_WIDTH: pong_storage_data_177 <= (fillup_transition == 1'b1) ? i_input_data[150 % IN_WIDTH] : pong_storage_data_177 ^ i_input_data[150 % IN_WIDTH];
                539 / IN_WIDTH: pong_storage_data_177 <= (fillup_transition == 1'b1) ? i_input_data[539 % IN_WIDTH] : pong_storage_data_177 ^ i_input_data[539 % IN_WIDTH];
                578 / IN_WIDTH: pong_storage_data_177 <= (fillup_transition == 1'b1) ? i_input_data[578 % IN_WIDTH] : pong_storage_data_177 ^ i_input_data[578 % IN_WIDTH];
                744 / IN_WIDTH: pong_storage_data_177 <= (fillup_transition == 1'b1) ? i_input_data[744 % IN_WIDTH] : pong_storage_data_177 ^ i_input_data[744 % IN_WIDTH];
                1125 / IN_WIDTH: pong_storage_data_177 <= (fillup_transition == 1'b1) ? i_input_data[1125 % IN_WIDTH] : pong_storage_data_177 ^ i_input_data[1125 % IN_WIDTH];
                default: pong_storage_data_177 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_177;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_177 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_177;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_177 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_177;
            end
        end
    end
end

logic ping_storage_data_178;
logic pong_storage_data_178;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_178 <= 1'b0;
        pong_storage_data_178 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                151 / IN_WIDTH: ping_storage_data_178 <= (fillup_transition == 1'b1) ? i_input_data[151 % IN_WIDTH] : ping_storage_data_178 ^ i_input_data[151 % IN_WIDTH];
                540 / IN_WIDTH: ping_storage_data_178 <= (fillup_transition == 1'b1) ? i_input_data[540 % IN_WIDTH] : ping_storage_data_178 ^ i_input_data[540 % IN_WIDTH];
                579 / IN_WIDTH: ping_storage_data_178 <= (fillup_transition == 1'b1) ? i_input_data[579 % IN_WIDTH] : ping_storage_data_178 ^ i_input_data[579 % IN_WIDTH];
                745 / IN_WIDTH: ping_storage_data_178 <= (fillup_transition == 1'b1) ? i_input_data[745 % IN_WIDTH] : ping_storage_data_178 ^ i_input_data[745 % IN_WIDTH];
                1126 / IN_WIDTH: ping_storage_data_178 <= (fillup_transition == 1'b1) ? i_input_data[1126 % IN_WIDTH] : ping_storage_data_178 ^ i_input_data[1126 % IN_WIDTH];
                default: ping_storage_data_178 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_178;
                endcase
            end else begin
                case (input_count)
                151 / IN_WIDTH: pong_storage_data_178 <= (fillup_transition == 1'b1) ? i_input_data[151 % IN_WIDTH] : pong_storage_data_178 ^ i_input_data[151 % IN_WIDTH];
                540 / IN_WIDTH: pong_storage_data_178 <= (fillup_transition == 1'b1) ? i_input_data[540 % IN_WIDTH] : pong_storage_data_178 ^ i_input_data[540 % IN_WIDTH];
                579 / IN_WIDTH: pong_storage_data_178 <= (fillup_transition == 1'b1) ? i_input_data[579 % IN_WIDTH] : pong_storage_data_178 ^ i_input_data[579 % IN_WIDTH];
                745 / IN_WIDTH: pong_storage_data_178 <= (fillup_transition == 1'b1) ? i_input_data[745 % IN_WIDTH] : pong_storage_data_178 ^ i_input_data[745 % IN_WIDTH];
                1126 / IN_WIDTH: pong_storage_data_178 <= (fillup_transition == 1'b1) ? i_input_data[1126 % IN_WIDTH] : pong_storage_data_178 ^ i_input_data[1126 % IN_WIDTH];
                default: pong_storage_data_178 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_178;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_178 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_178;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_178 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_178;
            end
        end
    end
end

logic ping_storage_data_179;
logic pong_storage_data_179;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_179 <= 1'b0;
        pong_storage_data_179 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                152 / IN_WIDTH: ping_storage_data_179 <= (fillup_transition == 1'b1) ? i_input_data[152 % IN_WIDTH] : ping_storage_data_179 ^ i_input_data[152 % IN_WIDTH];
                541 / IN_WIDTH: ping_storage_data_179 <= (fillup_transition == 1'b1) ? i_input_data[541 % IN_WIDTH] : ping_storage_data_179 ^ i_input_data[541 % IN_WIDTH];
                580 / IN_WIDTH: ping_storage_data_179 <= (fillup_transition == 1'b1) ? i_input_data[580 % IN_WIDTH] : ping_storage_data_179 ^ i_input_data[580 % IN_WIDTH];
                746 / IN_WIDTH: ping_storage_data_179 <= (fillup_transition == 1'b1) ? i_input_data[746 % IN_WIDTH] : ping_storage_data_179 ^ i_input_data[746 % IN_WIDTH];
                1127 / IN_WIDTH: ping_storage_data_179 <= (fillup_transition == 1'b1) ? i_input_data[1127 % IN_WIDTH] : ping_storage_data_179 ^ i_input_data[1127 % IN_WIDTH];
                default: ping_storage_data_179 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_179;
                endcase
            end else begin
                case (input_count)
                152 / IN_WIDTH: pong_storage_data_179 <= (fillup_transition == 1'b1) ? i_input_data[152 % IN_WIDTH] : pong_storage_data_179 ^ i_input_data[152 % IN_WIDTH];
                541 / IN_WIDTH: pong_storage_data_179 <= (fillup_transition == 1'b1) ? i_input_data[541 % IN_WIDTH] : pong_storage_data_179 ^ i_input_data[541 % IN_WIDTH];
                580 / IN_WIDTH: pong_storage_data_179 <= (fillup_transition == 1'b1) ? i_input_data[580 % IN_WIDTH] : pong_storage_data_179 ^ i_input_data[580 % IN_WIDTH];
                746 / IN_WIDTH: pong_storage_data_179 <= (fillup_transition == 1'b1) ? i_input_data[746 % IN_WIDTH] : pong_storage_data_179 ^ i_input_data[746 % IN_WIDTH];
                1127 / IN_WIDTH: pong_storage_data_179 <= (fillup_transition == 1'b1) ? i_input_data[1127 % IN_WIDTH] : pong_storage_data_179 ^ i_input_data[1127 % IN_WIDTH];
                default: pong_storage_data_179 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_179;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_179 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_179;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_179 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_179;
            end
        end
    end
end

logic ping_storage_data_180;
logic pong_storage_data_180;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_180 <= 1'b0;
        pong_storage_data_180 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                153 / IN_WIDTH: ping_storage_data_180 <= (fillup_transition == 1'b1) ? i_input_data[153 % IN_WIDTH] : ping_storage_data_180 ^ i_input_data[153 % IN_WIDTH];
                542 / IN_WIDTH: ping_storage_data_180 <= (fillup_transition == 1'b1) ? i_input_data[542 % IN_WIDTH] : ping_storage_data_180 ^ i_input_data[542 % IN_WIDTH];
                581 / IN_WIDTH: ping_storage_data_180 <= (fillup_transition == 1'b1) ? i_input_data[581 % IN_WIDTH] : ping_storage_data_180 ^ i_input_data[581 % IN_WIDTH];
                747 / IN_WIDTH: ping_storage_data_180 <= (fillup_transition == 1'b1) ? i_input_data[747 % IN_WIDTH] : ping_storage_data_180 ^ i_input_data[747 % IN_WIDTH];
                1128 / IN_WIDTH: ping_storage_data_180 <= (fillup_transition == 1'b1) ? i_input_data[1128 % IN_WIDTH] : ping_storage_data_180 ^ i_input_data[1128 % IN_WIDTH];
                default: ping_storage_data_180 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_180;
                endcase
            end else begin
                case (input_count)
                153 / IN_WIDTH: pong_storage_data_180 <= (fillup_transition == 1'b1) ? i_input_data[153 % IN_WIDTH] : pong_storage_data_180 ^ i_input_data[153 % IN_WIDTH];
                542 / IN_WIDTH: pong_storage_data_180 <= (fillup_transition == 1'b1) ? i_input_data[542 % IN_WIDTH] : pong_storage_data_180 ^ i_input_data[542 % IN_WIDTH];
                581 / IN_WIDTH: pong_storage_data_180 <= (fillup_transition == 1'b1) ? i_input_data[581 % IN_WIDTH] : pong_storage_data_180 ^ i_input_data[581 % IN_WIDTH];
                747 / IN_WIDTH: pong_storage_data_180 <= (fillup_transition == 1'b1) ? i_input_data[747 % IN_WIDTH] : pong_storage_data_180 ^ i_input_data[747 % IN_WIDTH];
                1128 / IN_WIDTH: pong_storage_data_180 <= (fillup_transition == 1'b1) ? i_input_data[1128 % IN_WIDTH] : pong_storage_data_180 ^ i_input_data[1128 % IN_WIDTH];
                default: pong_storage_data_180 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_180;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_180 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_180;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_180 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_180;
            end
        end
    end
end

logic ping_storage_data_181;
logic pong_storage_data_181;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_181 <= 1'b0;
        pong_storage_data_181 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                154 / IN_WIDTH: ping_storage_data_181 <= (fillup_transition == 1'b1) ? i_input_data[154 % IN_WIDTH] : ping_storage_data_181 ^ i_input_data[154 % IN_WIDTH];
                543 / IN_WIDTH: ping_storage_data_181 <= (fillup_transition == 1'b1) ? i_input_data[543 % IN_WIDTH] : ping_storage_data_181 ^ i_input_data[543 % IN_WIDTH];
                582 / IN_WIDTH: ping_storage_data_181 <= (fillup_transition == 1'b1) ? i_input_data[582 % IN_WIDTH] : ping_storage_data_181 ^ i_input_data[582 % IN_WIDTH];
                748 / IN_WIDTH: ping_storage_data_181 <= (fillup_transition == 1'b1) ? i_input_data[748 % IN_WIDTH] : ping_storage_data_181 ^ i_input_data[748 % IN_WIDTH];
                1129 / IN_WIDTH: ping_storage_data_181 <= (fillup_transition == 1'b1) ? i_input_data[1129 % IN_WIDTH] : ping_storage_data_181 ^ i_input_data[1129 % IN_WIDTH];
                default: ping_storage_data_181 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_181;
                endcase
            end else begin
                case (input_count)
                154 / IN_WIDTH: pong_storage_data_181 <= (fillup_transition == 1'b1) ? i_input_data[154 % IN_WIDTH] : pong_storage_data_181 ^ i_input_data[154 % IN_WIDTH];
                543 / IN_WIDTH: pong_storage_data_181 <= (fillup_transition == 1'b1) ? i_input_data[543 % IN_WIDTH] : pong_storage_data_181 ^ i_input_data[543 % IN_WIDTH];
                582 / IN_WIDTH: pong_storage_data_181 <= (fillup_transition == 1'b1) ? i_input_data[582 % IN_WIDTH] : pong_storage_data_181 ^ i_input_data[582 % IN_WIDTH];
                748 / IN_WIDTH: pong_storage_data_181 <= (fillup_transition == 1'b1) ? i_input_data[748 % IN_WIDTH] : pong_storage_data_181 ^ i_input_data[748 % IN_WIDTH];
                1129 / IN_WIDTH: pong_storage_data_181 <= (fillup_transition == 1'b1) ? i_input_data[1129 % IN_WIDTH] : pong_storage_data_181 ^ i_input_data[1129 % IN_WIDTH];
                default: pong_storage_data_181 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_181;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_181 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_181;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_181 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_181;
            end
        end
    end
end

logic ping_storage_data_182;
logic pong_storage_data_182;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_182 <= 1'b0;
        pong_storage_data_182 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                155 / IN_WIDTH: ping_storage_data_182 <= (fillup_transition == 1'b1) ? i_input_data[155 % IN_WIDTH] : ping_storage_data_182 ^ i_input_data[155 % IN_WIDTH];
                544 / IN_WIDTH: ping_storage_data_182 <= (fillup_transition == 1'b1) ? i_input_data[544 % IN_WIDTH] : ping_storage_data_182 ^ i_input_data[544 % IN_WIDTH];
                583 / IN_WIDTH: ping_storage_data_182 <= (fillup_transition == 1'b1) ? i_input_data[583 % IN_WIDTH] : ping_storage_data_182 ^ i_input_data[583 % IN_WIDTH];
                749 / IN_WIDTH: ping_storage_data_182 <= (fillup_transition == 1'b1) ? i_input_data[749 % IN_WIDTH] : ping_storage_data_182 ^ i_input_data[749 % IN_WIDTH];
                1130 / IN_WIDTH: ping_storage_data_182 <= (fillup_transition == 1'b1) ? i_input_data[1130 % IN_WIDTH] : ping_storage_data_182 ^ i_input_data[1130 % IN_WIDTH];
                default: ping_storage_data_182 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_182;
                endcase
            end else begin
                case (input_count)
                155 / IN_WIDTH: pong_storage_data_182 <= (fillup_transition == 1'b1) ? i_input_data[155 % IN_WIDTH] : pong_storage_data_182 ^ i_input_data[155 % IN_WIDTH];
                544 / IN_WIDTH: pong_storage_data_182 <= (fillup_transition == 1'b1) ? i_input_data[544 % IN_WIDTH] : pong_storage_data_182 ^ i_input_data[544 % IN_WIDTH];
                583 / IN_WIDTH: pong_storage_data_182 <= (fillup_transition == 1'b1) ? i_input_data[583 % IN_WIDTH] : pong_storage_data_182 ^ i_input_data[583 % IN_WIDTH];
                749 / IN_WIDTH: pong_storage_data_182 <= (fillup_transition == 1'b1) ? i_input_data[749 % IN_WIDTH] : pong_storage_data_182 ^ i_input_data[749 % IN_WIDTH];
                1130 / IN_WIDTH: pong_storage_data_182 <= (fillup_transition == 1'b1) ? i_input_data[1130 % IN_WIDTH] : pong_storage_data_182 ^ i_input_data[1130 % IN_WIDTH];
                default: pong_storage_data_182 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_182;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_182 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_182;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_182 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_182;
            end
        end
    end
end

logic ping_storage_data_183;
logic pong_storage_data_183;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_183 <= 1'b0;
        pong_storage_data_183 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                156 / IN_WIDTH: ping_storage_data_183 <= (fillup_transition == 1'b1) ? i_input_data[156 % IN_WIDTH] : ping_storage_data_183 ^ i_input_data[156 % IN_WIDTH];
                545 / IN_WIDTH: ping_storage_data_183 <= (fillup_transition == 1'b1) ? i_input_data[545 % IN_WIDTH] : ping_storage_data_183 ^ i_input_data[545 % IN_WIDTH];
                584 / IN_WIDTH: ping_storage_data_183 <= (fillup_transition == 1'b1) ? i_input_data[584 % IN_WIDTH] : ping_storage_data_183 ^ i_input_data[584 % IN_WIDTH];
                750 / IN_WIDTH: ping_storage_data_183 <= (fillup_transition == 1'b1) ? i_input_data[750 % IN_WIDTH] : ping_storage_data_183 ^ i_input_data[750 % IN_WIDTH];
                1131 / IN_WIDTH: ping_storage_data_183 <= (fillup_transition == 1'b1) ? i_input_data[1131 % IN_WIDTH] : ping_storage_data_183 ^ i_input_data[1131 % IN_WIDTH];
                default: ping_storage_data_183 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_183;
                endcase
            end else begin
                case (input_count)
                156 / IN_WIDTH: pong_storage_data_183 <= (fillup_transition == 1'b1) ? i_input_data[156 % IN_WIDTH] : pong_storage_data_183 ^ i_input_data[156 % IN_WIDTH];
                545 / IN_WIDTH: pong_storage_data_183 <= (fillup_transition == 1'b1) ? i_input_data[545 % IN_WIDTH] : pong_storage_data_183 ^ i_input_data[545 % IN_WIDTH];
                584 / IN_WIDTH: pong_storage_data_183 <= (fillup_transition == 1'b1) ? i_input_data[584 % IN_WIDTH] : pong_storage_data_183 ^ i_input_data[584 % IN_WIDTH];
                750 / IN_WIDTH: pong_storage_data_183 <= (fillup_transition == 1'b1) ? i_input_data[750 % IN_WIDTH] : pong_storage_data_183 ^ i_input_data[750 % IN_WIDTH];
                1131 / IN_WIDTH: pong_storage_data_183 <= (fillup_transition == 1'b1) ? i_input_data[1131 % IN_WIDTH] : pong_storage_data_183 ^ i_input_data[1131 % IN_WIDTH];
                default: pong_storage_data_183 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_183;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_183 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_183;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_183 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_183;
            end
        end
    end
end

logic ping_storage_data_184;
logic pong_storage_data_184;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_184 <= 1'b0;
        pong_storage_data_184 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                157 / IN_WIDTH: ping_storage_data_184 <= (fillup_transition == 1'b1) ? i_input_data[157 % IN_WIDTH] : ping_storage_data_184 ^ i_input_data[157 % IN_WIDTH];
                546 / IN_WIDTH: ping_storage_data_184 <= (fillup_transition == 1'b1) ? i_input_data[546 % IN_WIDTH] : ping_storage_data_184 ^ i_input_data[546 % IN_WIDTH];
                585 / IN_WIDTH: ping_storage_data_184 <= (fillup_transition == 1'b1) ? i_input_data[585 % IN_WIDTH] : ping_storage_data_184 ^ i_input_data[585 % IN_WIDTH];
                751 / IN_WIDTH: ping_storage_data_184 <= (fillup_transition == 1'b1) ? i_input_data[751 % IN_WIDTH] : ping_storage_data_184 ^ i_input_data[751 % IN_WIDTH];
                1132 / IN_WIDTH: ping_storage_data_184 <= (fillup_transition == 1'b1) ? i_input_data[1132 % IN_WIDTH] : ping_storage_data_184 ^ i_input_data[1132 % IN_WIDTH];
                default: ping_storage_data_184 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_184;
                endcase
            end else begin
                case (input_count)
                157 / IN_WIDTH: pong_storage_data_184 <= (fillup_transition == 1'b1) ? i_input_data[157 % IN_WIDTH] : pong_storage_data_184 ^ i_input_data[157 % IN_WIDTH];
                546 / IN_WIDTH: pong_storage_data_184 <= (fillup_transition == 1'b1) ? i_input_data[546 % IN_WIDTH] : pong_storage_data_184 ^ i_input_data[546 % IN_WIDTH];
                585 / IN_WIDTH: pong_storage_data_184 <= (fillup_transition == 1'b1) ? i_input_data[585 % IN_WIDTH] : pong_storage_data_184 ^ i_input_data[585 % IN_WIDTH];
                751 / IN_WIDTH: pong_storage_data_184 <= (fillup_transition == 1'b1) ? i_input_data[751 % IN_WIDTH] : pong_storage_data_184 ^ i_input_data[751 % IN_WIDTH];
                1132 / IN_WIDTH: pong_storage_data_184 <= (fillup_transition == 1'b1) ? i_input_data[1132 % IN_WIDTH] : pong_storage_data_184 ^ i_input_data[1132 % IN_WIDTH];
                default: pong_storage_data_184 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_184;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_184 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_184;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_184 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_184;
            end
        end
    end
end

logic ping_storage_data_185;
logic pong_storage_data_185;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_185 <= 1'b0;
        pong_storage_data_185 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                158 / IN_WIDTH: ping_storage_data_185 <= (fillup_transition == 1'b1) ? i_input_data[158 % IN_WIDTH] : ping_storage_data_185 ^ i_input_data[158 % IN_WIDTH];
                547 / IN_WIDTH: ping_storage_data_185 <= (fillup_transition == 1'b1) ? i_input_data[547 % IN_WIDTH] : ping_storage_data_185 ^ i_input_data[547 % IN_WIDTH];
                586 / IN_WIDTH: ping_storage_data_185 <= (fillup_transition == 1'b1) ? i_input_data[586 % IN_WIDTH] : ping_storage_data_185 ^ i_input_data[586 % IN_WIDTH];
                752 / IN_WIDTH: ping_storage_data_185 <= (fillup_transition == 1'b1) ? i_input_data[752 % IN_WIDTH] : ping_storage_data_185 ^ i_input_data[752 % IN_WIDTH];
                1133 / IN_WIDTH: ping_storage_data_185 <= (fillup_transition == 1'b1) ? i_input_data[1133 % IN_WIDTH] : ping_storage_data_185 ^ i_input_data[1133 % IN_WIDTH];
                default: ping_storage_data_185 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_185;
                endcase
            end else begin
                case (input_count)
                158 / IN_WIDTH: pong_storage_data_185 <= (fillup_transition == 1'b1) ? i_input_data[158 % IN_WIDTH] : pong_storage_data_185 ^ i_input_data[158 % IN_WIDTH];
                547 / IN_WIDTH: pong_storage_data_185 <= (fillup_transition == 1'b1) ? i_input_data[547 % IN_WIDTH] : pong_storage_data_185 ^ i_input_data[547 % IN_WIDTH];
                586 / IN_WIDTH: pong_storage_data_185 <= (fillup_transition == 1'b1) ? i_input_data[586 % IN_WIDTH] : pong_storage_data_185 ^ i_input_data[586 % IN_WIDTH];
                752 / IN_WIDTH: pong_storage_data_185 <= (fillup_transition == 1'b1) ? i_input_data[752 % IN_WIDTH] : pong_storage_data_185 ^ i_input_data[752 % IN_WIDTH];
                1133 / IN_WIDTH: pong_storage_data_185 <= (fillup_transition == 1'b1) ? i_input_data[1133 % IN_WIDTH] : pong_storage_data_185 ^ i_input_data[1133 % IN_WIDTH];
                default: pong_storage_data_185 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_185;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_185 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_185;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_185 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_185;
            end
        end
    end
end

logic ping_storage_data_186;
logic pong_storage_data_186;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_186 <= 1'b0;
        pong_storage_data_186 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                159 / IN_WIDTH: ping_storage_data_186 <= (fillup_transition == 1'b1) ? i_input_data[159 % IN_WIDTH] : ping_storage_data_186 ^ i_input_data[159 % IN_WIDTH];
                548 / IN_WIDTH: ping_storage_data_186 <= (fillup_transition == 1'b1) ? i_input_data[548 % IN_WIDTH] : ping_storage_data_186 ^ i_input_data[548 % IN_WIDTH];
                587 / IN_WIDTH: ping_storage_data_186 <= (fillup_transition == 1'b1) ? i_input_data[587 % IN_WIDTH] : ping_storage_data_186 ^ i_input_data[587 % IN_WIDTH];
                753 / IN_WIDTH: ping_storage_data_186 <= (fillup_transition == 1'b1) ? i_input_data[753 % IN_WIDTH] : ping_storage_data_186 ^ i_input_data[753 % IN_WIDTH];
                1134 / IN_WIDTH: ping_storage_data_186 <= (fillup_transition == 1'b1) ? i_input_data[1134 % IN_WIDTH] : ping_storage_data_186 ^ i_input_data[1134 % IN_WIDTH];
                default: ping_storage_data_186 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_186;
                endcase
            end else begin
                case (input_count)
                159 / IN_WIDTH: pong_storage_data_186 <= (fillup_transition == 1'b1) ? i_input_data[159 % IN_WIDTH] : pong_storage_data_186 ^ i_input_data[159 % IN_WIDTH];
                548 / IN_WIDTH: pong_storage_data_186 <= (fillup_transition == 1'b1) ? i_input_data[548 % IN_WIDTH] : pong_storage_data_186 ^ i_input_data[548 % IN_WIDTH];
                587 / IN_WIDTH: pong_storage_data_186 <= (fillup_transition == 1'b1) ? i_input_data[587 % IN_WIDTH] : pong_storage_data_186 ^ i_input_data[587 % IN_WIDTH];
                753 / IN_WIDTH: pong_storage_data_186 <= (fillup_transition == 1'b1) ? i_input_data[753 % IN_WIDTH] : pong_storage_data_186 ^ i_input_data[753 % IN_WIDTH];
                1134 / IN_WIDTH: pong_storage_data_186 <= (fillup_transition == 1'b1) ? i_input_data[1134 % IN_WIDTH] : pong_storage_data_186 ^ i_input_data[1134 % IN_WIDTH];
                default: pong_storage_data_186 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_186;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_186 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_186;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_186 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_186;
            end
        end
    end
end

logic ping_storage_data_187;
logic pong_storage_data_187;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_187 <= 1'b0;
        pong_storage_data_187 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                160 / IN_WIDTH: ping_storage_data_187 <= (fillup_transition == 1'b1) ? i_input_data[160 % IN_WIDTH] : ping_storage_data_187 ^ i_input_data[160 % IN_WIDTH];
                549 / IN_WIDTH: ping_storage_data_187 <= (fillup_transition == 1'b1) ? i_input_data[549 % IN_WIDTH] : ping_storage_data_187 ^ i_input_data[549 % IN_WIDTH];
                588 / IN_WIDTH: ping_storage_data_187 <= (fillup_transition == 1'b1) ? i_input_data[588 % IN_WIDTH] : ping_storage_data_187 ^ i_input_data[588 % IN_WIDTH];
                754 / IN_WIDTH: ping_storage_data_187 <= (fillup_transition == 1'b1) ? i_input_data[754 % IN_WIDTH] : ping_storage_data_187 ^ i_input_data[754 % IN_WIDTH];
                1135 / IN_WIDTH: ping_storage_data_187 <= (fillup_transition == 1'b1) ? i_input_data[1135 % IN_WIDTH] : ping_storage_data_187 ^ i_input_data[1135 % IN_WIDTH];
                default: ping_storage_data_187 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_187;
                endcase
            end else begin
                case (input_count)
                160 / IN_WIDTH: pong_storage_data_187 <= (fillup_transition == 1'b1) ? i_input_data[160 % IN_WIDTH] : pong_storage_data_187 ^ i_input_data[160 % IN_WIDTH];
                549 / IN_WIDTH: pong_storage_data_187 <= (fillup_transition == 1'b1) ? i_input_data[549 % IN_WIDTH] : pong_storage_data_187 ^ i_input_data[549 % IN_WIDTH];
                588 / IN_WIDTH: pong_storage_data_187 <= (fillup_transition == 1'b1) ? i_input_data[588 % IN_WIDTH] : pong_storage_data_187 ^ i_input_data[588 % IN_WIDTH];
                754 / IN_WIDTH: pong_storage_data_187 <= (fillup_transition == 1'b1) ? i_input_data[754 % IN_WIDTH] : pong_storage_data_187 ^ i_input_data[754 % IN_WIDTH];
                1135 / IN_WIDTH: pong_storage_data_187 <= (fillup_transition == 1'b1) ? i_input_data[1135 % IN_WIDTH] : pong_storage_data_187 ^ i_input_data[1135 % IN_WIDTH];
                default: pong_storage_data_187 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_187;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_187 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_187;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_187 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_187;
            end
        end
    end
end

logic ping_storage_data_188;
logic pong_storage_data_188;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_188 <= 1'b0;
        pong_storage_data_188 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                161 / IN_WIDTH: ping_storage_data_188 <= (fillup_transition == 1'b1) ? i_input_data[161 % IN_WIDTH] : ping_storage_data_188 ^ i_input_data[161 % IN_WIDTH];
                550 / IN_WIDTH: ping_storage_data_188 <= (fillup_transition == 1'b1) ? i_input_data[550 % IN_WIDTH] : ping_storage_data_188 ^ i_input_data[550 % IN_WIDTH];
                589 / IN_WIDTH: ping_storage_data_188 <= (fillup_transition == 1'b1) ? i_input_data[589 % IN_WIDTH] : ping_storage_data_188 ^ i_input_data[589 % IN_WIDTH];
                755 / IN_WIDTH: ping_storage_data_188 <= (fillup_transition == 1'b1) ? i_input_data[755 % IN_WIDTH] : ping_storage_data_188 ^ i_input_data[755 % IN_WIDTH];
                1136 / IN_WIDTH: ping_storage_data_188 <= (fillup_transition == 1'b1) ? i_input_data[1136 % IN_WIDTH] : ping_storage_data_188 ^ i_input_data[1136 % IN_WIDTH];
                default: ping_storage_data_188 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_188;
                endcase
            end else begin
                case (input_count)
                161 / IN_WIDTH: pong_storage_data_188 <= (fillup_transition == 1'b1) ? i_input_data[161 % IN_WIDTH] : pong_storage_data_188 ^ i_input_data[161 % IN_WIDTH];
                550 / IN_WIDTH: pong_storage_data_188 <= (fillup_transition == 1'b1) ? i_input_data[550 % IN_WIDTH] : pong_storage_data_188 ^ i_input_data[550 % IN_WIDTH];
                589 / IN_WIDTH: pong_storage_data_188 <= (fillup_transition == 1'b1) ? i_input_data[589 % IN_WIDTH] : pong_storage_data_188 ^ i_input_data[589 % IN_WIDTH];
                755 / IN_WIDTH: pong_storage_data_188 <= (fillup_transition == 1'b1) ? i_input_data[755 % IN_WIDTH] : pong_storage_data_188 ^ i_input_data[755 % IN_WIDTH];
                1136 / IN_WIDTH: pong_storage_data_188 <= (fillup_transition == 1'b1) ? i_input_data[1136 % IN_WIDTH] : pong_storage_data_188 ^ i_input_data[1136 % IN_WIDTH];
                default: pong_storage_data_188 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_188;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_188 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_188;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_188 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_188;
            end
        end
    end
end

logic ping_storage_data_189;
logic pong_storage_data_189;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_189 <= 1'b0;
        pong_storage_data_189 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                162 / IN_WIDTH: ping_storage_data_189 <= (fillup_transition == 1'b1) ? i_input_data[162 % IN_WIDTH] : ping_storage_data_189 ^ i_input_data[162 % IN_WIDTH];
                551 / IN_WIDTH: ping_storage_data_189 <= (fillup_transition == 1'b1) ? i_input_data[551 % IN_WIDTH] : ping_storage_data_189 ^ i_input_data[551 % IN_WIDTH];
                590 / IN_WIDTH: ping_storage_data_189 <= (fillup_transition == 1'b1) ? i_input_data[590 % IN_WIDTH] : ping_storage_data_189 ^ i_input_data[590 % IN_WIDTH];
                756 / IN_WIDTH: ping_storage_data_189 <= (fillup_transition == 1'b1) ? i_input_data[756 % IN_WIDTH] : ping_storage_data_189 ^ i_input_data[756 % IN_WIDTH];
                1137 / IN_WIDTH: ping_storage_data_189 <= (fillup_transition == 1'b1) ? i_input_data[1137 % IN_WIDTH] : ping_storage_data_189 ^ i_input_data[1137 % IN_WIDTH];
                default: ping_storage_data_189 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_189;
                endcase
            end else begin
                case (input_count)
                162 / IN_WIDTH: pong_storage_data_189 <= (fillup_transition == 1'b1) ? i_input_data[162 % IN_WIDTH] : pong_storage_data_189 ^ i_input_data[162 % IN_WIDTH];
                551 / IN_WIDTH: pong_storage_data_189 <= (fillup_transition == 1'b1) ? i_input_data[551 % IN_WIDTH] : pong_storage_data_189 ^ i_input_data[551 % IN_WIDTH];
                590 / IN_WIDTH: pong_storage_data_189 <= (fillup_transition == 1'b1) ? i_input_data[590 % IN_WIDTH] : pong_storage_data_189 ^ i_input_data[590 % IN_WIDTH];
                756 / IN_WIDTH: pong_storage_data_189 <= (fillup_transition == 1'b1) ? i_input_data[756 % IN_WIDTH] : pong_storage_data_189 ^ i_input_data[756 % IN_WIDTH];
                1137 / IN_WIDTH: pong_storage_data_189 <= (fillup_transition == 1'b1) ? i_input_data[1137 % IN_WIDTH] : pong_storage_data_189 ^ i_input_data[1137 % IN_WIDTH];
                default: pong_storage_data_189 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_189;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_189 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_189;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_189 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_189;
            end
        end
    end
end

logic ping_storage_data_190;
logic pong_storage_data_190;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_190 <= 1'b0;
        pong_storage_data_190 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                163 / IN_WIDTH: ping_storage_data_190 <= (fillup_transition == 1'b1) ? i_input_data[163 % IN_WIDTH] : ping_storage_data_190 ^ i_input_data[163 % IN_WIDTH];
                552 / IN_WIDTH: ping_storage_data_190 <= (fillup_transition == 1'b1) ? i_input_data[552 % IN_WIDTH] : ping_storage_data_190 ^ i_input_data[552 % IN_WIDTH];
                591 / IN_WIDTH: ping_storage_data_190 <= (fillup_transition == 1'b1) ? i_input_data[591 % IN_WIDTH] : ping_storage_data_190 ^ i_input_data[591 % IN_WIDTH];
                757 / IN_WIDTH: ping_storage_data_190 <= (fillup_transition == 1'b1) ? i_input_data[757 % IN_WIDTH] : ping_storage_data_190 ^ i_input_data[757 % IN_WIDTH];
                1138 / IN_WIDTH: ping_storage_data_190 <= (fillup_transition == 1'b1) ? i_input_data[1138 % IN_WIDTH] : ping_storage_data_190 ^ i_input_data[1138 % IN_WIDTH];
                default: ping_storage_data_190 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_190;
                endcase
            end else begin
                case (input_count)
                163 / IN_WIDTH: pong_storage_data_190 <= (fillup_transition == 1'b1) ? i_input_data[163 % IN_WIDTH] : pong_storage_data_190 ^ i_input_data[163 % IN_WIDTH];
                552 / IN_WIDTH: pong_storage_data_190 <= (fillup_transition == 1'b1) ? i_input_data[552 % IN_WIDTH] : pong_storage_data_190 ^ i_input_data[552 % IN_WIDTH];
                591 / IN_WIDTH: pong_storage_data_190 <= (fillup_transition == 1'b1) ? i_input_data[591 % IN_WIDTH] : pong_storage_data_190 ^ i_input_data[591 % IN_WIDTH];
                757 / IN_WIDTH: pong_storage_data_190 <= (fillup_transition == 1'b1) ? i_input_data[757 % IN_WIDTH] : pong_storage_data_190 ^ i_input_data[757 % IN_WIDTH];
                1138 / IN_WIDTH: pong_storage_data_190 <= (fillup_transition == 1'b1) ? i_input_data[1138 % IN_WIDTH] : pong_storage_data_190 ^ i_input_data[1138 % IN_WIDTH];
                default: pong_storage_data_190 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_190;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_190 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_190;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_190 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_190;
            end
        end
    end
end

logic ping_storage_data_191;
logic pong_storage_data_191;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_191 <= 1'b0;
        pong_storage_data_191 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                164 / IN_WIDTH: ping_storage_data_191 <= (fillup_transition == 1'b1) ? i_input_data[164 % IN_WIDTH] : ping_storage_data_191 ^ i_input_data[164 % IN_WIDTH];
                553 / IN_WIDTH: ping_storage_data_191 <= (fillup_transition == 1'b1) ? i_input_data[553 % IN_WIDTH] : ping_storage_data_191 ^ i_input_data[553 % IN_WIDTH];
                592 / IN_WIDTH: ping_storage_data_191 <= (fillup_transition == 1'b1) ? i_input_data[592 % IN_WIDTH] : ping_storage_data_191 ^ i_input_data[592 % IN_WIDTH];
                758 / IN_WIDTH: ping_storage_data_191 <= (fillup_transition == 1'b1) ? i_input_data[758 % IN_WIDTH] : ping_storage_data_191 ^ i_input_data[758 % IN_WIDTH];
                1139 / IN_WIDTH: ping_storage_data_191 <= (fillup_transition == 1'b1) ? i_input_data[1139 % IN_WIDTH] : ping_storage_data_191 ^ i_input_data[1139 % IN_WIDTH];
                default: ping_storage_data_191 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_191;
                endcase
            end else begin
                case (input_count)
                164 / IN_WIDTH: pong_storage_data_191 <= (fillup_transition == 1'b1) ? i_input_data[164 % IN_WIDTH] : pong_storage_data_191 ^ i_input_data[164 % IN_WIDTH];
                553 / IN_WIDTH: pong_storage_data_191 <= (fillup_transition == 1'b1) ? i_input_data[553 % IN_WIDTH] : pong_storage_data_191 ^ i_input_data[553 % IN_WIDTH];
                592 / IN_WIDTH: pong_storage_data_191 <= (fillup_transition == 1'b1) ? i_input_data[592 % IN_WIDTH] : pong_storage_data_191 ^ i_input_data[592 % IN_WIDTH];
                758 / IN_WIDTH: pong_storage_data_191 <= (fillup_transition == 1'b1) ? i_input_data[758 % IN_WIDTH] : pong_storage_data_191 ^ i_input_data[758 % IN_WIDTH];
                1139 / IN_WIDTH: pong_storage_data_191 <= (fillup_transition == 1'b1) ? i_input_data[1139 % IN_WIDTH] : pong_storage_data_191 ^ i_input_data[1139 % IN_WIDTH];
                default: pong_storage_data_191 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_191;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_191 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_191;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_191 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_191;
            end
        end
    end
end

logic ping_storage_data_192;
logic pong_storage_data_192;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_192 <= 1'b0;
        pong_storage_data_192 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                360 / IN_WIDTH: ping_storage_data_192 <= (fillup_transition == 1'b1) ? i_input_data[360 % IN_WIDTH] : ping_storage_data_192 ^ i_input_data[360 % IN_WIDTH];
                458 / IN_WIDTH: ping_storage_data_192 <= (fillup_transition == 1'b1) ? i_input_data[458 % IN_WIDTH] : ping_storage_data_192 ^ i_input_data[458 % IN_WIDTH];
                495 / IN_WIDTH: ping_storage_data_192 <= (fillup_transition == 1'b1) ? i_input_data[495 % IN_WIDTH] : ping_storage_data_192 ^ i_input_data[495 % IN_WIDTH];
                735 / IN_WIDTH: ping_storage_data_192 <= (fillup_transition == 1'b1) ? i_input_data[735 % IN_WIDTH] : ping_storage_data_192 ^ i_input_data[735 % IN_WIDTH];
                1056 / IN_WIDTH: ping_storage_data_192 <= (fillup_transition == 1'b1) ? i_input_data[1056 % IN_WIDTH] : ping_storage_data_192 ^ i_input_data[1056 % IN_WIDTH];
                default: ping_storage_data_192 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_192;
                endcase
            end else begin
                case (input_count)
                360 / IN_WIDTH: pong_storage_data_192 <= (fillup_transition == 1'b1) ? i_input_data[360 % IN_WIDTH] : pong_storage_data_192 ^ i_input_data[360 % IN_WIDTH];
                458 / IN_WIDTH: pong_storage_data_192 <= (fillup_transition == 1'b1) ? i_input_data[458 % IN_WIDTH] : pong_storage_data_192 ^ i_input_data[458 % IN_WIDTH];
                495 / IN_WIDTH: pong_storage_data_192 <= (fillup_transition == 1'b1) ? i_input_data[495 % IN_WIDTH] : pong_storage_data_192 ^ i_input_data[495 % IN_WIDTH];
                735 / IN_WIDTH: pong_storage_data_192 <= (fillup_transition == 1'b1) ? i_input_data[735 % IN_WIDTH] : pong_storage_data_192 ^ i_input_data[735 % IN_WIDTH];
                1056 / IN_WIDTH: pong_storage_data_192 <= (fillup_transition == 1'b1) ? i_input_data[1056 % IN_WIDTH] : pong_storage_data_192 ^ i_input_data[1056 % IN_WIDTH];
                default: pong_storage_data_192 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_192;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_192 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_192;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_192 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_192;
            end
        end
    end
end

logic ping_storage_data_193;
logic pong_storage_data_193;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_193 <= 1'b0;
        pong_storage_data_193 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                361 / IN_WIDTH: ping_storage_data_193 <= (fillup_transition == 1'b1) ? i_input_data[361 % IN_WIDTH] : ping_storage_data_193 ^ i_input_data[361 % IN_WIDTH];
                459 / IN_WIDTH: ping_storage_data_193 <= (fillup_transition == 1'b1) ? i_input_data[459 % IN_WIDTH] : ping_storage_data_193 ^ i_input_data[459 % IN_WIDTH];
                496 / IN_WIDTH: ping_storage_data_193 <= (fillup_transition == 1'b1) ? i_input_data[496 % IN_WIDTH] : ping_storage_data_193 ^ i_input_data[496 % IN_WIDTH];
                736 / IN_WIDTH: ping_storage_data_193 <= (fillup_transition == 1'b1) ? i_input_data[736 % IN_WIDTH] : ping_storage_data_193 ^ i_input_data[736 % IN_WIDTH];
                1057 / IN_WIDTH: ping_storage_data_193 <= (fillup_transition == 1'b1) ? i_input_data[1057 % IN_WIDTH] : ping_storage_data_193 ^ i_input_data[1057 % IN_WIDTH];
                default: ping_storage_data_193 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_193;
                endcase
            end else begin
                case (input_count)
                361 / IN_WIDTH: pong_storage_data_193 <= (fillup_transition == 1'b1) ? i_input_data[361 % IN_WIDTH] : pong_storage_data_193 ^ i_input_data[361 % IN_WIDTH];
                459 / IN_WIDTH: pong_storage_data_193 <= (fillup_transition == 1'b1) ? i_input_data[459 % IN_WIDTH] : pong_storage_data_193 ^ i_input_data[459 % IN_WIDTH];
                496 / IN_WIDTH: pong_storage_data_193 <= (fillup_transition == 1'b1) ? i_input_data[496 % IN_WIDTH] : pong_storage_data_193 ^ i_input_data[496 % IN_WIDTH];
                736 / IN_WIDTH: pong_storage_data_193 <= (fillup_transition == 1'b1) ? i_input_data[736 % IN_WIDTH] : pong_storage_data_193 ^ i_input_data[736 % IN_WIDTH];
                1057 / IN_WIDTH: pong_storage_data_193 <= (fillup_transition == 1'b1) ? i_input_data[1057 % IN_WIDTH] : pong_storage_data_193 ^ i_input_data[1057 % IN_WIDTH];
                default: pong_storage_data_193 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_193;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_193 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_193;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_193 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_193;
            end
        end
    end
end

logic ping_storage_data_194;
logic pong_storage_data_194;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_194 <= 1'b0;
        pong_storage_data_194 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                362 / IN_WIDTH: ping_storage_data_194 <= (fillup_transition == 1'b1) ? i_input_data[362 % IN_WIDTH] : ping_storage_data_194 ^ i_input_data[362 % IN_WIDTH];
                460 / IN_WIDTH: ping_storage_data_194 <= (fillup_transition == 1'b1) ? i_input_data[460 % IN_WIDTH] : ping_storage_data_194 ^ i_input_data[460 % IN_WIDTH];
                497 / IN_WIDTH: ping_storage_data_194 <= (fillup_transition == 1'b1) ? i_input_data[497 % IN_WIDTH] : ping_storage_data_194 ^ i_input_data[497 % IN_WIDTH];
                737 / IN_WIDTH: ping_storage_data_194 <= (fillup_transition == 1'b1) ? i_input_data[737 % IN_WIDTH] : ping_storage_data_194 ^ i_input_data[737 % IN_WIDTH];
                1058 / IN_WIDTH: ping_storage_data_194 <= (fillup_transition == 1'b1) ? i_input_data[1058 % IN_WIDTH] : ping_storage_data_194 ^ i_input_data[1058 % IN_WIDTH];
                default: ping_storage_data_194 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_194;
                endcase
            end else begin
                case (input_count)
                362 / IN_WIDTH: pong_storage_data_194 <= (fillup_transition == 1'b1) ? i_input_data[362 % IN_WIDTH] : pong_storage_data_194 ^ i_input_data[362 % IN_WIDTH];
                460 / IN_WIDTH: pong_storage_data_194 <= (fillup_transition == 1'b1) ? i_input_data[460 % IN_WIDTH] : pong_storage_data_194 ^ i_input_data[460 % IN_WIDTH];
                497 / IN_WIDTH: pong_storage_data_194 <= (fillup_transition == 1'b1) ? i_input_data[497 % IN_WIDTH] : pong_storage_data_194 ^ i_input_data[497 % IN_WIDTH];
                737 / IN_WIDTH: pong_storage_data_194 <= (fillup_transition == 1'b1) ? i_input_data[737 % IN_WIDTH] : pong_storage_data_194 ^ i_input_data[737 % IN_WIDTH];
                1058 / IN_WIDTH: pong_storage_data_194 <= (fillup_transition == 1'b1) ? i_input_data[1058 % IN_WIDTH] : pong_storage_data_194 ^ i_input_data[1058 % IN_WIDTH];
                default: pong_storage_data_194 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_194;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_194 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_194;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_194 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_194;
            end
        end
    end
end

logic ping_storage_data_195;
logic pong_storage_data_195;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_195 <= 1'b0;
        pong_storage_data_195 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                363 / IN_WIDTH: ping_storage_data_195 <= (fillup_transition == 1'b1) ? i_input_data[363 % IN_WIDTH] : ping_storage_data_195 ^ i_input_data[363 % IN_WIDTH];
                461 / IN_WIDTH: ping_storage_data_195 <= (fillup_transition == 1'b1) ? i_input_data[461 % IN_WIDTH] : ping_storage_data_195 ^ i_input_data[461 % IN_WIDTH];
                498 / IN_WIDTH: ping_storage_data_195 <= (fillup_transition == 1'b1) ? i_input_data[498 % IN_WIDTH] : ping_storage_data_195 ^ i_input_data[498 % IN_WIDTH];
                738 / IN_WIDTH: ping_storage_data_195 <= (fillup_transition == 1'b1) ? i_input_data[738 % IN_WIDTH] : ping_storage_data_195 ^ i_input_data[738 % IN_WIDTH];
                1059 / IN_WIDTH: ping_storage_data_195 <= (fillup_transition == 1'b1) ? i_input_data[1059 % IN_WIDTH] : ping_storage_data_195 ^ i_input_data[1059 % IN_WIDTH];
                default: ping_storage_data_195 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_195;
                endcase
            end else begin
                case (input_count)
                363 / IN_WIDTH: pong_storage_data_195 <= (fillup_transition == 1'b1) ? i_input_data[363 % IN_WIDTH] : pong_storage_data_195 ^ i_input_data[363 % IN_WIDTH];
                461 / IN_WIDTH: pong_storage_data_195 <= (fillup_transition == 1'b1) ? i_input_data[461 % IN_WIDTH] : pong_storage_data_195 ^ i_input_data[461 % IN_WIDTH];
                498 / IN_WIDTH: pong_storage_data_195 <= (fillup_transition == 1'b1) ? i_input_data[498 % IN_WIDTH] : pong_storage_data_195 ^ i_input_data[498 % IN_WIDTH];
                738 / IN_WIDTH: pong_storage_data_195 <= (fillup_transition == 1'b1) ? i_input_data[738 % IN_WIDTH] : pong_storage_data_195 ^ i_input_data[738 % IN_WIDTH];
                1059 / IN_WIDTH: pong_storage_data_195 <= (fillup_transition == 1'b1) ? i_input_data[1059 % IN_WIDTH] : pong_storage_data_195 ^ i_input_data[1059 % IN_WIDTH];
                default: pong_storage_data_195 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_195;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_195 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_195;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_195 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_195;
            end
        end
    end
end

logic ping_storage_data_196;
logic pong_storage_data_196;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_196 <= 1'b0;
        pong_storage_data_196 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                364 / IN_WIDTH: ping_storage_data_196 <= (fillup_transition == 1'b1) ? i_input_data[364 % IN_WIDTH] : ping_storage_data_196 ^ i_input_data[364 % IN_WIDTH];
                462 / IN_WIDTH: ping_storage_data_196 <= (fillup_transition == 1'b1) ? i_input_data[462 % IN_WIDTH] : ping_storage_data_196 ^ i_input_data[462 % IN_WIDTH];
                499 / IN_WIDTH: ping_storage_data_196 <= (fillup_transition == 1'b1) ? i_input_data[499 % IN_WIDTH] : ping_storage_data_196 ^ i_input_data[499 % IN_WIDTH];
                739 / IN_WIDTH: ping_storage_data_196 <= (fillup_transition == 1'b1) ? i_input_data[739 % IN_WIDTH] : ping_storage_data_196 ^ i_input_data[739 % IN_WIDTH];
                1060 / IN_WIDTH: ping_storage_data_196 <= (fillup_transition == 1'b1) ? i_input_data[1060 % IN_WIDTH] : ping_storage_data_196 ^ i_input_data[1060 % IN_WIDTH];
                default: ping_storage_data_196 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_196;
                endcase
            end else begin
                case (input_count)
                364 / IN_WIDTH: pong_storage_data_196 <= (fillup_transition == 1'b1) ? i_input_data[364 % IN_WIDTH] : pong_storage_data_196 ^ i_input_data[364 % IN_WIDTH];
                462 / IN_WIDTH: pong_storage_data_196 <= (fillup_transition == 1'b1) ? i_input_data[462 % IN_WIDTH] : pong_storage_data_196 ^ i_input_data[462 % IN_WIDTH];
                499 / IN_WIDTH: pong_storage_data_196 <= (fillup_transition == 1'b1) ? i_input_data[499 % IN_WIDTH] : pong_storage_data_196 ^ i_input_data[499 % IN_WIDTH];
                739 / IN_WIDTH: pong_storage_data_196 <= (fillup_transition == 1'b1) ? i_input_data[739 % IN_WIDTH] : pong_storage_data_196 ^ i_input_data[739 % IN_WIDTH];
                1060 / IN_WIDTH: pong_storage_data_196 <= (fillup_transition == 1'b1) ? i_input_data[1060 % IN_WIDTH] : pong_storage_data_196 ^ i_input_data[1060 % IN_WIDTH];
                default: pong_storage_data_196 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_196;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_196 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_196;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_196 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_196;
            end
        end
    end
end

logic ping_storage_data_197;
logic pong_storage_data_197;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_197 <= 1'b0;
        pong_storage_data_197 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                365 / IN_WIDTH: ping_storage_data_197 <= (fillup_transition == 1'b1) ? i_input_data[365 % IN_WIDTH] : ping_storage_data_197 ^ i_input_data[365 % IN_WIDTH];
                463 / IN_WIDTH: ping_storage_data_197 <= (fillup_transition == 1'b1) ? i_input_data[463 % IN_WIDTH] : ping_storage_data_197 ^ i_input_data[463 % IN_WIDTH];
                500 / IN_WIDTH: ping_storage_data_197 <= (fillup_transition == 1'b1) ? i_input_data[500 % IN_WIDTH] : ping_storage_data_197 ^ i_input_data[500 % IN_WIDTH];
                740 / IN_WIDTH: ping_storage_data_197 <= (fillup_transition == 1'b1) ? i_input_data[740 % IN_WIDTH] : ping_storage_data_197 ^ i_input_data[740 % IN_WIDTH];
                1061 / IN_WIDTH: ping_storage_data_197 <= (fillup_transition == 1'b1) ? i_input_data[1061 % IN_WIDTH] : ping_storage_data_197 ^ i_input_data[1061 % IN_WIDTH];
                default: ping_storage_data_197 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_197;
                endcase
            end else begin
                case (input_count)
                365 / IN_WIDTH: pong_storage_data_197 <= (fillup_transition == 1'b1) ? i_input_data[365 % IN_WIDTH] : pong_storage_data_197 ^ i_input_data[365 % IN_WIDTH];
                463 / IN_WIDTH: pong_storage_data_197 <= (fillup_transition == 1'b1) ? i_input_data[463 % IN_WIDTH] : pong_storage_data_197 ^ i_input_data[463 % IN_WIDTH];
                500 / IN_WIDTH: pong_storage_data_197 <= (fillup_transition == 1'b1) ? i_input_data[500 % IN_WIDTH] : pong_storage_data_197 ^ i_input_data[500 % IN_WIDTH];
                740 / IN_WIDTH: pong_storage_data_197 <= (fillup_transition == 1'b1) ? i_input_data[740 % IN_WIDTH] : pong_storage_data_197 ^ i_input_data[740 % IN_WIDTH];
                1061 / IN_WIDTH: pong_storage_data_197 <= (fillup_transition == 1'b1) ? i_input_data[1061 % IN_WIDTH] : pong_storage_data_197 ^ i_input_data[1061 % IN_WIDTH];
                default: pong_storage_data_197 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_197;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_197 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_197;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_197 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_197;
            end
        end
    end
end

logic ping_storage_data_198;
logic pong_storage_data_198;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_198 <= 1'b0;
        pong_storage_data_198 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                366 / IN_WIDTH: ping_storage_data_198 <= (fillup_transition == 1'b1) ? i_input_data[366 % IN_WIDTH] : ping_storage_data_198 ^ i_input_data[366 % IN_WIDTH];
                464 / IN_WIDTH: ping_storage_data_198 <= (fillup_transition == 1'b1) ? i_input_data[464 % IN_WIDTH] : ping_storage_data_198 ^ i_input_data[464 % IN_WIDTH];
                501 / IN_WIDTH: ping_storage_data_198 <= (fillup_transition == 1'b1) ? i_input_data[501 % IN_WIDTH] : ping_storage_data_198 ^ i_input_data[501 % IN_WIDTH];
                741 / IN_WIDTH: ping_storage_data_198 <= (fillup_transition == 1'b1) ? i_input_data[741 % IN_WIDTH] : ping_storage_data_198 ^ i_input_data[741 % IN_WIDTH];
                1062 / IN_WIDTH: ping_storage_data_198 <= (fillup_transition == 1'b1) ? i_input_data[1062 % IN_WIDTH] : ping_storage_data_198 ^ i_input_data[1062 % IN_WIDTH];
                default: ping_storage_data_198 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_198;
                endcase
            end else begin
                case (input_count)
                366 / IN_WIDTH: pong_storage_data_198 <= (fillup_transition == 1'b1) ? i_input_data[366 % IN_WIDTH] : pong_storage_data_198 ^ i_input_data[366 % IN_WIDTH];
                464 / IN_WIDTH: pong_storage_data_198 <= (fillup_transition == 1'b1) ? i_input_data[464 % IN_WIDTH] : pong_storage_data_198 ^ i_input_data[464 % IN_WIDTH];
                501 / IN_WIDTH: pong_storage_data_198 <= (fillup_transition == 1'b1) ? i_input_data[501 % IN_WIDTH] : pong_storage_data_198 ^ i_input_data[501 % IN_WIDTH];
                741 / IN_WIDTH: pong_storage_data_198 <= (fillup_transition == 1'b1) ? i_input_data[741 % IN_WIDTH] : pong_storage_data_198 ^ i_input_data[741 % IN_WIDTH];
                1062 / IN_WIDTH: pong_storage_data_198 <= (fillup_transition == 1'b1) ? i_input_data[1062 % IN_WIDTH] : pong_storage_data_198 ^ i_input_data[1062 % IN_WIDTH];
                default: pong_storage_data_198 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_198;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_198 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_198;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_198 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_198;
            end
        end
    end
end

logic ping_storage_data_199;
logic pong_storage_data_199;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_199 <= 1'b0;
        pong_storage_data_199 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                367 / IN_WIDTH: ping_storage_data_199 <= (fillup_transition == 1'b1) ? i_input_data[367 % IN_WIDTH] : ping_storage_data_199 ^ i_input_data[367 % IN_WIDTH];
                465 / IN_WIDTH: ping_storage_data_199 <= (fillup_transition == 1'b1) ? i_input_data[465 % IN_WIDTH] : ping_storage_data_199 ^ i_input_data[465 % IN_WIDTH];
                502 / IN_WIDTH: ping_storage_data_199 <= (fillup_transition == 1'b1) ? i_input_data[502 % IN_WIDTH] : ping_storage_data_199 ^ i_input_data[502 % IN_WIDTH];
                742 / IN_WIDTH: ping_storage_data_199 <= (fillup_transition == 1'b1) ? i_input_data[742 % IN_WIDTH] : ping_storage_data_199 ^ i_input_data[742 % IN_WIDTH];
                1063 / IN_WIDTH: ping_storage_data_199 <= (fillup_transition == 1'b1) ? i_input_data[1063 % IN_WIDTH] : ping_storage_data_199 ^ i_input_data[1063 % IN_WIDTH];
                default: ping_storage_data_199 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_199;
                endcase
            end else begin
                case (input_count)
                367 / IN_WIDTH: pong_storage_data_199 <= (fillup_transition == 1'b1) ? i_input_data[367 % IN_WIDTH] : pong_storage_data_199 ^ i_input_data[367 % IN_WIDTH];
                465 / IN_WIDTH: pong_storage_data_199 <= (fillup_transition == 1'b1) ? i_input_data[465 % IN_WIDTH] : pong_storage_data_199 ^ i_input_data[465 % IN_WIDTH];
                502 / IN_WIDTH: pong_storage_data_199 <= (fillup_transition == 1'b1) ? i_input_data[502 % IN_WIDTH] : pong_storage_data_199 ^ i_input_data[502 % IN_WIDTH];
                742 / IN_WIDTH: pong_storage_data_199 <= (fillup_transition == 1'b1) ? i_input_data[742 % IN_WIDTH] : pong_storage_data_199 ^ i_input_data[742 % IN_WIDTH];
                1063 / IN_WIDTH: pong_storage_data_199 <= (fillup_transition == 1'b1) ? i_input_data[1063 % IN_WIDTH] : pong_storage_data_199 ^ i_input_data[1063 % IN_WIDTH];
                default: pong_storage_data_199 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_199;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_199 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_199;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_199 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_199;
            end
        end
    end
end

logic ping_storage_data_200;
logic pong_storage_data_200;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_200 <= 1'b0;
        pong_storage_data_200 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                368 / IN_WIDTH: ping_storage_data_200 <= (fillup_transition == 1'b1) ? i_input_data[368 % IN_WIDTH] : ping_storage_data_200 ^ i_input_data[368 % IN_WIDTH];
                466 / IN_WIDTH: ping_storage_data_200 <= (fillup_transition == 1'b1) ? i_input_data[466 % IN_WIDTH] : ping_storage_data_200 ^ i_input_data[466 % IN_WIDTH];
                503 / IN_WIDTH: ping_storage_data_200 <= (fillup_transition == 1'b1) ? i_input_data[503 % IN_WIDTH] : ping_storage_data_200 ^ i_input_data[503 % IN_WIDTH];
                743 / IN_WIDTH: ping_storage_data_200 <= (fillup_transition == 1'b1) ? i_input_data[743 % IN_WIDTH] : ping_storage_data_200 ^ i_input_data[743 % IN_WIDTH];
                1064 / IN_WIDTH: ping_storage_data_200 <= (fillup_transition == 1'b1) ? i_input_data[1064 % IN_WIDTH] : ping_storage_data_200 ^ i_input_data[1064 % IN_WIDTH];
                default: ping_storage_data_200 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_200;
                endcase
            end else begin
                case (input_count)
                368 / IN_WIDTH: pong_storage_data_200 <= (fillup_transition == 1'b1) ? i_input_data[368 % IN_WIDTH] : pong_storage_data_200 ^ i_input_data[368 % IN_WIDTH];
                466 / IN_WIDTH: pong_storage_data_200 <= (fillup_transition == 1'b1) ? i_input_data[466 % IN_WIDTH] : pong_storage_data_200 ^ i_input_data[466 % IN_WIDTH];
                503 / IN_WIDTH: pong_storage_data_200 <= (fillup_transition == 1'b1) ? i_input_data[503 % IN_WIDTH] : pong_storage_data_200 ^ i_input_data[503 % IN_WIDTH];
                743 / IN_WIDTH: pong_storage_data_200 <= (fillup_transition == 1'b1) ? i_input_data[743 % IN_WIDTH] : pong_storage_data_200 ^ i_input_data[743 % IN_WIDTH];
                1064 / IN_WIDTH: pong_storage_data_200 <= (fillup_transition == 1'b1) ? i_input_data[1064 % IN_WIDTH] : pong_storage_data_200 ^ i_input_data[1064 % IN_WIDTH];
                default: pong_storage_data_200 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_200;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_200 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_200;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_200 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_200;
            end
        end
    end
end

logic ping_storage_data_201;
logic pong_storage_data_201;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_201 <= 1'b0;
        pong_storage_data_201 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                369 / IN_WIDTH: ping_storage_data_201 <= (fillup_transition == 1'b1) ? i_input_data[369 % IN_WIDTH] : ping_storage_data_201 ^ i_input_data[369 % IN_WIDTH];
                467 / IN_WIDTH: ping_storage_data_201 <= (fillup_transition == 1'b1) ? i_input_data[467 % IN_WIDTH] : ping_storage_data_201 ^ i_input_data[467 % IN_WIDTH];
                504 / IN_WIDTH: ping_storage_data_201 <= (fillup_transition == 1'b1) ? i_input_data[504 % IN_WIDTH] : ping_storage_data_201 ^ i_input_data[504 % IN_WIDTH];
                744 / IN_WIDTH: ping_storage_data_201 <= (fillup_transition == 1'b1) ? i_input_data[744 % IN_WIDTH] : ping_storage_data_201 ^ i_input_data[744 % IN_WIDTH];
                1065 / IN_WIDTH: ping_storage_data_201 <= (fillup_transition == 1'b1) ? i_input_data[1065 % IN_WIDTH] : ping_storage_data_201 ^ i_input_data[1065 % IN_WIDTH];
                default: ping_storage_data_201 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_201;
                endcase
            end else begin
                case (input_count)
                369 / IN_WIDTH: pong_storage_data_201 <= (fillup_transition == 1'b1) ? i_input_data[369 % IN_WIDTH] : pong_storage_data_201 ^ i_input_data[369 % IN_WIDTH];
                467 / IN_WIDTH: pong_storage_data_201 <= (fillup_transition == 1'b1) ? i_input_data[467 % IN_WIDTH] : pong_storage_data_201 ^ i_input_data[467 % IN_WIDTH];
                504 / IN_WIDTH: pong_storage_data_201 <= (fillup_transition == 1'b1) ? i_input_data[504 % IN_WIDTH] : pong_storage_data_201 ^ i_input_data[504 % IN_WIDTH];
                744 / IN_WIDTH: pong_storage_data_201 <= (fillup_transition == 1'b1) ? i_input_data[744 % IN_WIDTH] : pong_storage_data_201 ^ i_input_data[744 % IN_WIDTH];
                1065 / IN_WIDTH: pong_storage_data_201 <= (fillup_transition == 1'b1) ? i_input_data[1065 % IN_WIDTH] : pong_storage_data_201 ^ i_input_data[1065 % IN_WIDTH];
                default: pong_storage_data_201 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_201;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_201 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_201;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_201 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_201;
            end
        end
    end
end

logic ping_storage_data_202;
logic pong_storage_data_202;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_202 <= 1'b0;
        pong_storage_data_202 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                370 / IN_WIDTH: ping_storage_data_202 <= (fillup_transition == 1'b1) ? i_input_data[370 % IN_WIDTH] : ping_storage_data_202 ^ i_input_data[370 % IN_WIDTH];
                468 / IN_WIDTH: ping_storage_data_202 <= (fillup_transition == 1'b1) ? i_input_data[468 % IN_WIDTH] : ping_storage_data_202 ^ i_input_data[468 % IN_WIDTH];
                505 / IN_WIDTH: ping_storage_data_202 <= (fillup_transition == 1'b1) ? i_input_data[505 % IN_WIDTH] : ping_storage_data_202 ^ i_input_data[505 % IN_WIDTH];
                745 / IN_WIDTH: ping_storage_data_202 <= (fillup_transition == 1'b1) ? i_input_data[745 % IN_WIDTH] : ping_storage_data_202 ^ i_input_data[745 % IN_WIDTH];
                1066 / IN_WIDTH: ping_storage_data_202 <= (fillup_transition == 1'b1) ? i_input_data[1066 % IN_WIDTH] : ping_storage_data_202 ^ i_input_data[1066 % IN_WIDTH];
                default: ping_storage_data_202 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_202;
                endcase
            end else begin
                case (input_count)
                370 / IN_WIDTH: pong_storage_data_202 <= (fillup_transition == 1'b1) ? i_input_data[370 % IN_WIDTH] : pong_storage_data_202 ^ i_input_data[370 % IN_WIDTH];
                468 / IN_WIDTH: pong_storage_data_202 <= (fillup_transition == 1'b1) ? i_input_data[468 % IN_WIDTH] : pong_storage_data_202 ^ i_input_data[468 % IN_WIDTH];
                505 / IN_WIDTH: pong_storage_data_202 <= (fillup_transition == 1'b1) ? i_input_data[505 % IN_WIDTH] : pong_storage_data_202 ^ i_input_data[505 % IN_WIDTH];
                745 / IN_WIDTH: pong_storage_data_202 <= (fillup_transition == 1'b1) ? i_input_data[745 % IN_WIDTH] : pong_storage_data_202 ^ i_input_data[745 % IN_WIDTH];
                1066 / IN_WIDTH: pong_storage_data_202 <= (fillup_transition == 1'b1) ? i_input_data[1066 % IN_WIDTH] : pong_storage_data_202 ^ i_input_data[1066 % IN_WIDTH];
                default: pong_storage_data_202 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_202;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_202 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_202;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_202 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_202;
            end
        end
    end
end

logic ping_storage_data_203;
logic pong_storage_data_203;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_203 <= 1'b0;
        pong_storage_data_203 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                371 / IN_WIDTH: ping_storage_data_203 <= (fillup_transition == 1'b1) ? i_input_data[371 % IN_WIDTH] : ping_storage_data_203 ^ i_input_data[371 % IN_WIDTH];
                469 / IN_WIDTH: ping_storage_data_203 <= (fillup_transition == 1'b1) ? i_input_data[469 % IN_WIDTH] : ping_storage_data_203 ^ i_input_data[469 % IN_WIDTH];
                506 / IN_WIDTH: ping_storage_data_203 <= (fillup_transition == 1'b1) ? i_input_data[506 % IN_WIDTH] : ping_storage_data_203 ^ i_input_data[506 % IN_WIDTH];
                746 / IN_WIDTH: ping_storage_data_203 <= (fillup_transition == 1'b1) ? i_input_data[746 % IN_WIDTH] : ping_storage_data_203 ^ i_input_data[746 % IN_WIDTH];
                1067 / IN_WIDTH: ping_storage_data_203 <= (fillup_transition == 1'b1) ? i_input_data[1067 % IN_WIDTH] : ping_storage_data_203 ^ i_input_data[1067 % IN_WIDTH];
                default: ping_storage_data_203 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_203;
                endcase
            end else begin
                case (input_count)
                371 / IN_WIDTH: pong_storage_data_203 <= (fillup_transition == 1'b1) ? i_input_data[371 % IN_WIDTH] : pong_storage_data_203 ^ i_input_data[371 % IN_WIDTH];
                469 / IN_WIDTH: pong_storage_data_203 <= (fillup_transition == 1'b1) ? i_input_data[469 % IN_WIDTH] : pong_storage_data_203 ^ i_input_data[469 % IN_WIDTH];
                506 / IN_WIDTH: pong_storage_data_203 <= (fillup_transition == 1'b1) ? i_input_data[506 % IN_WIDTH] : pong_storage_data_203 ^ i_input_data[506 % IN_WIDTH];
                746 / IN_WIDTH: pong_storage_data_203 <= (fillup_transition == 1'b1) ? i_input_data[746 % IN_WIDTH] : pong_storage_data_203 ^ i_input_data[746 % IN_WIDTH];
                1067 / IN_WIDTH: pong_storage_data_203 <= (fillup_transition == 1'b1) ? i_input_data[1067 % IN_WIDTH] : pong_storage_data_203 ^ i_input_data[1067 % IN_WIDTH];
                default: pong_storage_data_203 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_203;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_203 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_203;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_203 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_203;
            end
        end
    end
end

logic ping_storage_data_204;
logic pong_storage_data_204;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_204 <= 1'b0;
        pong_storage_data_204 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                372 / IN_WIDTH: ping_storage_data_204 <= (fillup_transition == 1'b1) ? i_input_data[372 % IN_WIDTH] : ping_storage_data_204 ^ i_input_data[372 % IN_WIDTH];
                470 / IN_WIDTH: ping_storage_data_204 <= (fillup_transition == 1'b1) ? i_input_data[470 % IN_WIDTH] : ping_storage_data_204 ^ i_input_data[470 % IN_WIDTH];
                507 / IN_WIDTH: ping_storage_data_204 <= (fillup_transition == 1'b1) ? i_input_data[507 % IN_WIDTH] : ping_storage_data_204 ^ i_input_data[507 % IN_WIDTH];
                747 / IN_WIDTH: ping_storage_data_204 <= (fillup_transition == 1'b1) ? i_input_data[747 % IN_WIDTH] : ping_storage_data_204 ^ i_input_data[747 % IN_WIDTH];
                1068 / IN_WIDTH: ping_storage_data_204 <= (fillup_transition == 1'b1) ? i_input_data[1068 % IN_WIDTH] : ping_storage_data_204 ^ i_input_data[1068 % IN_WIDTH];
                default: ping_storage_data_204 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_204;
                endcase
            end else begin
                case (input_count)
                372 / IN_WIDTH: pong_storage_data_204 <= (fillup_transition == 1'b1) ? i_input_data[372 % IN_WIDTH] : pong_storage_data_204 ^ i_input_data[372 % IN_WIDTH];
                470 / IN_WIDTH: pong_storage_data_204 <= (fillup_transition == 1'b1) ? i_input_data[470 % IN_WIDTH] : pong_storage_data_204 ^ i_input_data[470 % IN_WIDTH];
                507 / IN_WIDTH: pong_storage_data_204 <= (fillup_transition == 1'b1) ? i_input_data[507 % IN_WIDTH] : pong_storage_data_204 ^ i_input_data[507 % IN_WIDTH];
                747 / IN_WIDTH: pong_storage_data_204 <= (fillup_transition == 1'b1) ? i_input_data[747 % IN_WIDTH] : pong_storage_data_204 ^ i_input_data[747 % IN_WIDTH];
                1068 / IN_WIDTH: pong_storage_data_204 <= (fillup_transition == 1'b1) ? i_input_data[1068 % IN_WIDTH] : pong_storage_data_204 ^ i_input_data[1068 % IN_WIDTH];
                default: pong_storage_data_204 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_204;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_204 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_204;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_204 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_204;
            end
        end
    end
end

logic ping_storage_data_205;
logic pong_storage_data_205;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_205 <= 1'b0;
        pong_storage_data_205 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                373 / IN_WIDTH: ping_storage_data_205 <= (fillup_transition == 1'b1) ? i_input_data[373 % IN_WIDTH] : ping_storage_data_205 ^ i_input_data[373 % IN_WIDTH];
                471 / IN_WIDTH: ping_storage_data_205 <= (fillup_transition == 1'b1) ? i_input_data[471 % IN_WIDTH] : ping_storage_data_205 ^ i_input_data[471 % IN_WIDTH];
                508 / IN_WIDTH: ping_storage_data_205 <= (fillup_transition == 1'b1) ? i_input_data[508 % IN_WIDTH] : ping_storage_data_205 ^ i_input_data[508 % IN_WIDTH];
                748 / IN_WIDTH: ping_storage_data_205 <= (fillup_transition == 1'b1) ? i_input_data[748 % IN_WIDTH] : ping_storage_data_205 ^ i_input_data[748 % IN_WIDTH];
                1069 / IN_WIDTH: ping_storage_data_205 <= (fillup_transition == 1'b1) ? i_input_data[1069 % IN_WIDTH] : ping_storage_data_205 ^ i_input_data[1069 % IN_WIDTH];
                default: ping_storage_data_205 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_205;
                endcase
            end else begin
                case (input_count)
                373 / IN_WIDTH: pong_storage_data_205 <= (fillup_transition == 1'b1) ? i_input_data[373 % IN_WIDTH] : pong_storage_data_205 ^ i_input_data[373 % IN_WIDTH];
                471 / IN_WIDTH: pong_storage_data_205 <= (fillup_transition == 1'b1) ? i_input_data[471 % IN_WIDTH] : pong_storage_data_205 ^ i_input_data[471 % IN_WIDTH];
                508 / IN_WIDTH: pong_storage_data_205 <= (fillup_transition == 1'b1) ? i_input_data[508 % IN_WIDTH] : pong_storage_data_205 ^ i_input_data[508 % IN_WIDTH];
                748 / IN_WIDTH: pong_storage_data_205 <= (fillup_transition == 1'b1) ? i_input_data[748 % IN_WIDTH] : pong_storage_data_205 ^ i_input_data[748 % IN_WIDTH];
                1069 / IN_WIDTH: pong_storage_data_205 <= (fillup_transition == 1'b1) ? i_input_data[1069 % IN_WIDTH] : pong_storage_data_205 ^ i_input_data[1069 % IN_WIDTH];
                default: pong_storage_data_205 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_205;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_205 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_205;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_205 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_205;
            end
        end
    end
end

logic ping_storage_data_206;
logic pong_storage_data_206;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_206 <= 1'b0;
        pong_storage_data_206 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                374 / IN_WIDTH: ping_storage_data_206 <= (fillup_transition == 1'b1) ? i_input_data[374 % IN_WIDTH] : ping_storage_data_206 ^ i_input_data[374 % IN_WIDTH];
                472 / IN_WIDTH: ping_storage_data_206 <= (fillup_transition == 1'b1) ? i_input_data[472 % IN_WIDTH] : ping_storage_data_206 ^ i_input_data[472 % IN_WIDTH];
                509 / IN_WIDTH: ping_storage_data_206 <= (fillup_transition == 1'b1) ? i_input_data[509 % IN_WIDTH] : ping_storage_data_206 ^ i_input_data[509 % IN_WIDTH];
                749 / IN_WIDTH: ping_storage_data_206 <= (fillup_transition == 1'b1) ? i_input_data[749 % IN_WIDTH] : ping_storage_data_206 ^ i_input_data[749 % IN_WIDTH];
                1070 / IN_WIDTH: ping_storage_data_206 <= (fillup_transition == 1'b1) ? i_input_data[1070 % IN_WIDTH] : ping_storage_data_206 ^ i_input_data[1070 % IN_WIDTH];
                default: ping_storage_data_206 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_206;
                endcase
            end else begin
                case (input_count)
                374 / IN_WIDTH: pong_storage_data_206 <= (fillup_transition == 1'b1) ? i_input_data[374 % IN_WIDTH] : pong_storage_data_206 ^ i_input_data[374 % IN_WIDTH];
                472 / IN_WIDTH: pong_storage_data_206 <= (fillup_transition == 1'b1) ? i_input_data[472 % IN_WIDTH] : pong_storage_data_206 ^ i_input_data[472 % IN_WIDTH];
                509 / IN_WIDTH: pong_storage_data_206 <= (fillup_transition == 1'b1) ? i_input_data[509 % IN_WIDTH] : pong_storage_data_206 ^ i_input_data[509 % IN_WIDTH];
                749 / IN_WIDTH: pong_storage_data_206 <= (fillup_transition == 1'b1) ? i_input_data[749 % IN_WIDTH] : pong_storage_data_206 ^ i_input_data[749 % IN_WIDTH];
                1070 / IN_WIDTH: pong_storage_data_206 <= (fillup_transition == 1'b1) ? i_input_data[1070 % IN_WIDTH] : pong_storage_data_206 ^ i_input_data[1070 % IN_WIDTH];
                default: pong_storage_data_206 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_206;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_206 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_206;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_206 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_206;
            end
        end
    end
end

logic ping_storage_data_207;
logic pong_storage_data_207;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_207 <= 1'b0;
        pong_storage_data_207 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                375 / IN_WIDTH: ping_storage_data_207 <= (fillup_transition == 1'b1) ? i_input_data[375 % IN_WIDTH] : ping_storage_data_207 ^ i_input_data[375 % IN_WIDTH];
                473 / IN_WIDTH: ping_storage_data_207 <= (fillup_transition == 1'b1) ? i_input_data[473 % IN_WIDTH] : ping_storage_data_207 ^ i_input_data[473 % IN_WIDTH];
                510 / IN_WIDTH: ping_storage_data_207 <= (fillup_transition == 1'b1) ? i_input_data[510 % IN_WIDTH] : ping_storage_data_207 ^ i_input_data[510 % IN_WIDTH];
                750 / IN_WIDTH: ping_storage_data_207 <= (fillup_transition == 1'b1) ? i_input_data[750 % IN_WIDTH] : ping_storage_data_207 ^ i_input_data[750 % IN_WIDTH];
                1071 / IN_WIDTH: ping_storage_data_207 <= (fillup_transition == 1'b1) ? i_input_data[1071 % IN_WIDTH] : ping_storage_data_207 ^ i_input_data[1071 % IN_WIDTH];
                default: ping_storage_data_207 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_207;
                endcase
            end else begin
                case (input_count)
                375 / IN_WIDTH: pong_storage_data_207 <= (fillup_transition == 1'b1) ? i_input_data[375 % IN_WIDTH] : pong_storage_data_207 ^ i_input_data[375 % IN_WIDTH];
                473 / IN_WIDTH: pong_storage_data_207 <= (fillup_transition == 1'b1) ? i_input_data[473 % IN_WIDTH] : pong_storage_data_207 ^ i_input_data[473 % IN_WIDTH];
                510 / IN_WIDTH: pong_storage_data_207 <= (fillup_transition == 1'b1) ? i_input_data[510 % IN_WIDTH] : pong_storage_data_207 ^ i_input_data[510 % IN_WIDTH];
                750 / IN_WIDTH: pong_storage_data_207 <= (fillup_transition == 1'b1) ? i_input_data[750 % IN_WIDTH] : pong_storage_data_207 ^ i_input_data[750 % IN_WIDTH];
                1071 / IN_WIDTH: pong_storage_data_207 <= (fillup_transition == 1'b1) ? i_input_data[1071 % IN_WIDTH] : pong_storage_data_207 ^ i_input_data[1071 % IN_WIDTH];
                default: pong_storage_data_207 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_207;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_207 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_207;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_207 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_207;
            end
        end
    end
end

logic ping_storage_data_208;
logic pong_storage_data_208;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_208 <= 1'b0;
        pong_storage_data_208 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                376 / IN_WIDTH: ping_storage_data_208 <= (fillup_transition == 1'b1) ? i_input_data[376 % IN_WIDTH] : ping_storage_data_208 ^ i_input_data[376 % IN_WIDTH];
                474 / IN_WIDTH: ping_storage_data_208 <= (fillup_transition == 1'b1) ? i_input_data[474 % IN_WIDTH] : ping_storage_data_208 ^ i_input_data[474 % IN_WIDTH];
                511 / IN_WIDTH: ping_storage_data_208 <= (fillup_transition == 1'b1) ? i_input_data[511 % IN_WIDTH] : ping_storage_data_208 ^ i_input_data[511 % IN_WIDTH];
                751 / IN_WIDTH: ping_storage_data_208 <= (fillup_transition == 1'b1) ? i_input_data[751 % IN_WIDTH] : ping_storage_data_208 ^ i_input_data[751 % IN_WIDTH];
                1072 / IN_WIDTH: ping_storage_data_208 <= (fillup_transition == 1'b1) ? i_input_data[1072 % IN_WIDTH] : ping_storage_data_208 ^ i_input_data[1072 % IN_WIDTH];
                default: ping_storage_data_208 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_208;
                endcase
            end else begin
                case (input_count)
                376 / IN_WIDTH: pong_storage_data_208 <= (fillup_transition == 1'b1) ? i_input_data[376 % IN_WIDTH] : pong_storage_data_208 ^ i_input_data[376 % IN_WIDTH];
                474 / IN_WIDTH: pong_storage_data_208 <= (fillup_transition == 1'b1) ? i_input_data[474 % IN_WIDTH] : pong_storage_data_208 ^ i_input_data[474 % IN_WIDTH];
                511 / IN_WIDTH: pong_storage_data_208 <= (fillup_transition == 1'b1) ? i_input_data[511 % IN_WIDTH] : pong_storage_data_208 ^ i_input_data[511 % IN_WIDTH];
                751 / IN_WIDTH: pong_storage_data_208 <= (fillup_transition == 1'b1) ? i_input_data[751 % IN_WIDTH] : pong_storage_data_208 ^ i_input_data[751 % IN_WIDTH];
                1072 / IN_WIDTH: pong_storage_data_208 <= (fillup_transition == 1'b1) ? i_input_data[1072 % IN_WIDTH] : pong_storage_data_208 ^ i_input_data[1072 % IN_WIDTH];
                default: pong_storage_data_208 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_208;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_208 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_208;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_208 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_208;
            end
        end
    end
end

logic ping_storage_data_209;
logic pong_storage_data_209;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_209 <= 1'b0;
        pong_storage_data_209 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                377 / IN_WIDTH: ping_storage_data_209 <= (fillup_transition == 1'b1) ? i_input_data[377 % IN_WIDTH] : ping_storage_data_209 ^ i_input_data[377 % IN_WIDTH];
                475 / IN_WIDTH: ping_storage_data_209 <= (fillup_transition == 1'b1) ? i_input_data[475 % IN_WIDTH] : ping_storage_data_209 ^ i_input_data[475 % IN_WIDTH];
                512 / IN_WIDTH: ping_storage_data_209 <= (fillup_transition == 1'b1) ? i_input_data[512 % IN_WIDTH] : ping_storage_data_209 ^ i_input_data[512 % IN_WIDTH];
                752 / IN_WIDTH: ping_storage_data_209 <= (fillup_transition == 1'b1) ? i_input_data[752 % IN_WIDTH] : ping_storage_data_209 ^ i_input_data[752 % IN_WIDTH];
                1073 / IN_WIDTH: ping_storage_data_209 <= (fillup_transition == 1'b1) ? i_input_data[1073 % IN_WIDTH] : ping_storage_data_209 ^ i_input_data[1073 % IN_WIDTH];
                default: ping_storage_data_209 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_209;
                endcase
            end else begin
                case (input_count)
                377 / IN_WIDTH: pong_storage_data_209 <= (fillup_transition == 1'b1) ? i_input_data[377 % IN_WIDTH] : pong_storage_data_209 ^ i_input_data[377 % IN_WIDTH];
                475 / IN_WIDTH: pong_storage_data_209 <= (fillup_transition == 1'b1) ? i_input_data[475 % IN_WIDTH] : pong_storage_data_209 ^ i_input_data[475 % IN_WIDTH];
                512 / IN_WIDTH: pong_storage_data_209 <= (fillup_transition == 1'b1) ? i_input_data[512 % IN_WIDTH] : pong_storage_data_209 ^ i_input_data[512 % IN_WIDTH];
                752 / IN_WIDTH: pong_storage_data_209 <= (fillup_transition == 1'b1) ? i_input_data[752 % IN_WIDTH] : pong_storage_data_209 ^ i_input_data[752 % IN_WIDTH];
                1073 / IN_WIDTH: pong_storage_data_209 <= (fillup_transition == 1'b1) ? i_input_data[1073 % IN_WIDTH] : pong_storage_data_209 ^ i_input_data[1073 % IN_WIDTH];
                default: pong_storage_data_209 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_209;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_209 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_209;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_209 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_209;
            end
        end
    end
end

logic ping_storage_data_210;
logic pong_storage_data_210;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_210 <= 1'b0;
        pong_storage_data_210 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                378 / IN_WIDTH: ping_storage_data_210 <= (fillup_transition == 1'b1) ? i_input_data[378 % IN_WIDTH] : ping_storage_data_210 ^ i_input_data[378 % IN_WIDTH];
                476 / IN_WIDTH: ping_storage_data_210 <= (fillup_transition == 1'b1) ? i_input_data[476 % IN_WIDTH] : ping_storage_data_210 ^ i_input_data[476 % IN_WIDTH];
                513 / IN_WIDTH: ping_storage_data_210 <= (fillup_transition == 1'b1) ? i_input_data[513 % IN_WIDTH] : ping_storage_data_210 ^ i_input_data[513 % IN_WIDTH];
                753 / IN_WIDTH: ping_storage_data_210 <= (fillup_transition == 1'b1) ? i_input_data[753 % IN_WIDTH] : ping_storage_data_210 ^ i_input_data[753 % IN_WIDTH];
                1074 / IN_WIDTH: ping_storage_data_210 <= (fillup_transition == 1'b1) ? i_input_data[1074 % IN_WIDTH] : ping_storage_data_210 ^ i_input_data[1074 % IN_WIDTH];
                default: ping_storage_data_210 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_210;
                endcase
            end else begin
                case (input_count)
                378 / IN_WIDTH: pong_storage_data_210 <= (fillup_transition == 1'b1) ? i_input_data[378 % IN_WIDTH] : pong_storage_data_210 ^ i_input_data[378 % IN_WIDTH];
                476 / IN_WIDTH: pong_storage_data_210 <= (fillup_transition == 1'b1) ? i_input_data[476 % IN_WIDTH] : pong_storage_data_210 ^ i_input_data[476 % IN_WIDTH];
                513 / IN_WIDTH: pong_storage_data_210 <= (fillup_transition == 1'b1) ? i_input_data[513 % IN_WIDTH] : pong_storage_data_210 ^ i_input_data[513 % IN_WIDTH];
                753 / IN_WIDTH: pong_storage_data_210 <= (fillup_transition == 1'b1) ? i_input_data[753 % IN_WIDTH] : pong_storage_data_210 ^ i_input_data[753 % IN_WIDTH];
                1074 / IN_WIDTH: pong_storage_data_210 <= (fillup_transition == 1'b1) ? i_input_data[1074 % IN_WIDTH] : pong_storage_data_210 ^ i_input_data[1074 % IN_WIDTH];
                default: pong_storage_data_210 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_210;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_210 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_210;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_210 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_210;
            end
        end
    end
end

logic ping_storage_data_211;
logic pong_storage_data_211;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_211 <= 1'b0;
        pong_storage_data_211 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                379 / IN_WIDTH: ping_storage_data_211 <= (fillup_transition == 1'b1) ? i_input_data[379 % IN_WIDTH] : ping_storage_data_211 ^ i_input_data[379 % IN_WIDTH];
                477 / IN_WIDTH: ping_storage_data_211 <= (fillup_transition == 1'b1) ? i_input_data[477 % IN_WIDTH] : ping_storage_data_211 ^ i_input_data[477 % IN_WIDTH];
                514 / IN_WIDTH: ping_storage_data_211 <= (fillup_transition == 1'b1) ? i_input_data[514 % IN_WIDTH] : ping_storage_data_211 ^ i_input_data[514 % IN_WIDTH];
                754 / IN_WIDTH: ping_storage_data_211 <= (fillup_transition == 1'b1) ? i_input_data[754 % IN_WIDTH] : ping_storage_data_211 ^ i_input_data[754 % IN_WIDTH];
                1075 / IN_WIDTH: ping_storage_data_211 <= (fillup_transition == 1'b1) ? i_input_data[1075 % IN_WIDTH] : ping_storage_data_211 ^ i_input_data[1075 % IN_WIDTH];
                default: ping_storage_data_211 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_211;
                endcase
            end else begin
                case (input_count)
                379 / IN_WIDTH: pong_storage_data_211 <= (fillup_transition == 1'b1) ? i_input_data[379 % IN_WIDTH] : pong_storage_data_211 ^ i_input_data[379 % IN_WIDTH];
                477 / IN_WIDTH: pong_storage_data_211 <= (fillup_transition == 1'b1) ? i_input_data[477 % IN_WIDTH] : pong_storage_data_211 ^ i_input_data[477 % IN_WIDTH];
                514 / IN_WIDTH: pong_storage_data_211 <= (fillup_transition == 1'b1) ? i_input_data[514 % IN_WIDTH] : pong_storage_data_211 ^ i_input_data[514 % IN_WIDTH];
                754 / IN_WIDTH: pong_storage_data_211 <= (fillup_transition == 1'b1) ? i_input_data[754 % IN_WIDTH] : pong_storage_data_211 ^ i_input_data[754 % IN_WIDTH];
                1075 / IN_WIDTH: pong_storage_data_211 <= (fillup_transition == 1'b1) ? i_input_data[1075 % IN_WIDTH] : pong_storage_data_211 ^ i_input_data[1075 % IN_WIDTH];
                default: pong_storage_data_211 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_211;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_211 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_211;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_211 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_211;
            end
        end
    end
end

logic ping_storage_data_212;
logic pong_storage_data_212;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_212 <= 1'b0;
        pong_storage_data_212 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                380 / IN_WIDTH: ping_storage_data_212 <= (fillup_transition == 1'b1) ? i_input_data[380 % IN_WIDTH] : ping_storage_data_212 ^ i_input_data[380 % IN_WIDTH];
                478 / IN_WIDTH: ping_storage_data_212 <= (fillup_transition == 1'b1) ? i_input_data[478 % IN_WIDTH] : ping_storage_data_212 ^ i_input_data[478 % IN_WIDTH];
                515 / IN_WIDTH: ping_storage_data_212 <= (fillup_transition == 1'b1) ? i_input_data[515 % IN_WIDTH] : ping_storage_data_212 ^ i_input_data[515 % IN_WIDTH];
                755 / IN_WIDTH: ping_storage_data_212 <= (fillup_transition == 1'b1) ? i_input_data[755 % IN_WIDTH] : ping_storage_data_212 ^ i_input_data[755 % IN_WIDTH];
                1076 / IN_WIDTH: ping_storage_data_212 <= (fillup_transition == 1'b1) ? i_input_data[1076 % IN_WIDTH] : ping_storage_data_212 ^ i_input_data[1076 % IN_WIDTH];
                default: ping_storage_data_212 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_212;
                endcase
            end else begin
                case (input_count)
                380 / IN_WIDTH: pong_storage_data_212 <= (fillup_transition == 1'b1) ? i_input_data[380 % IN_WIDTH] : pong_storage_data_212 ^ i_input_data[380 % IN_WIDTH];
                478 / IN_WIDTH: pong_storage_data_212 <= (fillup_transition == 1'b1) ? i_input_data[478 % IN_WIDTH] : pong_storage_data_212 ^ i_input_data[478 % IN_WIDTH];
                515 / IN_WIDTH: pong_storage_data_212 <= (fillup_transition == 1'b1) ? i_input_data[515 % IN_WIDTH] : pong_storage_data_212 ^ i_input_data[515 % IN_WIDTH];
                755 / IN_WIDTH: pong_storage_data_212 <= (fillup_transition == 1'b1) ? i_input_data[755 % IN_WIDTH] : pong_storage_data_212 ^ i_input_data[755 % IN_WIDTH];
                1076 / IN_WIDTH: pong_storage_data_212 <= (fillup_transition == 1'b1) ? i_input_data[1076 % IN_WIDTH] : pong_storage_data_212 ^ i_input_data[1076 % IN_WIDTH];
                default: pong_storage_data_212 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_212;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_212 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_212;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_212 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_212;
            end
        end
    end
end

logic ping_storage_data_213;
logic pong_storage_data_213;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_213 <= 1'b0;
        pong_storage_data_213 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                381 / IN_WIDTH: ping_storage_data_213 <= (fillup_transition == 1'b1) ? i_input_data[381 % IN_WIDTH] : ping_storage_data_213 ^ i_input_data[381 % IN_WIDTH];
                479 / IN_WIDTH: ping_storage_data_213 <= (fillup_transition == 1'b1) ? i_input_data[479 % IN_WIDTH] : ping_storage_data_213 ^ i_input_data[479 % IN_WIDTH];
                516 / IN_WIDTH: ping_storage_data_213 <= (fillup_transition == 1'b1) ? i_input_data[516 % IN_WIDTH] : ping_storage_data_213 ^ i_input_data[516 % IN_WIDTH];
                756 / IN_WIDTH: ping_storage_data_213 <= (fillup_transition == 1'b1) ? i_input_data[756 % IN_WIDTH] : ping_storage_data_213 ^ i_input_data[756 % IN_WIDTH];
                1077 / IN_WIDTH: ping_storage_data_213 <= (fillup_transition == 1'b1) ? i_input_data[1077 % IN_WIDTH] : ping_storage_data_213 ^ i_input_data[1077 % IN_WIDTH];
                default: ping_storage_data_213 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_213;
                endcase
            end else begin
                case (input_count)
                381 / IN_WIDTH: pong_storage_data_213 <= (fillup_transition == 1'b1) ? i_input_data[381 % IN_WIDTH] : pong_storage_data_213 ^ i_input_data[381 % IN_WIDTH];
                479 / IN_WIDTH: pong_storage_data_213 <= (fillup_transition == 1'b1) ? i_input_data[479 % IN_WIDTH] : pong_storage_data_213 ^ i_input_data[479 % IN_WIDTH];
                516 / IN_WIDTH: pong_storage_data_213 <= (fillup_transition == 1'b1) ? i_input_data[516 % IN_WIDTH] : pong_storage_data_213 ^ i_input_data[516 % IN_WIDTH];
                756 / IN_WIDTH: pong_storage_data_213 <= (fillup_transition == 1'b1) ? i_input_data[756 % IN_WIDTH] : pong_storage_data_213 ^ i_input_data[756 % IN_WIDTH];
                1077 / IN_WIDTH: pong_storage_data_213 <= (fillup_transition == 1'b1) ? i_input_data[1077 % IN_WIDTH] : pong_storage_data_213 ^ i_input_data[1077 % IN_WIDTH];
                default: pong_storage_data_213 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_213;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_213 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_213;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_213 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_213;
            end
        end
    end
end

logic ping_storage_data_214;
logic pong_storage_data_214;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_214 <= 1'b0;
        pong_storage_data_214 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                382 / IN_WIDTH: ping_storage_data_214 <= (fillup_transition == 1'b1) ? i_input_data[382 % IN_WIDTH] : ping_storage_data_214 ^ i_input_data[382 % IN_WIDTH];
                384 / IN_WIDTH: ping_storage_data_214 <= (fillup_transition == 1'b1) ? i_input_data[384 % IN_WIDTH] : ping_storage_data_214 ^ i_input_data[384 % IN_WIDTH];
                517 / IN_WIDTH: ping_storage_data_214 <= (fillup_transition == 1'b1) ? i_input_data[517 % IN_WIDTH] : ping_storage_data_214 ^ i_input_data[517 % IN_WIDTH];
                757 / IN_WIDTH: ping_storage_data_214 <= (fillup_transition == 1'b1) ? i_input_data[757 % IN_WIDTH] : ping_storage_data_214 ^ i_input_data[757 % IN_WIDTH];
                1078 / IN_WIDTH: ping_storage_data_214 <= (fillup_transition == 1'b1) ? i_input_data[1078 % IN_WIDTH] : ping_storage_data_214 ^ i_input_data[1078 % IN_WIDTH];
                default: ping_storage_data_214 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_214;
                endcase
            end else begin
                case (input_count)
                382 / IN_WIDTH: pong_storage_data_214 <= (fillup_transition == 1'b1) ? i_input_data[382 % IN_WIDTH] : pong_storage_data_214 ^ i_input_data[382 % IN_WIDTH];
                384 / IN_WIDTH: pong_storage_data_214 <= (fillup_transition == 1'b1) ? i_input_data[384 % IN_WIDTH] : pong_storage_data_214 ^ i_input_data[384 % IN_WIDTH];
                517 / IN_WIDTH: pong_storage_data_214 <= (fillup_transition == 1'b1) ? i_input_data[517 % IN_WIDTH] : pong_storage_data_214 ^ i_input_data[517 % IN_WIDTH];
                757 / IN_WIDTH: pong_storage_data_214 <= (fillup_transition == 1'b1) ? i_input_data[757 % IN_WIDTH] : pong_storage_data_214 ^ i_input_data[757 % IN_WIDTH];
                1078 / IN_WIDTH: pong_storage_data_214 <= (fillup_transition == 1'b1) ? i_input_data[1078 % IN_WIDTH] : pong_storage_data_214 ^ i_input_data[1078 % IN_WIDTH];
                default: pong_storage_data_214 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_214;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_214 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_214;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_214 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_214;
            end
        end
    end
end

logic ping_storage_data_215;
logic pong_storage_data_215;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_215 <= 1'b0;
        pong_storage_data_215 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                383 / IN_WIDTH: ping_storage_data_215 <= (fillup_transition == 1'b1) ? i_input_data[383 % IN_WIDTH] : ping_storage_data_215 ^ i_input_data[383 % IN_WIDTH];
                385 / IN_WIDTH: ping_storage_data_215 <= (fillup_transition == 1'b1) ? i_input_data[385 % IN_WIDTH] : ping_storage_data_215 ^ i_input_data[385 % IN_WIDTH];
                518 / IN_WIDTH: ping_storage_data_215 <= (fillup_transition == 1'b1) ? i_input_data[518 % IN_WIDTH] : ping_storage_data_215 ^ i_input_data[518 % IN_WIDTH];
                758 / IN_WIDTH: ping_storage_data_215 <= (fillup_transition == 1'b1) ? i_input_data[758 % IN_WIDTH] : ping_storage_data_215 ^ i_input_data[758 % IN_WIDTH];
                1079 / IN_WIDTH: ping_storage_data_215 <= (fillup_transition == 1'b1) ? i_input_data[1079 % IN_WIDTH] : ping_storage_data_215 ^ i_input_data[1079 % IN_WIDTH];
                default: ping_storage_data_215 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_215;
                endcase
            end else begin
                case (input_count)
                383 / IN_WIDTH: pong_storage_data_215 <= (fillup_transition == 1'b1) ? i_input_data[383 % IN_WIDTH] : pong_storage_data_215 ^ i_input_data[383 % IN_WIDTH];
                385 / IN_WIDTH: pong_storage_data_215 <= (fillup_transition == 1'b1) ? i_input_data[385 % IN_WIDTH] : pong_storage_data_215 ^ i_input_data[385 % IN_WIDTH];
                518 / IN_WIDTH: pong_storage_data_215 <= (fillup_transition == 1'b1) ? i_input_data[518 % IN_WIDTH] : pong_storage_data_215 ^ i_input_data[518 % IN_WIDTH];
                758 / IN_WIDTH: pong_storage_data_215 <= (fillup_transition == 1'b1) ? i_input_data[758 % IN_WIDTH] : pong_storage_data_215 ^ i_input_data[758 % IN_WIDTH];
                1079 / IN_WIDTH: pong_storage_data_215 <= (fillup_transition == 1'b1) ? i_input_data[1079 % IN_WIDTH] : pong_storage_data_215 ^ i_input_data[1079 % IN_WIDTH];
                default: pong_storage_data_215 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_215;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_215 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_215;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_215 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_215;
            end
        end
    end
end

logic ping_storage_data_216;
logic pong_storage_data_216;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_216 <= 1'b0;
        pong_storage_data_216 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                288 / IN_WIDTH: ping_storage_data_216 <= (fillup_transition == 1'b1) ? i_input_data[288 % IN_WIDTH] : ping_storage_data_216 ^ i_input_data[288 % IN_WIDTH];
                386 / IN_WIDTH: ping_storage_data_216 <= (fillup_transition == 1'b1) ? i_input_data[386 % IN_WIDTH] : ping_storage_data_216 ^ i_input_data[386 % IN_WIDTH];
                519 / IN_WIDTH: ping_storage_data_216 <= (fillup_transition == 1'b1) ? i_input_data[519 % IN_WIDTH] : ping_storage_data_216 ^ i_input_data[519 % IN_WIDTH];
                759 / IN_WIDTH: ping_storage_data_216 <= (fillup_transition == 1'b1) ? i_input_data[759 % IN_WIDTH] : ping_storage_data_216 ^ i_input_data[759 % IN_WIDTH];
                1080 / IN_WIDTH: ping_storage_data_216 <= (fillup_transition == 1'b1) ? i_input_data[1080 % IN_WIDTH] : ping_storage_data_216 ^ i_input_data[1080 % IN_WIDTH];
                default: ping_storage_data_216 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_216;
                endcase
            end else begin
                case (input_count)
                288 / IN_WIDTH: pong_storage_data_216 <= (fillup_transition == 1'b1) ? i_input_data[288 % IN_WIDTH] : pong_storage_data_216 ^ i_input_data[288 % IN_WIDTH];
                386 / IN_WIDTH: pong_storage_data_216 <= (fillup_transition == 1'b1) ? i_input_data[386 % IN_WIDTH] : pong_storage_data_216 ^ i_input_data[386 % IN_WIDTH];
                519 / IN_WIDTH: pong_storage_data_216 <= (fillup_transition == 1'b1) ? i_input_data[519 % IN_WIDTH] : pong_storage_data_216 ^ i_input_data[519 % IN_WIDTH];
                759 / IN_WIDTH: pong_storage_data_216 <= (fillup_transition == 1'b1) ? i_input_data[759 % IN_WIDTH] : pong_storage_data_216 ^ i_input_data[759 % IN_WIDTH];
                1080 / IN_WIDTH: pong_storage_data_216 <= (fillup_transition == 1'b1) ? i_input_data[1080 % IN_WIDTH] : pong_storage_data_216 ^ i_input_data[1080 % IN_WIDTH];
                default: pong_storage_data_216 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_216;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_216 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_216;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_216 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_216;
            end
        end
    end
end

logic ping_storage_data_217;
logic pong_storage_data_217;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_217 <= 1'b0;
        pong_storage_data_217 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                289 / IN_WIDTH: ping_storage_data_217 <= (fillup_transition == 1'b1) ? i_input_data[289 % IN_WIDTH] : ping_storage_data_217 ^ i_input_data[289 % IN_WIDTH];
                387 / IN_WIDTH: ping_storage_data_217 <= (fillup_transition == 1'b1) ? i_input_data[387 % IN_WIDTH] : ping_storage_data_217 ^ i_input_data[387 % IN_WIDTH];
                520 / IN_WIDTH: ping_storage_data_217 <= (fillup_transition == 1'b1) ? i_input_data[520 % IN_WIDTH] : ping_storage_data_217 ^ i_input_data[520 % IN_WIDTH];
                760 / IN_WIDTH: ping_storage_data_217 <= (fillup_transition == 1'b1) ? i_input_data[760 % IN_WIDTH] : ping_storage_data_217 ^ i_input_data[760 % IN_WIDTH];
                1081 / IN_WIDTH: ping_storage_data_217 <= (fillup_transition == 1'b1) ? i_input_data[1081 % IN_WIDTH] : ping_storage_data_217 ^ i_input_data[1081 % IN_WIDTH];
                default: ping_storage_data_217 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_217;
                endcase
            end else begin
                case (input_count)
                289 / IN_WIDTH: pong_storage_data_217 <= (fillup_transition == 1'b1) ? i_input_data[289 % IN_WIDTH] : pong_storage_data_217 ^ i_input_data[289 % IN_WIDTH];
                387 / IN_WIDTH: pong_storage_data_217 <= (fillup_transition == 1'b1) ? i_input_data[387 % IN_WIDTH] : pong_storage_data_217 ^ i_input_data[387 % IN_WIDTH];
                520 / IN_WIDTH: pong_storage_data_217 <= (fillup_transition == 1'b1) ? i_input_data[520 % IN_WIDTH] : pong_storage_data_217 ^ i_input_data[520 % IN_WIDTH];
                760 / IN_WIDTH: pong_storage_data_217 <= (fillup_transition == 1'b1) ? i_input_data[760 % IN_WIDTH] : pong_storage_data_217 ^ i_input_data[760 % IN_WIDTH];
                1081 / IN_WIDTH: pong_storage_data_217 <= (fillup_transition == 1'b1) ? i_input_data[1081 % IN_WIDTH] : pong_storage_data_217 ^ i_input_data[1081 % IN_WIDTH];
                default: pong_storage_data_217 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_217;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_217 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_217;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_217 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_217;
            end
        end
    end
end

logic ping_storage_data_218;
logic pong_storage_data_218;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_218 <= 1'b0;
        pong_storage_data_218 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                290 / IN_WIDTH: ping_storage_data_218 <= (fillup_transition == 1'b1) ? i_input_data[290 % IN_WIDTH] : ping_storage_data_218 ^ i_input_data[290 % IN_WIDTH];
                388 / IN_WIDTH: ping_storage_data_218 <= (fillup_transition == 1'b1) ? i_input_data[388 % IN_WIDTH] : ping_storage_data_218 ^ i_input_data[388 % IN_WIDTH];
                521 / IN_WIDTH: ping_storage_data_218 <= (fillup_transition == 1'b1) ? i_input_data[521 % IN_WIDTH] : ping_storage_data_218 ^ i_input_data[521 % IN_WIDTH];
                761 / IN_WIDTH: ping_storage_data_218 <= (fillup_transition == 1'b1) ? i_input_data[761 % IN_WIDTH] : ping_storage_data_218 ^ i_input_data[761 % IN_WIDTH];
                1082 / IN_WIDTH: ping_storage_data_218 <= (fillup_transition == 1'b1) ? i_input_data[1082 % IN_WIDTH] : ping_storage_data_218 ^ i_input_data[1082 % IN_WIDTH];
                default: ping_storage_data_218 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_218;
                endcase
            end else begin
                case (input_count)
                290 / IN_WIDTH: pong_storage_data_218 <= (fillup_transition == 1'b1) ? i_input_data[290 % IN_WIDTH] : pong_storage_data_218 ^ i_input_data[290 % IN_WIDTH];
                388 / IN_WIDTH: pong_storage_data_218 <= (fillup_transition == 1'b1) ? i_input_data[388 % IN_WIDTH] : pong_storage_data_218 ^ i_input_data[388 % IN_WIDTH];
                521 / IN_WIDTH: pong_storage_data_218 <= (fillup_transition == 1'b1) ? i_input_data[521 % IN_WIDTH] : pong_storage_data_218 ^ i_input_data[521 % IN_WIDTH];
                761 / IN_WIDTH: pong_storage_data_218 <= (fillup_transition == 1'b1) ? i_input_data[761 % IN_WIDTH] : pong_storage_data_218 ^ i_input_data[761 % IN_WIDTH];
                1082 / IN_WIDTH: pong_storage_data_218 <= (fillup_transition == 1'b1) ? i_input_data[1082 % IN_WIDTH] : pong_storage_data_218 ^ i_input_data[1082 % IN_WIDTH];
                default: pong_storage_data_218 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_218;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_218 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_218;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_218 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_218;
            end
        end
    end
end

logic ping_storage_data_219;
logic pong_storage_data_219;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_219 <= 1'b0;
        pong_storage_data_219 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                291 / IN_WIDTH: ping_storage_data_219 <= (fillup_transition == 1'b1) ? i_input_data[291 % IN_WIDTH] : ping_storage_data_219 ^ i_input_data[291 % IN_WIDTH];
                389 / IN_WIDTH: ping_storage_data_219 <= (fillup_transition == 1'b1) ? i_input_data[389 % IN_WIDTH] : ping_storage_data_219 ^ i_input_data[389 % IN_WIDTH];
                522 / IN_WIDTH: ping_storage_data_219 <= (fillup_transition == 1'b1) ? i_input_data[522 % IN_WIDTH] : ping_storage_data_219 ^ i_input_data[522 % IN_WIDTH];
                762 / IN_WIDTH: ping_storage_data_219 <= (fillup_transition == 1'b1) ? i_input_data[762 % IN_WIDTH] : ping_storage_data_219 ^ i_input_data[762 % IN_WIDTH];
                1083 / IN_WIDTH: ping_storage_data_219 <= (fillup_transition == 1'b1) ? i_input_data[1083 % IN_WIDTH] : ping_storage_data_219 ^ i_input_data[1083 % IN_WIDTH];
                default: ping_storage_data_219 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_219;
                endcase
            end else begin
                case (input_count)
                291 / IN_WIDTH: pong_storage_data_219 <= (fillup_transition == 1'b1) ? i_input_data[291 % IN_WIDTH] : pong_storage_data_219 ^ i_input_data[291 % IN_WIDTH];
                389 / IN_WIDTH: pong_storage_data_219 <= (fillup_transition == 1'b1) ? i_input_data[389 % IN_WIDTH] : pong_storage_data_219 ^ i_input_data[389 % IN_WIDTH];
                522 / IN_WIDTH: pong_storage_data_219 <= (fillup_transition == 1'b1) ? i_input_data[522 % IN_WIDTH] : pong_storage_data_219 ^ i_input_data[522 % IN_WIDTH];
                762 / IN_WIDTH: pong_storage_data_219 <= (fillup_transition == 1'b1) ? i_input_data[762 % IN_WIDTH] : pong_storage_data_219 ^ i_input_data[762 % IN_WIDTH];
                1083 / IN_WIDTH: pong_storage_data_219 <= (fillup_transition == 1'b1) ? i_input_data[1083 % IN_WIDTH] : pong_storage_data_219 ^ i_input_data[1083 % IN_WIDTH];
                default: pong_storage_data_219 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_219;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_219 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_219;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_219 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_219;
            end
        end
    end
end

logic ping_storage_data_220;
logic pong_storage_data_220;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_220 <= 1'b0;
        pong_storage_data_220 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                292 / IN_WIDTH: ping_storage_data_220 <= (fillup_transition == 1'b1) ? i_input_data[292 % IN_WIDTH] : ping_storage_data_220 ^ i_input_data[292 % IN_WIDTH];
                390 / IN_WIDTH: ping_storage_data_220 <= (fillup_transition == 1'b1) ? i_input_data[390 % IN_WIDTH] : ping_storage_data_220 ^ i_input_data[390 % IN_WIDTH];
                523 / IN_WIDTH: ping_storage_data_220 <= (fillup_transition == 1'b1) ? i_input_data[523 % IN_WIDTH] : ping_storage_data_220 ^ i_input_data[523 % IN_WIDTH];
                763 / IN_WIDTH: ping_storage_data_220 <= (fillup_transition == 1'b1) ? i_input_data[763 % IN_WIDTH] : ping_storage_data_220 ^ i_input_data[763 % IN_WIDTH];
                1084 / IN_WIDTH: ping_storage_data_220 <= (fillup_transition == 1'b1) ? i_input_data[1084 % IN_WIDTH] : ping_storage_data_220 ^ i_input_data[1084 % IN_WIDTH];
                default: ping_storage_data_220 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_220;
                endcase
            end else begin
                case (input_count)
                292 / IN_WIDTH: pong_storage_data_220 <= (fillup_transition == 1'b1) ? i_input_data[292 % IN_WIDTH] : pong_storage_data_220 ^ i_input_data[292 % IN_WIDTH];
                390 / IN_WIDTH: pong_storage_data_220 <= (fillup_transition == 1'b1) ? i_input_data[390 % IN_WIDTH] : pong_storage_data_220 ^ i_input_data[390 % IN_WIDTH];
                523 / IN_WIDTH: pong_storage_data_220 <= (fillup_transition == 1'b1) ? i_input_data[523 % IN_WIDTH] : pong_storage_data_220 ^ i_input_data[523 % IN_WIDTH];
                763 / IN_WIDTH: pong_storage_data_220 <= (fillup_transition == 1'b1) ? i_input_data[763 % IN_WIDTH] : pong_storage_data_220 ^ i_input_data[763 % IN_WIDTH];
                1084 / IN_WIDTH: pong_storage_data_220 <= (fillup_transition == 1'b1) ? i_input_data[1084 % IN_WIDTH] : pong_storage_data_220 ^ i_input_data[1084 % IN_WIDTH];
                default: pong_storage_data_220 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_220;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_220 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_220;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_220 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_220;
            end
        end
    end
end

logic ping_storage_data_221;
logic pong_storage_data_221;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_221 <= 1'b0;
        pong_storage_data_221 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                293 / IN_WIDTH: ping_storage_data_221 <= (fillup_transition == 1'b1) ? i_input_data[293 % IN_WIDTH] : ping_storage_data_221 ^ i_input_data[293 % IN_WIDTH];
                391 / IN_WIDTH: ping_storage_data_221 <= (fillup_transition == 1'b1) ? i_input_data[391 % IN_WIDTH] : ping_storage_data_221 ^ i_input_data[391 % IN_WIDTH];
                524 / IN_WIDTH: ping_storage_data_221 <= (fillup_transition == 1'b1) ? i_input_data[524 % IN_WIDTH] : ping_storage_data_221 ^ i_input_data[524 % IN_WIDTH];
                764 / IN_WIDTH: ping_storage_data_221 <= (fillup_transition == 1'b1) ? i_input_data[764 % IN_WIDTH] : ping_storage_data_221 ^ i_input_data[764 % IN_WIDTH];
                1085 / IN_WIDTH: ping_storage_data_221 <= (fillup_transition == 1'b1) ? i_input_data[1085 % IN_WIDTH] : ping_storage_data_221 ^ i_input_data[1085 % IN_WIDTH];
                default: ping_storage_data_221 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_221;
                endcase
            end else begin
                case (input_count)
                293 / IN_WIDTH: pong_storage_data_221 <= (fillup_transition == 1'b1) ? i_input_data[293 % IN_WIDTH] : pong_storage_data_221 ^ i_input_data[293 % IN_WIDTH];
                391 / IN_WIDTH: pong_storage_data_221 <= (fillup_transition == 1'b1) ? i_input_data[391 % IN_WIDTH] : pong_storage_data_221 ^ i_input_data[391 % IN_WIDTH];
                524 / IN_WIDTH: pong_storage_data_221 <= (fillup_transition == 1'b1) ? i_input_data[524 % IN_WIDTH] : pong_storage_data_221 ^ i_input_data[524 % IN_WIDTH];
                764 / IN_WIDTH: pong_storage_data_221 <= (fillup_transition == 1'b1) ? i_input_data[764 % IN_WIDTH] : pong_storage_data_221 ^ i_input_data[764 % IN_WIDTH];
                1085 / IN_WIDTH: pong_storage_data_221 <= (fillup_transition == 1'b1) ? i_input_data[1085 % IN_WIDTH] : pong_storage_data_221 ^ i_input_data[1085 % IN_WIDTH];
                default: pong_storage_data_221 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_221;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_221 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_221;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_221 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_221;
            end
        end
    end
end

logic ping_storage_data_222;
logic pong_storage_data_222;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_222 <= 1'b0;
        pong_storage_data_222 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                294 / IN_WIDTH: ping_storage_data_222 <= (fillup_transition == 1'b1) ? i_input_data[294 % IN_WIDTH] : ping_storage_data_222 ^ i_input_data[294 % IN_WIDTH];
                392 / IN_WIDTH: ping_storage_data_222 <= (fillup_transition == 1'b1) ? i_input_data[392 % IN_WIDTH] : ping_storage_data_222 ^ i_input_data[392 % IN_WIDTH];
                525 / IN_WIDTH: ping_storage_data_222 <= (fillup_transition == 1'b1) ? i_input_data[525 % IN_WIDTH] : ping_storage_data_222 ^ i_input_data[525 % IN_WIDTH];
                765 / IN_WIDTH: ping_storage_data_222 <= (fillup_transition == 1'b1) ? i_input_data[765 % IN_WIDTH] : ping_storage_data_222 ^ i_input_data[765 % IN_WIDTH];
                1086 / IN_WIDTH: ping_storage_data_222 <= (fillup_transition == 1'b1) ? i_input_data[1086 % IN_WIDTH] : ping_storage_data_222 ^ i_input_data[1086 % IN_WIDTH];
                default: ping_storage_data_222 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_222;
                endcase
            end else begin
                case (input_count)
                294 / IN_WIDTH: pong_storage_data_222 <= (fillup_transition == 1'b1) ? i_input_data[294 % IN_WIDTH] : pong_storage_data_222 ^ i_input_data[294 % IN_WIDTH];
                392 / IN_WIDTH: pong_storage_data_222 <= (fillup_transition == 1'b1) ? i_input_data[392 % IN_WIDTH] : pong_storage_data_222 ^ i_input_data[392 % IN_WIDTH];
                525 / IN_WIDTH: pong_storage_data_222 <= (fillup_transition == 1'b1) ? i_input_data[525 % IN_WIDTH] : pong_storage_data_222 ^ i_input_data[525 % IN_WIDTH];
                765 / IN_WIDTH: pong_storage_data_222 <= (fillup_transition == 1'b1) ? i_input_data[765 % IN_WIDTH] : pong_storage_data_222 ^ i_input_data[765 % IN_WIDTH];
                1086 / IN_WIDTH: pong_storage_data_222 <= (fillup_transition == 1'b1) ? i_input_data[1086 % IN_WIDTH] : pong_storage_data_222 ^ i_input_data[1086 % IN_WIDTH];
                default: pong_storage_data_222 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_222;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_222 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_222;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_222 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_222;
            end
        end
    end
end

logic ping_storage_data_223;
logic pong_storage_data_223;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_223 <= 1'b0;
        pong_storage_data_223 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                295 / IN_WIDTH: ping_storage_data_223 <= (fillup_transition == 1'b1) ? i_input_data[295 % IN_WIDTH] : ping_storage_data_223 ^ i_input_data[295 % IN_WIDTH];
                393 / IN_WIDTH: ping_storage_data_223 <= (fillup_transition == 1'b1) ? i_input_data[393 % IN_WIDTH] : ping_storage_data_223 ^ i_input_data[393 % IN_WIDTH];
                526 / IN_WIDTH: ping_storage_data_223 <= (fillup_transition == 1'b1) ? i_input_data[526 % IN_WIDTH] : ping_storage_data_223 ^ i_input_data[526 % IN_WIDTH];
                766 / IN_WIDTH: ping_storage_data_223 <= (fillup_transition == 1'b1) ? i_input_data[766 % IN_WIDTH] : ping_storage_data_223 ^ i_input_data[766 % IN_WIDTH];
                1087 / IN_WIDTH: ping_storage_data_223 <= (fillup_transition == 1'b1) ? i_input_data[1087 % IN_WIDTH] : ping_storage_data_223 ^ i_input_data[1087 % IN_WIDTH];
                default: ping_storage_data_223 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_223;
                endcase
            end else begin
                case (input_count)
                295 / IN_WIDTH: pong_storage_data_223 <= (fillup_transition == 1'b1) ? i_input_data[295 % IN_WIDTH] : pong_storage_data_223 ^ i_input_data[295 % IN_WIDTH];
                393 / IN_WIDTH: pong_storage_data_223 <= (fillup_transition == 1'b1) ? i_input_data[393 % IN_WIDTH] : pong_storage_data_223 ^ i_input_data[393 % IN_WIDTH];
                526 / IN_WIDTH: pong_storage_data_223 <= (fillup_transition == 1'b1) ? i_input_data[526 % IN_WIDTH] : pong_storage_data_223 ^ i_input_data[526 % IN_WIDTH];
                766 / IN_WIDTH: pong_storage_data_223 <= (fillup_transition == 1'b1) ? i_input_data[766 % IN_WIDTH] : pong_storage_data_223 ^ i_input_data[766 % IN_WIDTH];
                1087 / IN_WIDTH: pong_storage_data_223 <= (fillup_transition == 1'b1) ? i_input_data[1087 % IN_WIDTH] : pong_storage_data_223 ^ i_input_data[1087 % IN_WIDTH];
                default: pong_storage_data_223 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_223;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_223 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_223;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_223 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_223;
            end
        end
    end
end

logic ping_storage_data_224;
logic pong_storage_data_224;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_224 <= 1'b0;
        pong_storage_data_224 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                296 / IN_WIDTH: ping_storage_data_224 <= (fillup_transition == 1'b1) ? i_input_data[296 % IN_WIDTH] : ping_storage_data_224 ^ i_input_data[296 % IN_WIDTH];
                394 / IN_WIDTH: ping_storage_data_224 <= (fillup_transition == 1'b1) ? i_input_data[394 % IN_WIDTH] : ping_storage_data_224 ^ i_input_data[394 % IN_WIDTH];
                527 / IN_WIDTH: ping_storage_data_224 <= (fillup_transition == 1'b1) ? i_input_data[527 % IN_WIDTH] : ping_storage_data_224 ^ i_input_data[527 % IN_WIDTH];
                767 / IN_WIDTH: ping_storage_data_224 <= (fillup_transition == 1'b1) ? i_input_data[767 % IN_WIDTH] : ping_storage_data_224 ^ i_input_data[767 % IN_WIDTH];
                1088 / IN_WIDTH: ping_storage_data_224 <= (fillup_transition == 1'b1) ? i_input_data[1088 % IN_WIDTH] : ping_storage_data_224 ^ i_input_data[1088 % IN_WIDTH];
                default: ping_storage_data_224 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_224;
                endcase
            end else begin
                case (input_count)
                296 / IN_WIDTH: pong_storage_data_224 <= (fillup_transition == 1'b1) ? i_input_data[296 % IN_WIDTH] : pong_storage_data_224 ^ i_input_data[296 % IN_WIDTH];
                394 / IN_WIDTH: pong_storage_data_224 <= (fillup_transition == 1'b1) ? i_input_data[394 % IN_WIDTH] : pong_storage_data_224 ^ i_input_data[394 % IN_WIDTH];
                527 / IN_WIDTH: pong_storage_data_224 <= (fillup_transition == 1'b1) ? i_input_data[527 % IN_WIDTH] : pong_storage_data_224 ^ i_input_data[527 % IN_WIDTH];
                767 / IN_WIDTH: pong_storage_data_224 <= (fillup_transition == 1'b1) ? i_input_data[767 % IN_WIDTH] : pong_storage_data_224 ^ i_input_data[767 % IN_WIDTH];
                1088 / IN_WIDTH: pong_storage_data_224 <= (fillup_transition == 1'b1) ? i_input_data[1088 % IN_WIDTH] : pong_storage_data_224 ^ i_input_data[1088 % IN_WIDTH];
                default: pong_storage_data_224 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_224;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_224 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_224;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_224 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_224;
            end
        end
    end
end

logic ping_storage_data_225;
logic pong_storage_data_225;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_225 <= 1'b0;
        pong_storage_data_225 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                297 / IN_WIDTH: ping_storage_data_225 <= (fillup_transition == 1'b1) ? i_input_data[297 % IN_WIDTH] : ping_storage_data_225 ^ i_input_data[297 % IN_WIDTH];
                395 / IN_WIDTH: ping_storage_data_225 <= (fillup_transition == 1'b1) ? i_input_data[395 % IN_WIDTH] : ping_storage_data_225 ^ i_input_data[395 % IN_WIDTH];
                528 / IN_WIDTH: ping_storage_data_225 <= (fillup_transition == 1'b1) ? i_input_data[528 % IN_WIDTH] : ping_storage_data_225 ^ i_input_data[528 % IN_WIDTH];
                672 / IN_WIDTH: ping_storage_data_225 <= (fillup_transition == 1'b1) ? i_input_data[672 % IN_WIDTH] : ping_storage_data_225 ^ i_input_data[672 % IN_WIDTH];
                1089 / IN_WIDTH: ping_storage_data_225 <= (fillup_transition == 1'b1) ? i_input_data[1089 % IN_WIDTH] : ping_storage_data_225 ^ i_input_data[1089 % IN_WIDTH];
                default: ping_storage_data_225 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_225;
                endcase
            end else begin
                case (input_count)
                297 / IN_WIDTH: pong_storage_data_225 <= (fillup_transition == 1'b1) ? i_input_data[297 % IN_WIDTH] : pong_storage_data_225 ^ i_input_data[297 % IN_WIDTH];
                395 / IN_WIDTH: pong_storage_data_225 <= (fillup_transition == 1'b1) ? i_input_data[395 % IN_WIDTH] : pong_storage_data_225 ^ i_input_data[395 % IN_WIDTH];
                528 / IN_WIDTH: pong_storage_data_225 <= (fillup_transition == 1'b1) ? i_input_data[528 % IN_WIDTH] : pong_storage_data_225 ^ i_input_data[528 % IN_WIDTH];
                672 / IN_WIDTH: pong_storage_data_225 <= (fillup_transition == 1'b1) ? i_input_data[672 % IN_WIDTH] : pong_storage_data_225 ^ i_input_data[672 % IN_WIDTH];
                1089 / IN_WIDTH: pong_storage_data_225 <= (fillup_transition == 1'b1) ? i_input_data[1089 % IN_WIDTH] : pong_storage_data_225 ^ i_input_data[1089 % IN_WIDTH];
                default: pong_storage_data_225 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_225;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_225 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_225;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_225 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_225;
            end
        end
    end
end

logic ping_storage_data_226;
logic pong_storage_data_226;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_226 <= 1'b0;
        pong_storage_data_226 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                298 / IN_WIDTH: ping_storage_data_226 <= (fillup_transition == 1'b1) ? i_input_data[298 % IN_WIDTH] : ping_storage_data_226 ^ i_input_data[298 % IN_WIDTH];
                396 / IN_WIDTH: ping_storage_data_226 <= (fillup_transition == 1'b1) ? i_input_data[396 % IN_WIDTH] : ping_storage_data_226 ^ i_input_data[396 % IN_WIDTH];
                529 / IN_WIDTH: ping_storage_data_226 <= (fillup_transition == 1'b1) ? i_input_data[529 % IN_WIDTH] : ping_storage_data_226 ^ i_input_data[529 % IN_WIDTH];
                673 / IN_WIDTH: ping_storage_data_226 <= (fillup_transition == 1'b1) ? i_input_data[673 % IN_WIDTH] : ping_storage_data_226 ^ i_input_data[673 % IN_WIDTH];
                1090 / IN_WIDTH: ping_storage_data_226 <= (fillup_transition == 1'b1) ? i_input_data[1090 % IN_WIDTH] : ping_storage_data_226 ^ i_input_data[1090 % IN_WIDTH];
                default: ping_storage_data_226 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_226;
                endcase
            end else begin
                case (input_count)
                298 / IN_WIDTH: pong_storage_data_226 <= (fillup_transition == 1'b1) ? i_input_data[298 % IN_WIDTH] : pong_storage_data_226 ^ i_input_data[298 % IN_WIDTH];
                396 / IN_WIDTH: pong_storage_data_226 <= (fillup_transition == 1'b1) ? i_input_data[396 % IN_WIDTH] : pong_storage_data_226 ^ i_input_data[396 % IN_WIDTH];
                529 / IN_WIDTH: pong_storage_data_226 <= (fillup_transition == 1'b1) ? i_input_data[529 % IN_WIDTH] : pong_storage_data_226 ^ i_input_data[529 % IN_WIDTH];
                673 / IN_WIDTH: pong_storage_data_226 <= (fillup_transition == 1'b1) ? i_input_data[673 % IN_WIDTH] : pong_storage_data_226 ^ i_input_data[673 % IN_WIDTH];
                1090 / IN_WIDTH: pong_storage_data_226 <= (fillup_transition == 1'b1) ? i_input_data[1090 % IN_WIDTH] : pong_storage_data_226 ^ i_input_data[1090 % IN_WIDTH];
                default: pong_storage_data_226 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_226;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_226 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_226;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_226 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_226;
            end
        end
    end
end

logic ping_storage_data_227;
logic pong_storage_data_227;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_227 <= 1'b0;
        pong_storage_data_227 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                299 / IN_WIDTH: ping_storage_data_227 <= (fillup_transition == 1'b1) ? i_input_data[299 % IN_WIDTH] : ping_storage_data_227 ^ i_input_data[299 % IN_WIDTH];
                397 / IN_WIDTH: ping_storage_data_227 <= (fillup_transition == 1'b1) ? i_input_data[397 % IN_WIDTH] : ping_storage_data_227 ^ i_input_data[397 % IN_WIDTH];
                530 / IN_WIDTH: ping_storage_data_227 <= (fillup_transition == 1'b1) ? i_input_data[530 % IN_WIDTH] : ping_storage_data_227 ^ i_input_data[530 % IN_WIDTH];
                674 / IN_WIDTH: ping_storage_data_227 <= (fillup_transition == 1'b1) ? i_input_data[674 % IN_WIDTH] : ping_storage_data_227 ^ i_input_data[674 % IN_WIDTH];
                1091 / IN_WIDTH: ping_storage_data_227 <= (fillup_transition == 1'b1) ? i_input_data[1091 % IN_WIDTH] : ping_storage_data_227 ^ i_input_data[1091 % IN_WIDTH];
                default: ping_storage_data_227 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_227;
                endcase
            end else begin
                case (input_count)
                299 / IN_WIDTH: pong_storage_data_227 <= (fillup_transition == 1'b1) ? i_input_data[299 % IN_WIDTH] : pong_storage_data_227 ^ i_input_data[299 % IN_WIDTH];
                397 / IN_WIDTH: pong_storage_data_227 <= (fillup_transition == 1'b1) ? i_input_data[397 % IN_WIDTH] : pong_storage_data_227 ^ i_input_data[397 % IN_WIDTH];
                530 / IN_WIDTH: pong_storage_data_227 <= (fillup_transition == 1'b1) ? i_input_data[530 % IN_WIDTH] : pong_storage_data_227 ^ i_input_data[530 % IN_WIDTH];
                674 / IN_WIDTH: pong_storage_data_227 <= (fillup_transition == 1'b1) ? i_input_data[674 % IN_WIDTH] : pong_storage_data_227 ^ i_input_data[674 % IN_WIDTH];
                1091 / IN_WIDTH: pong_storage_data_227 <= (fillup_transition == 1'b1) ? i_input_data[1091 % IN_WIDTH] : pong_storage_data_227 ^ i_input_data[1091 % IN_WIDTH];
                default: pong_storage_data_227 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_227;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_227 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_227;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_227 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_227;
            end
        end
    end
end

logic ping_storage_data_228;
logic pong_storage_data_228;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_228 <= 1'b0;
        pong_storage_data_228 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                300 / IN_WIDTH: ping_storage_data_228 <= (fillup_transition == 1'b1) ? i_input_data[300 % IN_WIDTH] : ping_storage_data_228 ^ i_input_data[300 % IN_WIDTH];
                398 / IN_WIDTH: ping_storage_data_228 <= (fillup_transition == 1'b1) ? i_input_data[398 % IN_WIDTH] : ping_storage_data_228 ^ i_input_data[398 % IN_WIDTH];
                531 / IN_WIDTH: ping_storage_data_228 <= (fillup_transition == 1'b1) ? i_input_data[531 % IN_WIDTH] : ping_storage_data_228 ^ i_input_data[531 % IN_WIDTH];
                675 / IN_WIDTH: ping_storage_data_228 <= (fillup_transition == 1'b1) ? i_input_data[675 % IN_WIDTH] : ping_storage_data_228 ^ i_input_data[675 % IN_WIDTH];
                1092 / IN_WIDTH: ping_storage_data_228 <= (fillup_transition == 1'b1) ? i_input_data[1092 % IN_WIDTH] : ping_storage_data_228 ^ i_input_data[1092 % IN_WIDTH];
                default: ping_storage_data_228 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_228;
                endcase
            end else begin
                case (input_count)
                300 / IN_WIDTH: pong_storage_data_228 <= (fillup_transition == 1'b1) ? i_input_data[300 % IN_WIDTH] : pong_storage_data_228 ^ i_input_data[300 % IN_WIDTH];
                398 / IN_WIDTH: pong_storage_data_228 <= (fillup_transition == 1'b1) ? i_input_data[398 % IN_WIDTH] : pong_storage_data_228 ^ i_input_data[398 % IN_WIDTH];
                531 / IN_WIDTH: pong_storage_data_228 <= (fillup_transition == 1'b1) ? i_input_data[531 % IN_WIDTH] : pong_storage_data_228 ^ i_input_data[531 % IN_WIDTH];
                675 / IN_WIDTH: pong_storage_data_228 <= (fillup_transition == 1'b1) ? i_input_data[675 % IN_WIDTH] : pong_storage_data_228 ^ i_input_data[675 % IN_WIDTH];
                1092 / IN_WIDTH: pong_storage_data_228 <= (fillup_transition == 1'b1) ? i_input_data[1092 % IN_WIDTH] : pong_storage_data_228 ^ i_input_data[1092 % IN_WIDTH];
                default: pong_storage_data_228 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_228;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_228 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_228;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_228 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_228;
            end
        end
    end
end

logic ping_storage_data_229;
logic pong_storage_data_229;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_229 <= 1'b0;
        pong_storage_data_229 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                301 / IN_WIDTH: ping_storage_data_229 <= (fillup_transition == 1'b1) ? i_input_data[301 % IN_WIDTH] : ping_storage_data_229 ^ i_input_data[301 % IN_WIDTH];
                399 / IN_WIDTH: ping_storage_data_229 <= (fillup_transition == 1'b1) ? i_input_data[399 % IN_WIDTH] : ping_storage_data_229 ^ i_input_data[399 % IN_WIDTH];
                532 / IN_WIDTH: ping_storage_data_229 <= (fillup_transition == 1'b1) ? i_input_data[532 % IN_WIDTH] : ping_storage_data_229 ^ i_input_data[532 % IN_WIDTH];
                676 / IN_WIDTH: ping_storage_data_229 <= (fillup_transition == 1'b1) ? i_input_data[676 % IN_WIDTH] : ping_storage_data_229 ^ i_input_data[676 % IN_WIDTH];
                1093 / IN_WIDTH: ping_storage_data_229 <= (fillup_transition == 1'b1) ? i_input_data[1093 % IN_WIDTH] : ping_storage_data_229 ^ i_input_data[1093 % IN_WIDTH];
                default: ping_storage_data_229 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_229;
                endcase
            end else begin
                case (input_count)
                301 / IN_WIDTH: pong_storage_data_229 <= (fillup_transition == 1'b1) ? i_input_data[301 % IN_WIDTH] : pong_storage_data_229 ^ i_input_data[301 % IN_WIDTH];
                399 / IN_WIDTH: pong_storage_data_229 <= (fillup_transition == 1'b1) ? i_input_data[399 % IN_WIDTH] : pong_storage_data_229 ^ i_input_data[399 % IN_WIDTH];
                532 / IN_WIDTH: pong_storage_data_229 <= (fillup_transition == 1'b1) ? i_input_data[532 % IN_WIDTH] : pong_storage_data_229 ^ i_input_data[532 % IN_WIDTH];
                676 / IN_WIDTH: pong_storage_data_229 <= (fillup_transition == 1'b1) ? i_input_data[676 % IN_WIDTH] : pong_storage_data_229 ^ i_input_data[676 % IN_WIDTH];
                1093 / IN_WIDTH: pong_storage_data_229 <= (fillup_transition == 1'b1) ? i_input_data[1093 % IN_WIDTH] : pong_storage_data_229 ^ i_input_data[1093 % IN_WIDTH];
                default: pong_storage_data_229 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_229;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_229 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_229;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_229 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_229;
            end
        end
    end
end

logic ping_storage_data_230;
logic pong_storage_data_230;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_230 <= 1'b0;
        pong_storage_data_230 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                302 / IN_WIDTH: ping_storage_data_230 <= (fillup_transition == 1'b1) ? i_input_data[302 % IN_WIDTH] : ping_storage_data_230 ^ i_input_data[302 % IN_WIDTH];
                400 / IN_WIDTH: ping_storage_data_230 <= (fillup_transition == 1'b1) ? i_input_data[400 % IN_WIDTH] : ping_storage_data_230 ^ i_input_data[400 % IN_WIDTH];
                533 / IN_WIDTH: ping_storage_data_230 <= (fillup_transition == 1'b1) ? i_input_data[533 % IN_WIDTH] : ping_storage_data_230 ^ i_input_data[533 % IN_WIDTH];
                677 / IN_WIDTH: ping_storage_data_230 <= (fillup_transition == 1'b1) ? i_input_data[677 % IN_WIDTH] : ping_storage_data_230 ^ i_input_data[677 % IN_WIDTH];
                1094 / IN_WIDTH: ping_storage_data_230 <= (fillup_transition == 1'b1) ? i_input_data[1094 % IN_WIDTH] : ping_storage_data_230 ^ i_input_data[1094 % IN_WIDTH];
                default: ping_storage_data_230 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_230;
                endcase
            end else begin
                case (input_count)
                302 / IN_WIDTH: pong_storage_data_230 <= (fillup_transition == 1'b1) ? i_input_data[302 % IN_WIDTH] : pong_storage_data_230 ^ i_input_data[302 % IN_WIDTH];
                400 / IN_WIDTH: pong_storage_data_230 <= (fillup_transition == 1'b1) ? i_input_data[400 % IN_WIDTH] : pong_storage_data_230 ^ i_input_data[400 % IN_WIDTH];
                533 / IN_WIDTH: pong_storage_data_230 <= (fillup_transition == 1'b1) ? i_input_data[533 % IN_WIDTH] : pong_storage_data_230 ^ i_input_data[533 % IN_WIDTH];
                677 / IN_WIDTH: pong_storage_data_230 <= (fillup_transition == 1'b1) ? i_input_data[677 % IN_WIDTH] : pong_storage_data_230 ^ i_input_data[677 % IN_WIDTH];
                1094 / IN_WIDTH: pong_storage_data_230 <= (fillup_transition == 1'b1) ? i_input_data[1094 % IN_WIDTH] : pong_storage_data_230 ^ i_input_data[1094 % IN_WIDTH];
                default: pong_storage_data_230 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_230;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_230 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_230;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_230 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_230;
            end
        end
    end
end

logic ping_storage_data_231;
logic pong_storage_data_231;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_231 <= 1'b0;
        pong_storage_data_231 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                303 / IN_WIDTH: ping_storage_data_231 <= (fillup_transition == 1'b1) ? i_input_data[303 % IN_WIDTH] : ping_storage_data_231 ^ i_input_data[303 % IN_WIDTH];
                401 / IN_WIDTH: ping_storage_data_231 <= (fillup_transition == 1'b1) ? i_input_data[401 % IN_WIDTH] : ping_storage_data_231 ^ i_input_data[401 % IN_WIDTH];
                534 / IN_WIDTH: ping_storage_data_231 <= (fillup_transition == 1'b1) ? i_input_data[534 % IN_WIDTH] : ping_storage_data_231 ^ i_input_data[534 % IN_WIDTH];
                678 / IN_WIDTH: ping_storage_data_231 <= (fillup_transition == 1'b1) ? i_input_data[678 % IN_WIDTH] : ping_storage_data_231 ^ i_input_data[678 % IN_WIDTH];
                1095 / IN_WIDTH: ping_storage_data_231 <= (fillup_transition == 1'b1) ? i_input_data[1095 % IN_WIDTH] : ping_storage_data_231 ^ i_input_data[1095 % IN_WIDTH];
                default: ping_storage_data_231 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_231;
                endcase
            end else begin
                case (input_count)
                303 / IN_WIDTH: pong_storage_data_231 <= (fillup_transition == 1'b1) ? i_input_data[303 % IN_WIDTH] : pong_storage_data_231 ^ i_input_data[303 % IN_WIDTH];
                401 / IN_WIDTH: pong_storage_data_231 <= (fillup_transition == 1'b1) ? i_input_data[401 % IN_WIDTH] : pong_storage_data_231 ^ i_input_data[401 % IN_WIDTH];
                534 / IN_WIDTH: pong_storage_data_231 <= (fillup_transition == 1'b1) ? i_input_data[534 % IN_WIDTH] : pong_storage_data_231 ^ i_input_data[534 % IN_WIDTH];
                678 / IN_WIDTH: pong_storage_data_231 <= (fillup_transition == 1'b1) ? i_input_data[678 % IN_WIDTH] : pong_storage_data_231 ^ i_input_data[678 % IN_WIDTH];
                1095 / IN_WIDTH: pong_storage_data_231 <= (fillup_transition == 1'b1) ? i_input_data[1095 % IN_WIDTH] : pong_storage_data_231 ^ i_input_data[1095 % IN_WIDTH];
                default: pong_storage_data_231 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_231;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_231 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_231;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_231 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_231;
            end
        end
    end
end

logic ping_storage_data_232;
logic pong_storage_data_232;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_232 <= 1'b0;
        pong_storage_data_232 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                304 / IN_WIDTH: ping_storage_data_232 <= (fillup_transition == 1'b1) ? i_input_data[304 % IN_WIDTH] : ping_storage_data_232 ^ i_input_data[304 % IN_WIDTH];
                402 / IN_WIDTH: ping_storage_data_232 <= (fillup_transition == 1'b1) ? i_input_data[402 % IN_WIDTH] : ping_storage_data_232 ^ i_input_data[402 % IN_WIDTH];
                535 / IN_WIDTH: ping_storage_data_232 <= (fillup_transition == 1'b1) ? i_input_data[535 % IN_WIDTH] : ping_storage_data_232 ^ i_input_data[535 % IN_WIDTH];
                679 / IN_WIDTH: ping_storage_data_232 <= (fillup_transition == 1'b1) ? i_input_data[679 % IN_WIDTH] : ping_storage_data_232 ^ i_input_data[679 % IN_WIDTH];
                1096 / IN_WIDTH: ping_storage_data_232 <= (fillup_transition == 1'b1) ? i_input_data[1096 % IN_WIDTH] : ping_storage_data_232 ^ i_input_data[1096 % IN_WIDTH];
                default: ping_storage_data_232 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_232;
                endcase
            end else begin
                case (input_count)
                304 / IN_WIDTH: pong_storage_data_232 <= (fillup_transition == 1'b1) ? i_input_data[304 % IN_WIDTH] : pong_storage_data_232 ^ i_input_data[304 % IN_WIDTH];
                402 / IN_WIDTH: pong_storage_data_232 <= (fillup_transition == 1'b1) ? i_input_data[402 % IN_WIDTH] : pong_storage_data_232 ^ i_input_data[402 % IN_WIDTH];
                535 / IN_WIDTH: pong_storage_data_232 <= (fillup_transition == 1'b1) ? i_input_data[535 % IN_WIDTH] : pong_storage_data_232 ^ i_input_data[535 % IN_WIDTH];
                679 / IN_WIDTH: pong_storage_data_232 <= (fillup_transition == 1'b1) ? i_input_data[679 % IN_WIDTH] : pong_storage_data_232 ^ i_input_data[679 % IN_WIDTH];
                1096 / IN_WIDTH: pong_storage_data_232 <= (fillup_transition == 1'b1) ? i_input_data[1096 % IN_WIDTH] : pong_storage_data_232 ^ i_input_data[1096 % IN_WIDTH];
                default: pong_storage_data_232 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_232;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_232 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_232;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_232 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_232;
            end
        end
    end
end

logic ping_storage_data_233;
logic pong_storage_data_233;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_233 <= 1'b0;
        pong_storage_data_233 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                305 / IN_WIDTH: ping_storage_data_233 <= (fillup_transition == 1'b1) ? i_input_data[305 % IN_WIDTH] : ping_storage_data_233 ^ i_input_data[305 % IN_WIDTH];
                403 / IN_WIDTH: ping_storage_data_233 <= (fillup_transition == 1'b1) ? i_input_data[403 % IN_WIDTH] : ping_storage_data_233 ^ i_input_data[403 % IN_WIDTH];
                536 / IN_WIDTH: ping_storage_data_233 <= (fillup_transition == 1'b1) ? i_input_data[536 % IN_WIDTH] : ping_storage_data_233 ^ i_input_data[536 % IN_WIDTH];
                680 / IN_WIDTH: ping_storage_data_233 <= (fillup_transition == 1'b1) ? i_input_data[680 % IN_WIDTH] : ping_storage_data_233 ^ i_input_data[680 % IN_WIDTH];
                1097 / IN_WIDTH: ping_storage_data_233 <= (fillup_transition == 1'b1) ? i_input_data[1097 % IN_WIDTH] : ping_storage_data_233 ^ i_input_data[1097 % IN_WIDTH];
                default: ping_storage_data_233 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_233;
                endcase
            end else begin
                case (input_count)
                305 / IN_WIDTH: pong_storage_data_233 <= (fillup_transition == 1'b1) ? i_input_data[305 % IN_WIDTH] : pong_storage_data_233 ^ i_input_data[305 % IN_WIDTH];
                403 / IN_WIDTH: pong_storage_data_233 <= (fillup_transition == 1'b1) ? i_input_data[403 % IN_WIDTH] : pong_storage_data_233 ^ i_input_data[403 % IN_WIDTH];
                536 / IN_WIDTH: pong_storage_data_233 <= (fillup_transition == 1'b1) ? i_input_data[536 % IN_WIDTH] : pong_storage_data_233 ^ i_input_data[536 % IN_WIDTH];
                680 / IN_WIDTH: pong_storage_data_233 <= (fillup_transition == 1'b1) ? i_input_data[680 % IN_WIDTH] : pong_storage_data_233 ^ i_input_data[680 % IN_WIDTH];
                1097 / IN_WIDTH: pong_storage_data_233 <= (fillup_transition == 1'b1) ? i_input_data[1097 % IN_WIDTH] : pong_storage_data_233 ^ i_input_data[1097 % IN_WIDTH];
                default: pong_storage_data_233 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_233;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_233 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_233;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_233 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_233;
            end
        end
    end
end

logic ping_storage_data_234;
logic pong_storage_data_234;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_234 <= 1'b0;
        pong_storage_data_234 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                306 / IN_WIDTH: ping_storage_data_234 <= (fillup_transition == 1'b1) ? i_input_data[306 % IN_WIDTH] : ping_storage_data_234 ^ i_input_data[306 % IN_WIDTH];
                404 / IN_WIDTH: ping_storage_data_234 <= (fillup_transition == 1'b1) ? i_input_data[404 % IN_WIDTH] : ping_storage_data_234 ^ i_input_data[404 % IN_WIDTH];
                537 / IN_WIDTH: ping_storage_data_234 <= (fillup_transition == 1'b1) ? i_input_data[537 % IN_WIDTH] : ping_storage_data_234 ^ i_input_data[537 % IN_WIDTH];
                681 / IN_WIDTH: ping_storage_data_234 <= (fillup_transition == 1'b1) ? i_input_data[681 % IN_WIDTH] : ping_storage_data_234 ^ i_input_data[681 % IN_WIDTH];
                1098 / IN_WIDTH: ping_storage_data_234 <= (fillup_transition == 1'b1) ? i_input_data[1098 % IN_WIDTH] : ping_storage_data_234 ^ i_input_data[1098 % IN_WIDTH];
                default: ping_storage_data_234 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_234;
                endcase
            end else begin
                case (input_count)
                306 / IN_WIDTH: pong_storage_data_234 <= (fillup_transition == 1'b1) ? i_input_data[306 % IN_WIDTH] : pong_storage_data_234 ^ i_input_data[306 % IN_WIDTH];
                404 / IN_WIDTH: pong_storage_data_234 <= (fillup_transition == 1'b1) ? i_input_data[404 % IN_WIDTH] : pong_storage_data_234 ^ i_input_data[404 % IN_WIDTH];
                537 / IN_WIDTH: pong_storage_data_234 <= (fillup_transition == 1'b1) ? i_input_data[537 % IN_WIDTH] : pong_storage_data_234 ^ i_input_data[537 % IN_WIDTH];
                681 / IN_WIDTH: pong_storage_data_234 <= (fillup_transition == 1'b1) ? i_input_data[681 % IN_WIDTH] : pong_storage_data_234 ^ i_input_data[681 % IN_WIDTH];
                1098 / IN_WIDTH: pong_storage_data_234 <= (fillup_transition == 1'b1) ? i_input_data[1098 % IN_WIDTH] : pong_storage_data_234 ^ i_input_data[1098 % IN_WIDTH];
                default: pong_storage_data_234 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_234;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_234 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_234;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_234 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_234;
            end
        end
    end
end

logic ping_storage_data_235;
logic pong_storage_data_235;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_235 <= 1'b0;
        pong_storage_data_235 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                307 / IN_WIDTH: ping_storage_data_235 <= (fillup_transition == 1'b1) ? i_input_data[307 % IN_WIDTH] : ping_storage_data_235 ^ i_input_data[307 % IN_WIDTH];
                405 / IN_WIDTH: ping_storage_data_235 <= (fillup_transition == 1'b1) ? i_input_data[405 % IN_WIDTH] : ping_storage_data_235 ^ i_input_data[405 % IN_WIDTH];
                538 / IN_WIDTH: ping_storage_data_235 <= (fillup_transition == 1'b1) ? i_input_data[538 % IN_WIDTH] : ping_storage_data_235 ^ i_input_data[538 % IN_WIDTH];
                682 / IN_WIDTH: ping_storage_data_235 <= (fillup_transition == 1'b1) ? i_input_data[682 % IN_WIDTH] : ping_storage_data_235 ^ i_input_data[682 % IN_WIDTH];
                1099 / IN_WIDTH: ping_storage_data_235 <= (fillup_transition == 1'b1) ? i_input_data[1099 % IN_WIDTH] : ping_storage_data_235 ^ i_input_data[1099 % IN_WIDTH];
                default: ping_storage_data_235 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_235;
                endcase
            end else begin
                case (input_count)
                307 / IN_WIDTH: pong_storage_data_235 <= (fillup_transition == 1'b1) ? i_input_data[307 % IN_WIDTH] : pong_storage_data_235 ^ i_input_data[307 % IN_WIDTH];
                405 / IN_WIDTH: pong_storage_data_235 <= (fillup_transition == 1'b1) ? i_input_data[405 % IN_WIDTH] : pong_storage_data_235 ^ i_input_data[405 % IN_WIDTH];
                538 / IN_WIDTH: pong_storage_data_235 <= (fillup_transition == 1'b1) ? i_input_data[538 % IN_WIDTH] : pong_storage_data_235 ^ i_input_data[538 % IN_WIDTH];
                682 / IN_WIDTH: pong_storage_data_235 <= (fillup_transition == 1'b1) ? i_input_data[682 % IN_WIDTH] : pong_storage_data_235 ^ i_input_data[682 % IN_WIDTH];
                1099 / IN_WIDTH: pong_storage_data_235 <= (fillup_transition == 1'b1) ? i_input_data[1099 % IN_WIDTH] : pong_storage_data_235 ^ i_input_data[1099 % IN_WIDTH];
                default: pong_storage_data_235 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_235;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_235 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_235;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_235 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_235;
            end
        end
    end
end

logic ping_storage_data_236;
logic pong_storage_data_236;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_236 <= 1'b0;
        pong_storage_data_236 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                308 / IN_WIDTH: ping_storage_data_236 <= (fillup_transition == 1'b1) ? i_input_data[308 % IN_WIDTH] : ping_storage_data_236 ^ i_input_data[308 % IN_WIDTH];
                406 / IN_WIDTH: ping_storage_data_236 <= (fillup_transition == 1'b1) ? i_input_data[406 % IN_WIDTH] : ping_storage_data_236 ^ i_input_data[406 % IN_WIDTH];
                539 / IN_WIDTH: ping_storage_data_236 <= (fillup_transition == 1'b1) ? i_input_data[539 % IN_WIDTH] : ping_storage_data_236 ^ i_input_data[539 % IN_WIDTH];
                683 / IN_WIDTH: ping_storage_data_236 <= (fillup_transition == 1'b1) ? i_input_data[683 % IN_WIDTH] : ping_storage_data_236 ^ i_input_data[683 % IN_WIDTH];
                1100 / IN_WIDTH: ping_storage_data_236 <= (fillup_transition == 1'b1) ? i_input_data[1100 % IN_WIDTH] : ping_storage_data_236 ^ i_input_data[1100 % IN_WIDTH];
                default: ping_storage_data_236 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_236;
                endcase
            end else begin
                case (input_count)
                308 / IN_WIDTH: pong_storage_data_236 <= (fillup_transition == 1'b1) ? i_input_data[308 % IN_WIDTH] : pong_storage_data_236 ^ i_input_data[308 % IN_WIDTH];
                406 / IN_WIDTH: pong_storage_data_236 <= (fillup_transition == 1'b1) ? i_input_data[406 % IN_WIDTH] : pong_storage_data_236 ^ i_input_data[406 % IN_WIDTH];
                539 / IN_WIDTH: pong_storage_data_236 <= (fillup_transition == 1'b1) ? i_input_data[539 % IN_WIDTH] : pong_storage_data_236 ^ i_input_data[539 % IN_WIDTH];
                683 / IN_WIDTH: pong_storage_data_236 <= (fillup_transition == 1'b1) ? i_input_data[683 % IN_WIDTH] : pong_storage_data_236 ^ i_input_data[683 % IN_WIDTH];
                1100 / IN_WIDTH: pong_storage_data_236 <= (fillup_transition == 1'b1) ? i_input_data[1100 % IN_WIDTH] : pong_storage_data_236 ^ i_input_data[1100 % IN_WIDTH];
                default: pong_storage_data_236 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_236;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_236 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_236;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_236 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_236;
            end
        end
    end
end

logic ping_storage_data_237;
logic pong_storage_data_237;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_237 <= 1'b0;
        pong_storage_data_237 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                309 / IN_WIDTH: ping_storage_data_237 <= (fillup_transition == 1'b1) ? i_input_data[309 % IN_WIDTH] : ping_storage_data_237 ^ i_input_data[309 % IN_WIDTH];
                407 / IN_WIDTH: ping_storage_data_237 <= (fillup_transition == 1'b1) ? i_input_data[407 % IN_WIDTH] : ping_storage_data_237 ^ i_input_data[407 % IN_WIDTH];
                540 / IN_WIDTH: ping_storage_data_237 <= (fillup_transition == 1'b1) ? i_input_data[540 % IN_WIDTH] : ping_storage_data_237 ^ i_input_data[540 % IN_WIDTH];
                684 / IN_WIDTH: ping_storage_data_237 <= (fillup_transition == 1'b1) ? i_input_data[684 % IN_WIDTH] : ping_storage_data_237 ^ i_input_data[684 % IN_WIDTH];
                1101 / IN_WIDTH: ping_storage_data_237 <= (fillup_transition == 1'b1) ? i_input_data[1101 % IN_WIDTH] : ping_storage_data_237 ^ i_input_data[1101 % IN_WIDTH];
                default: ping_storage_data_237 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_237;
                endcase
            end else begin
                case (input_count)
                309 / IN_WIDTH: pong_storage_data_237 <= (fillup_transition == 1'b1) ? i_input_data[309 % IN_WIDTH] : pong_storage_data_237 ^ i_input_data[309 % IN_WIDTH];
                407 / IN_WIDTH: pong_storage_data_237 <= (fillup_transition == 1'b1) ? i_input_data[407 % IN_WIDTH] : pong_storage_data_237 ^ i_input_data[407 % IN_WIDTH];
                540 / IN_WIDTH: pong_storage_data_237 <= (fillup_transition == 1'b1) ? i_input_data[540 % IN_WIDTH] : pong_storage_data_237 ^ i_input_data[540 % IN_WIDTH];
                684 / IN_WIDTH: pong_storage_data_237 <= (fillup_transition == 1'b1) ? i_input_data[684 % IN_WIDTH] : pong_storage_data_237 ^ i_input_data[684 % IN_WIDTH];
                1101 / IN_WIDTH: pong_storage_data_237 <= (fillup_transition == 1'b1) ? i_input_data[1101 % IN_WIDTH] : pong_storage_data_237 ^ i_input_data[1101 % IN_WIDTH];
                default: pong_storage_data_237 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_237;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_237 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_237;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_237 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_237;
            end
        end
    end
end

logic ping_storage_data_238;
logic pong_storage_data_238;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_238 <= 1'b0;
        pong_storage_data_238 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                310 / IN_WIDTH: ping_storage_data_238 <= (fillup_transition == 1'b1) ? i_input_data[310 % IN_WIDTH] : ping_storage_data_238 ^ i_input_data[310 % IN_WIDTH];
                408 / IN_WIDTH: ping_storage_data_238 <= (fillup_transition == 1'b1) ? i_input_data[408 % IN_WIDTH] : ping_storage_data_238 ^ i_input_data[408 % IN_WIDTH];
                541 / IN_WIDTH: ping_storage_data_238 <= (fillup_transition == 1'b1) ? i_input_data[541 % IN_WIDTH] : ping_storage_data_238 ^ i_input_data[541 % IN_WIDTH];
                685 / IN_WIDTH: ping_storage_data_238 <= (fillup_transition == 1'b1) ? i_input_data[685 % IN_WIDTH] : ping_storage_data_238 ^ i_input_data[685 % IN_WIDTH];
                1102 / IN_WIDTH: ping_storage_data_238 <= (fillup_transition == 1'b1) ? i_input_data[1102 % IN_WIDTH] : ping_storage_data_238 ^ i_input_data[1102 % IN_WIDTH];
                default: ping_storage_data_238 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_238;
                endcase
            end else begin
                case (input_count)
                310 / IN_WIDTH: pong_storage_data_238 <= (fillup_transition == 1'b1) ? i_input_data[310 % IN_WIDTH] : pong_storage_data_238 ^ i_input_data[310 % IN_WIDTH];
                408 / IN_WIDTH: pong_storage_data_238 <= (fillup_transition == 1'b1) ? i_input_data[408 % IN_WIDTH] : pong_storage_data_238 ^ i_input_data[408 % IN_WIDTH];
                541 / IN_WIDTH: pong_storage_data_238 <= (fillup_transition == 1'b1) ? i_input_data[541 % IN_WIDTH] : pong_storage_data_238 ^ i_input_data[541 % IN_WIDTH];
                685 / IN_WIDTH: pong_storage_data_238 <= (fillup_transition == 1'b1) ? i_input_data[685 % IN_WIDTH] : pong_storage_data_238 ^ i_input_data[685 % IN_WIDTH];
                1102 / IN_WIDTH: pong_storage_data_238 <= (fillup_transition == 1'b1) ? i_input_data[1102 % IN_WIDTH] : pong_storage_data_238 ^ i_input_data[1102 % IN_WIDTH];
                default: pong_storage_data_238 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_238;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_238 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_238;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_238 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_238;
            end
        end
    end
end

logic ping_storage_data_239;
logic pong_storage_data_239;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_239 <= 1'b0;
        pong_storage_data_239 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                311 / IN_WIDTH: ping_storage_data_239 <= (fillup_transition == 1'b1) ? i_input_data[311 % IN_WIDTH] : ping_storage_data_239 ^ i_input_data[311 % IN_WIDTH];
                409 / IN_WIDTH: ping_storage_data_239 <= (fillup_transition == 1'b1) ? i_input_data[409 % IN_WIDTH] : ping_storage_data_239 ^ i_input_data[409 % IN_WIDTH];
                542 / IN_WIDTH: ping_storage_data_239 <= (fillup_transition == 1'b1) ? i_input_data[542 % IN_WIDTH] : ping_storage_data_239 ^ i_input_data[542 % IN_WIDTH];
                686 / IN_WIDTH: ping_storage_data_239 <= (fillup_transition == 1'b1) ? i_input_data[686 % IN_WIDTH] : ping_storage_data_239 ^ i_input_data[686 % IN_WIDTH];
                1103 / IN_WIDTH: ping_storage_data_239 <= (fillup_transition == 1'b1) ? i_input_data[1103 % IN_WIDTH] : ping_storage_data_239 ^ i_input_data[1103 % IN_WIDTH];
                default: ping_storage_data_239 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_239;
                endcase
            end else begin
                case (input_count)
                311 / IN_WIDTH: pong_storage_data_239 <= (fillup_transition == 1'b1) ? i_input_data[311 % IN_WIDTH] : pong_storage_data_239 ^ i_input_data[311 % IN_WIDTH];
                409 / IN_WIDTH: pong_storage_data_239 <= (fillup_transition == 1'b1) ? i_input_data[409 % IN_WIDTH] : pong_storage_data_239 ^ i_input_data[409 % IN_WIDTH];
                542 / IN_WIDTH: pong_storage_data_239 <= (fillup_transition == 1'b1) ? i_input_data[542 % IN_WIDTH] : pong_storage_data_239 ^ i_input_data[542 % IN_WIDTH];
                686 / IN_WIDTH: pong_storage_data_239 <= (fillup_transition == 1'b1) ? i_input_data[686 % IN_WIDTH] : pong_storage_data_239 ^ i_input_data[686 % IN_WIDTH];
                1103 / IN_WIDTH: pong_storage_data_239 <= (fillup_transition == 1'b1) ? i_input_data[1103 % IN_WIDTH] : pong_storage_data_239 ^ i_input_data[1103 % IN_WIDTH];
                default: pong_storage_data_239 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_239;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_239 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_239;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_239 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_239;
            end
        end
    end
end

logic ping_storage_data_240;
logic pong_storage_data_240;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_240 <= 1'b0;
        pong_storage_data_240 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                312 / IN_WIDTH: ping_storage_data_240 <= (fillup_transition == 1'b1) ? i_input_data[312 % IN_WIDTH] : ping_storage_data_240 ^ i_input_data[312 % IN_WIDTH];
                410 / IN_WIDTH: ping_storage_data_240 <= (fillup_transition == 1'b1) ? i_input_data[410 % IN_WIDTH] : ping_storage_data_240 ^ i_input_data[410 % IN_WIDTH];
                543 / IN_WIDTH: ping_storage_data_240 <= (fillup_transition == 1'b1) ? i_input_data[543 % IN_WIDTH] : ping_storage_data_240 ^ i_input_data[543 % IN_WIDTH];
                687 / IN_WIDTH: ping_storage_data_240 <= (fillup_transition == 1'b1) ? i_input_data[687 % IN_WIDTH] : ping_storage_data_240 ^ i_input_data[687 % IN_WIDTH];
                1104 / IN_WIDTH: ping_storage_data_240 <= (fillup_transition == 1'b1) ? i_input_data[1104 % IN_WIDTH] : ping_storage_data_240 ^ i_input_data[1104 % IN_WIDTH];
                default: ping_storage_data_240 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_240;
                endcase
            end else begin
                case (input_count)
                312 / IN_WIDTH: pong_storage_data_240 <= (fillup_transition == 1'b1) ? i_input_data[312 % IN_WIDTH] : pong_storage_data_240 ^ i_input_data[312 % IN_WIDTH];
                410 / IN_WIDTH: pong_storage_data_240 <= (fillup_transition == 1'b1) ? i_input_data[410 % IN_WIDTH] : pong_storage_data_240 ^ i_input_data[410 % IN_WIDTH];
                543 / IN_WIDTH: pong_storage_data_240 <= (fillup_transition == 1'b1) ? i_input_data[543 % IN_WIDTH] : pong_storage_data_240 ^ i_input_data[543 % IN_WIDTH];
                687 / IN_WIDTH: pong_storage_data_240 <= (fillup_transition == 1'b1) ? i_input_data[687 % IN_WIDTH] : pong_storage_data_240 ^ i_input_data[687 % IN_WIDTH];
                1104 / IN_WIDTH: pong_storage_data_240 <= (fillup_transition == 1'b1) ? i_input_data[1104 % IN_WIDTH] : pong_storage_data_240 ^ i_input_data[1104 % IN_WIDTH];
                default: pong_storage_data_240 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_240;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_240 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_240;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_240 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_240;
            end
        end
    end
end

logic ping_storage_data_241;
logic pong_storage_data_241;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_241 <= 1'b0;
        pong_storage_data_241 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                313 / IN_WIDTH: ping_storage_data_241 <= (fillup_transition == 1'b1) ? i_input_data[313 % IN_WIDTH] : ping_storage_data_241 ^ i_input_data[313 % IN_WIDTH];
                411 / IN_WIDTH: ping_storage_data_241 <= (fillup_transition == 1'b1) ? i_input_data[411 % IN_WIDTH] : ping_storage_data_241 ^ i_input_data[411 % IN_WIDTH];
                544 / IN_WIDTH: ping_storage_data_241 <= (fillup_transition == 1'b1) ? i_input_data[544 % IN_WIDTH] : ping_storage_data_241 ^ i_input_data[544 % IN_WIDTH];
                688 / IN_WIDTH: ping_storage_data_241 <= (fillup_transition == 1'b1) ? i_input_data[688 % IN_WIDTH] : ping_storage_data_241 ^ i_input_data[688 % IN_WIDTH];
                1105 / IN_WIDTH: ping_storage_data_241 <= (fillup_transition == 1'b1) ? i_input_data[1105 % IN_WIDTH] : ping_storage_data_241 ^ i_input_data[1105 % IN_WIDTH];
                default: ping_storage_data_241 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_241;
                endcase
            end else begin
                case (input_count)
                313 / IN_WIDTH: pong_storage_data_241 <= (fillup_transition == 1'b1) ? i_input_data[313 % IN_WIDTH] : pong_storage_data_241 ^ i_input_data[313 % IN_WIDTH];
                411 / IN_WIDTH: pong_storage_data_241 <= (fillup_transition == 1'b1) ? i_input_data[411 % IN_WIDTH] : pong_storage_data_241 ^ i_input_data[411 % IN_WIDTH];
                544 / IN_WIDTH: pong_storage_data_241 <= (fillup_transition == 1'b1) ? i_input_data[544 % IN_WIDTH] : pong_storage_data_241 ^ i_input_data[544 % IN_WIDTH];
                688 / IN_WIDTH: pong_storage_data_241 <= (fillup_transition == 1'b1) ? i_input_data[688 % IN_WIDTH] : pong_storage_data_241 ^ i_input_data[688 % IN_WIDTH];
                1105 / IN_WIDTH: pong_storage_data_241 <= (fillup_transition == 1'b1) ? i_input_data[1105 % IN_WIDTH] : pong_storage_data_241 ^ i_input_data[1105 % IN_WIDTH];
                default: pong_storage_data_241 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_241;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_241 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_241;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_241 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_241;
            end
        end
    end
end

logic ping_storage_data_242;
logic pong_storage_data_242;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_242 <= 1'b0;
        pong_storage_data_242 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                314 / IN_WIDTH: ping_storage_data_242 <= (fillup_transition == 1'b1) ? i_input_data[314 % IN_WIDTH] : ping_storage_data_242 ^ i_input_data[314 % IN_WIDTH];
                412 / IN_WIDTH: ping_storage_data_242 <= (fillup_transition == 1'b1) ? i_input_data[412 % IN_WIDTH] : ping_storage_data_242 ^ i_input_data[412 % IN_WIDTH];
                545 / IN_WIDTH: ping_storage_data_242 <= (fillup_transition == 1'b1) ? i_input_data[545 % IN_WIDTH] : ping_storage_data_242 ^ i_input_data[545 % IN_WIDTH];
                689 / IN_WIDTH: ping_storage_data_242 <= (fillup_transition == 1'b1) ? i_input_data[689 % IN_WIDTH] : ping_storage_data_242 ^ i_input_data[689 % IN_WIDTH];
                1106 / IN_WIDTH: ping_storage_data_242 <= (fillup_transition == 1'b1) ? i_input_data[1106 % IN_WIDTH] : ping_storage_data_242 ^ i_input_data[1106 % IN_WIDTH];
                default: ping_storage_data_242 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_242;
                endcase
            end else begin
                case (input_count)
                314 / IN_WIDTH: pong_storage_data_242 <= (fillup_transition == 1'b1) ? i_input_data[314 % IN_WIDTH] : pong_storage_data_242 ^ i_input_data[314 % IN_WIDTH];
                412 / IN_WIDTH: pong_storage_data_242 <= (fillup_transition == 1'b1) ? i_input_data[412 % IN_WIDTH] : pong_storage_data_242 ^ i_input_data[412 % IN_WIDTH];
                545 / IN_WIDTH: pong_storage_data_242 <= (fillup_transition == 1'b1) ? i_input_data[545 % IN_WIDTH] : pong_storage_data_242 ^ i_input_data[545 % IN_WIDTH];
                689 / IN_WIDTH: pong_storage_data_242 <= (fillup_transition == 1'b1) ? i_input_data[689 % IN_WIDTH] : pong_storage_data_242 ^ i_input_data[689 % IN_WIDTH];
                1106 / IN_WIDTH: pong_storage_data_242 <= (fillup_transition == 1'b1) ? i_input_data[1106 % IN_WIDTH] : pong_storage_data_242 ^ i_input_data[1106 % IN_WIDTH];
                default: pong_storage_data_242 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_242;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_242 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_242;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_242 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_242;
            end
        end
    end
end

logic ping_storage_data_243;
logic pong_storage_data_243;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_243 <= 1'b0;
        pong_storage_data_243 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                315 / IN_WIDTH: ping_storage_data_243 <= (fillup_transition == 1'b1) ? i_input_data[315 % IN_WIDTH] : ping_storage_data_243 ^ i_input_data[315 % IN_WIDTH];
                413 / IN_WIDTH: ping_storage_data_243 <= (fillup_transition == 1'b1) ? i_input_data[413 % IN_WIDTH] : ping_storage_data_243 ^ i_input_data[413 % IN_WIDTH];
                546 / IN_WIDTH: ping_storage_data_243 <= (fillup_transition == 1'b1) ? i_input_data[546 % IN_WIDTH] : ping_storage_data_243 ^ i_input_data[546 % IN_WIDTH];
                690 / IN_WIDTH: ping_storage_data_243 <= (fillup_transition == 1'b1) ? i_input_data[690 % IN_WIDTH] : ping_storage_data_243 ^ i_input_data[690 % IN_WIDTH];
                1107 / IN_WIDTH: ping_storage_data_243 <= (fillup_transition == 1'b1) ? i_input_data[1107 % IN_WIDTH] : ping_storage_data_243 ^ i_input_data[1107 % IN_WIDTH];
                default: ping_storage_data_243 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_243;
                endcase
            end else begin
                case (input_count)
                315 / IN_WIDTH: pong_storage_data_243 <= (fillup_transition == 1'b1) ? i_input_data[315 % IN_WIDTH] : pong_storage_data_243 ^ i_input_data[315 % IN_WIDTH];
                413 / IN_WIDTH: pong_storage_data_243 <= (fillup_transition == 1'b1) ? i_input_data[413 % IN_WIDTH] : pong_storage_data_243 ^ i_input_data[413 % IN_WIDTH];
                546 / IN_WIDTH: pong_storage_data_243 <= (fillup_transition == 1'b1) ? i_input_data[546 % IN_WIDTH] : pong_storage_data_243 ^ i_input_data[546 % IN_WIDTH];
                690 / IN_WIDTH: pong_storage_data_243 <= (fillup_transition == 1'b1) ? i_input_data[690 % IN_WIDTH] : pong_storage_data_243 ^ i_input_data[690 % IN_WIDTH];
                1107 / IN_WIDTH: pong_storage_data_243 <= (fillup_transition == 1'b1) ? i_input_data[1107 % IN_WIDTH] : pong_storage_data_243 ^ i_input_data[1107 % IN_WIDTH];
                default: pong_storage_data_243 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_243;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_243 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_243;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_243 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_243;
            end
        end
    end
end

logic ping_storage_data_244;
logic pong_storage_data_244;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_244 <= 1'b0;
        pong_storage_data_244 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                316 / IN_WIDTH: ping_storage_data_244 <= (fillup_transition == 1'b1) ? i_input_data[316 % IN_WIDTH] : ping_storage_data_244 ^ i_input_data[316 % IN_WIDTH];
                414 / IN_WIDTH: ping_storage_data_244 <= (fillup_transition == 1'b1) ? i_input_data[414 % IN_WIDTH] : ping_storage_data_244 ^ i_input_data[414 % IN_WIDTH];
                547 / IN_WIDTH: ping_storage_data_244 <= (fillup_transition == 1'b1) ? i_input_data[547 % IN_WIDTH] : ping_storage_data_244 ^ i_input_data[547 % IN_WIDTH];
                691 / IN_WIDTH: ping_storage_data_244 <= (fillup_transition == 1'b1) ? i_input_data[691 % IN_WIDTH] : ping_storage_data_244 ^ i_input_data[691 % IN_WIDTH];
                1108 / IN_WIDTH: ping_storage_data_244 <= (fillup_transition == 1'b1) ? i_input_data[1108 % IN_WIDTH] : ping_storage_data_244 ^ i_input_data[1108 % IN_WIDTH];
                default: ping_storage_data_244 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_244;
                endcase
            end else begin
                case (input_count)
                316 / IN_WIDTH: pong_storage_data_244 <= (fillup_transition == 1'b1) ? i_input_data[316 % IN_WIDTH] : pong_storage_data_244 ^ i_input_data[316 % IN_WIDTH];
                414 / IN_WIDTH: pong_storage_data_244 <= (fillup_transition == 1'b1) ? i_input_data[414 % IN_WIDTH] : pong_storage_data_244 ^ i_input_data[414 % IN_WIDTH];
                547 / IN_WIDTH: pong_storage_data_244 <= (fillup_transition == 1'b1) ? i_input_data[547 % IN_WIDTH] : pong_storage_data_244 ^ i_input_data[547 % IN_WIDTH];
                691 / IN_WIDTH: pong_storage_data_244 <= (fillup_transition == 1'b1) ? i_input_data[691 % IN_WIDTH] : pong_storage_data_244 ^ i_input_data[691 % IN_WIDTH];
                1108 / IN_WIDTH: pong_storage_data_244 <= (fillup_transition == 1'b1) ? i_input_data[1108 % IN_WIDTH] : pong_storage_data_244 ^ i_input_data[1108 % IN_WIDTH];
                default: pong_storage_data_244 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_244;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_244 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_244;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_244 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_244;
            end
        end
    end
end

logic ping_storage_data_245;
logic pong_storage_data_245;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_245 <= 1'b0;
        pong_storage_data_245 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                317 / IN_WIDTH: ping_storage_data_245 <= (fillup_transition == 1'b1) ? i_input_data[317 % IN_WIDTH] : ping_storage_data_245 ^ i_input_data[317 % IN_WIDTH];
                415 / IN_WIDTH: ping_storage_data_245 <= (fillup_transition == 1'b1) ? i_input_data[415 % IN_WIDTH] : ping_storage_data_245 ^ i_input_data[415 % IN_WIDTH];
                548 / IN_WIDTH: ping_storage_data_245 <= (fillup_transition == 1'b1) ? i_input_data[548 % IN_WIDTH] : ping_storage_data_245 ^ i_input_data[548 % IN_WIDTH];
                692 / IN_WIDTH: ping_storage_data_245 <= (fillup_transition == 1'b1) ? i_input_data[692 % IN_WIDTH] : ping_storage_data_245 ^ i_input_data[692 % IN_WIDTH];
                1109 / IN_WIDTH: ping_storage_data_245 <= (fillup_transition == 1'b1) ? i_input_data[1109 % IN_WIDTH] : ping_storage_data_245 ^ i_input_data[1109 % IN_WIDTH];
                default: ping_storage_data_245 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_245;
                endcase
            end else begin
                case (input_count)
                317 / IN_WIDTH: pong_storage_data_245 <= (fillup_transition == 1'b1) ? i_input_data[317 % IN_WIDTH] : pong_storage_data_245 ^ i_input_data[317 % IN_WIDTH];
                415 / IN_WIDTH: pong_storage_data_245 <= (fillup_transition == 1'b1) ? i_input_data[415 % IN_WIDTH] : pong_storage_data_245 ^ i_input_data[415 % IN_WIDTH];
                548 / IN_WIDTH: pong_storage_data_245 <= (fillup_transition == 1'b1) ? i_input_data[548 % IN_WIDTH] : pong_storage_data_245 ^ i_input_data[548 % IN_WIDTH];
                692 / IN_WIDTH: pong_storage_data_245 <= (fillup_transition == 1'b1) ? i_input_data[692 % IN_WIDTH] : pong_storage_data_245 ^ i_input_data[692 % IN_WIDTH];
                1109 / IN_WIDTH: pong_storage_data_245 <= (fillup_transition == 1'b1) ? i_input_data[1109 % IN_WIDTH] : pong_storage_data_245 ^ i_input_data[1109 % IN_WIDTH];
                default: pong_storage_data_245 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_245;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_245 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_245;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_245 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_245;
            end
        end
    end
end

logic ping_storage_data_246;
logic pong_storage_data_246;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_246 <= 1'b0;
        pong_storage_data_246 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                318 / IN_WIDTH: ping_storage_data_246 <= (fillup_transition == 1'b1) ? i_input_data[318 % IN_WIDTH] : ping_storage_data_246 ^ i_input_data[318 % IN_WIDTH];
                416 / IN_WIDTH: ping_storage_data_246 <= (fillup_transition == 1'b1) ? i_input_data[416 % IN_WIDTH] : ping_storage_data_246 ^ i_input_data[416 % IN_WIDTH];
                549 / IN_WIDTH: ping_storage_data_246 <= (fillup_transition == 1'b1) ? i_input_data[549 % IN_WIDTH] : ping_storage_data_246 ^ i_input_data[549 % IN_WIDTH];
                693 / IN_WIDTH: ping_storage_data_246 <= (fillup_transition == 1'b1) ? i_input_data[693 % IN_WIDTH] : ping_storage_data_246 ^ i_input_data[693 % IN_WIDTH];
                1110 / IN_WIDTH: ping_storage_data_246 <= (fillup_transition == 1'b1) ? i_input_data[1110 % IN_WIDTH] : ping_storage_data_246 ^ i_input_data[1110 % IN_WIDTH];
                default: ping_storage_data_246 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_246;
                endcase
            end else begin
                case (input_count)
                318 / IN_WIDTH: pong_storage_data_246 <= (fillup_transition == 1'b1) ? i_input_data[318 % IN_WIDTH] : pong_storage_data_246 ^ i_input_data[318 % IN_WIDTH];
                416 / IN_WIDTH: pong_storage_data_246 <= (fillup_transition == 1'b1) ? i_input_data[416 % IN_WIDTH] : pong_storage_data_246 ^ i_input_data[416 % IN_WIDTH];
                549 / IN_WIDTH: pong_storage_data_246 <= (fillup_transition == 1'b1) ? i_input_data[549 % IN_WIDTH] : pong_storage_data_246 ^ i_input_data[549 % IN_WIDTH];
                693 / IN_WIDTH: pong_storage_data_246 <= (fillup_transition == 1'b1) ? i_input_data[693 % IN_WIDTH] : pong_storage_data_246 ^ i_input_data[693 % IN_WIDTH];
                1110 / IN_WIDTH: pong_storage_data_246 <= (fillup_transition == 1'b1) ? i_input_data[1110 % IN_WIDTH] : pong_storage_data_246 ^ i_input_data[1110 % IN_WIDTH];
                default: pong_storage_data_246 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_246;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_246 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_246;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_246 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_246;
            end
        end
    end
end

logic ping_storage_data_247;
logic pong_storage_data_247;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_247 <= 1'b0;
        pong_storage_data_247 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                319 / IN_WIDTH: ping_storage_data_247 <= (fillup_transition == 1'b1) ? i_input_data[319 % IN_WIDTH] : ping_storage_data_247 ^ i_input_data[319 % IN_WIDTH];
                417 / IN_WIDTH: ping_storage_data_247 <= (fillup_transition == 1'b1) ? i_input_data[417 % IN_WIDTH] : ping_storage_data_247 ^ i_input_data[417 % IN_WIDTH];
                550 / IN_WIDTH: ping_storage_data_247 <= (fillup_transition == 1'b1) ? i_input_data[550 % IN_WIDTH] : ping_storage_data_247 ^ i_input_data[550 % IN_WIDTH];
                694 / IN_WIDTH: ping_storage_data_247 <= (fillup_transition == 1'b1) ? i_input_data[694 % IN_WIDTH] : ping_storage_data_247 ^ i_input_data[694 % IN_WIDTH];
                1111 / IN_WIDTH: ping_storage_data_247 <= (fillup_transition == 1'b1) ? i_input_data[1111 % IN_WIDTH] : ping_storage_data_247 ^ i_input_data[1111 % IN_WIDTH];
                default: ping_storage_data_247 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_247;
                endcase
            end else begin
                case (input_count)
                319 / IN_WIDTH: pong_storage_data_247 <= (fillup_transition == 1'b1) ? i_input_data[319 % IN_WIDTH] : pong_storage_data_247 ^ i_input_data[319 % IN_WIDTH];
                417 / IN_WIDTH: pong_storage_data_247 <= (fillup_transition == 1'b1) ? i_input_data[417 % IN_WIDTH] : pong_storage_data_247 ^ i_input_data[417 % IN_WIDTH];
                550 / IN_WIDTH: pong_storage_data_247 <= (fillup_transition == 1'b1) ? i_input_data[550 % IN_WIDTH] : pong_storage_data_247 ^ i_input_data[550 % IN_WIDTH];
                694 / IN_WIDTH: pong_storage_data_247 <= (fillup_transition == 1'b1) ? i_input_data[694 % IN_WIDTH] : pong_storage_data_247 ^ i_input_data[694 % IN_WIDTH];
                1111 / IN_WIDTH: pong_storage_data_247 <= (fillup_transition == 1'b1) ? i_input_data[1111 % IN_WIDTH] : pong_storage_data_247 ^ i_input_data[1111 % IN_WIDTH];
                default: pong_storage_data_247 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_247;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_247 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_247;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_247 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_247;
            end
        end
    end
end

logic ping_storage_data_248;
logic pong_storage_data_248;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_248 <= 1'b0;
        pong_storage_data_248 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                320 / IN_WIDTH: ping_storage_data_248 <= (fillup_transition == 1'b1) ? i_input_data[320 % IN_WIDTH] : ping_storage_data_248 ^ i_input_data[320 % IN_WIDTH];
                418 / IN_WIDTH: ping_storage_data_248 <= (fillup_transition == 1'b1) ? i_input_data[418 % IN_WIDTH] : ping_storage_data_248 ^ i_input_data[418 % IN_WIDTH];
                551 / IN_WIDTH: ping_storage_data_248 <= (fillup_transition == 1'b1) ? i_input_data[551 % IN_WIDTH] : ping_storage_data_248 ^ i_input_data[551 % IN_WIDTH];
                695 / IN_WIDTH: ping_storage_data_248 <= (fillup_transition == 1'b1) ? i_input_data[695 % IN_WIDTH] : ping_storage_data_248 ^ i_input_data[695 % IN_WIDTH];
                1112 / IN_WIDTH: ping_storage_data_248 <= (fillup_transition == 1'b1) ? i_input_data[1112 % IN_WIDTH] : ping_storage_data_248 ^ i_input_data[1112 % IN_WIDTH];
                default: ping_storage_data_248 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_248;
                endcase
            end else begin
                case (input_count)
                320 / IN_WIDTH: pong_storage_data_248 <= (fillup_transition == 1'b1) ? i_input_data[320 % IN_WIDTH] : pong_storage_data_248 ^ i_input_data[320 % IN_WIDTH];
                418 / IN_WIDTH: pong_storage_data_248 <= (fillup_transition == 1'b1) ? i_input_data[418 % IN_WIDTH] : pong_storage_data_248 ^ i_input_data[418 % IN_WIDTH];
                551 / IN_WIDTH: pong_storage_data_248 <= (fillup_transition == 1'b1) ? i_input_data[551 % IN_WIDTH] : pong_storage_data_248 ^ i_input_data[551 % IN_WIDTH];
                695 / IN_WIDTH: pong_storage_data_248 <= (fillup_transition == 1'b1) ? i_input_data[695 % IN_WIDTH] : pong_storage_data_248 ^ i_input_data[695 % IN_WIDTH];
                1112 / IN_WIDTH: pong_storage_data_248 <= (fillup_transition == 1'b1) ? i_input_data[1112 % IN_WIDTH] : pong_storage_data_248 ^ i_input_data[1112 % IN_WIDTH];
                default: pong_storage_data_248 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_248;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_248 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_248;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_248 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_248;
            end
        end
    end
end

logic ping_storage_data_249;
logic pong_storage_data_249;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_249 <= 1'b0;
        pong_storage_data_249 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                321 / IN_WIDTH: ping_storage_data_249 <= (fillup_transition == 1'b1) ? i_input_data[321 % IN_WIDTH] : ping_storage_data_249 ^ i_input_data[321 % IN_WIDTH];
                419 / IN_WIDTH: ping_storage_data_249 <= (fillup_transition == 1'b1) ? i_input_data[419 % IN_WIDTH] : ping_storage_data_249 ^ i_input_data[419 % IN_WIDTH];
                552 / IN_WIDTH: ping_storage_data_249 <= (fillup_transition == 1'b1) ? i_input_data[552 % IN_WIDTH] : ping_storage_data_249 ^ i_input_data[552 % IN_WIDTH];
                696 / IN_WIDTH: ping_storage_data_249 <= (fillup_transition == 1'b1) ? i_input_data[696 % IN_WIDTH] : ping_storage_data_249 ^ i_input_data[696 % IN_WIDTH];
                1113 / IN_WIDTH: ping_storage_data_249 <= (fillup_transition == 1'b1) ? i_input_data[1113 % IN_WIDTH] : ping_storage_data_249 ^ i_input_data[1113 % IN_WIDTH];
                default: ping_storage_data_249 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_249;
                endcase
            end else begin
                case (input_count)
                321 / IN_WIDTH: pong_storage_data_249 <= (fillup_transition == 1'b1) ? i_input_data[321 % IN_WIDTH] : pong_storage_data_249 ^ i_input_data[321 % IN_WIDTH];
                419 / IN_WIDTH: pong_storage_data_249 <= (fillup_transition == 1'b1) ? i_input_data[419 % IN_WIDTH] : pong_storage_data_249 ^ i_input_data[419 % IN_WIDTH];
                552 / IN_WIDTH: pong_storage_data_249 <= (fillup_transition == 1'b1) ? i_input_data[552 % IN_WIDTH] : pong_storage_data_249 ^ i_input_data[552 % IN_WIDTH];
                696 / IN_WIDTH: pong_storage_data_249 <= (fillup_transition == 1'b1) ? i_input_data[696 % IN_WIDTH] : pong_storage_data_249 ^ i_input_data[696 % IN_WIDTH];
                1113 / IN_WIDTH: pong_storage_data_249 <= (fillup_transition == 1'b1) ? i_input_data[1113 % IN_WIDTH] : pong_storage_data_249 ^ i_input_data[1113 % IN_WIDTH];
                default: pong_storage_data_249 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_249;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_249 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_249;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_249 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_249;
            end
        end
    end
end

logic ping_storage_data_250;
logic pong_storage_data_250;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_250 <= 1'b0;
        pong_storage_data_250 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                322 / IN_WIDTH: ping_storage_data_250 <= (fillup_transition == 1'b1) ? i_input_data[322 % IN_WIDTH] : ping_storage_data_250 ^ i_input_data[322 % IN_WIDTH];
                420 / IN_WIDTH: ping_storage_data_250 <= (fillup_transition == 1'b1) ? i_input_data[420 % IN_WIDTH] : ping_storage_data_250 ^ i_input_data[420 % IN_WIDTH];
                553 / IN_WIDTH: ping_storage_data_250 <= (fillup_transition == 1'b1) ? i_input_data[553 % IN_WIDTH] : ping_storage_data_250 ^ i_input_data[553 % IN_WIDTH];
                697 / IN_WIDTH: ping_storage_data_250 <= (fillup_transition == 1'b1) ? i_input_data[697 % IN_WIDTH] : ping_storage_data_250 ^ i_input_data[697 % IN_WIDTH];
                1114 / IN_WIDTH: ping_storage_data_250 <= (fillup_transition == 1'b1) ? i_input_data[1114 % IN_WIDTH] : ping_storage_data_250 ^ i_input_data[1114 % IN_WIDTH];
                default: ping_storage_data_250 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_250;
                endcase
            end else begin
                case (input_count)
                322 / IN_WIDTH: pong_storage_data_250 <= (fillup_transition == 1'b1) ? i_input_data[322 % IN_WIDTH] : pong_storage_data_250 ^ i_input_data[322 % IN_WIDTH];
                420 / IN_WIDTH: pong_storage_data_250 <= (fillup_transition == 1'b1) ? i_input_data[420 % IN_WIDTH] : pong_storage_data_250 ^ i_input_data[420 % IN_WIDTH];
                553 / IN_WIDTH: pong_storage_data_250 <= (fillup_transition == 1'b1) ? i_input_data[553 % IN_WIDTH] : pong_storage_data_250 ^ i_input_data[553 % IN_WIDTH];
                697 / IN_WIDTH: pong_storage_data_250 <= (fillup_transition == 1'b1) ? i_input_data[697 % IN_WIDTH] : pong_storage_data_250 ^ i_input_data[697 % IN_WIDTH];
                1114 / IN_WIDTH: pong_storage_data_250 <= (fillup_transition == 1'b1) ? i_input_data[1114 % IN_WIDTH] : pong_storage_data_250 ^ i_input_data[1114 % IN_WIDTH];
                default: pong_storage_data_250 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_250;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_250 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_250;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_250 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_250;
            end
        end
    end
end

logic ping_storage_data_251;
logic pong_storage_data_251;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_251 <= 1'b0;
        pong_storage_data_251 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                323 / IN_WIDTH: ping_storage_data_251 <= (fillup_transition == 1'b1) ? i_input_data[323 % IN_WIDTH] : ping_storage_data_251 ^ i_input_data[323 % IN_WIDTH];
                421 / IN_WIDTH: ping_storage_data_251 <= (fillup_transition == 1'b1) ? i_input_data[421 % IN_WIDTH] : ping_storage_data_251 ^ i_input_data[421 % IN_WIDTH];
                554 / IN_WIDTH: ping_storage_data_251 <= (fillup_transition == 1'b1) ? i_input_data[554 % IN_WIDTH] : ping_storage_data_251 ^ i_input_data[554 % IN_WIDTH];
                698 / IN_WIDTH: ping_storage_data_251 <= (fillup_transition == 1'b1) ? i_input_data[698 % IN_WIDTH] : ping_storage_data_251 ^ i_input_data[698 % IN_WIDTH];
                1115 / IN_WIDTH: ping_storage_data_251 <= (fillup_transition == 1'b1) ? i_input_data[1115 % IN_WIDTH] : ping_storage_data_251 ^ i_input_data[1115 % IN_WIDTH];
                default: ping_storage_data_251 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_251;
                endcase
            end else begin
                case (input_count)
                323 / IN_WIDTH: pong_storage_data_251 <= (fillup_transition == 1'b1) ? i_input_data[323 % IN_WIDTH] : pong_storage_data_251 ^ i_input_data[323 % IN_WIDTH];
                421 / IN_WIDTH: pong_storage_data_251 <= (fillup_transition == 1'b1) ? i_input_data[421 % IN_WIDTH] : pong_storage_data_251 ^ i_input_data[421 % IN_WIDTH];
                554 / IN_WIDTH: pong_storage_data_251 <= (fillup_transition == 1'b1) ? i_input_data[554 % IN_WIDTH] : pong_storage_data_251 ^ i_input_data[554 % IN_WIDTH];
                698 / IN_WIDTH: pong_storage_data_251 <= (fillup_transition == 1'b1) ? i_input_data[698 % IN_WIDTH] : pong_storage_data_251 ^ i_input_data[698 % IN_WIDTH];
                1115 / IN_WIDTH: pong_storage_data_251 <= (fillup_transition == 1'b1) ? i_input_data[1115 % IN_WIDTH] : pong_storage_data_251 ^ i_input_data[1115 % IN_WIDTH];
                default: pong_storage_data_251 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_251;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_251 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_251;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_251 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_251;
            end
        end
    end
end

logic ping_storage_data_252;
logic pong_storage_data_252;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_252 <= 1'b0;
        pong_storage_data_252 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                324 / IN_WIDTH: ping_storage_data_252 <= (fillup_transition == 1'b1) ? i_input_data[324 % IN_WIDTH] : ping_storage_data_252 ^ i_input_data[324 % IN_WIDTH];
                422 / IN_WIDTH: ping_storage_data_252 <= (fillup_transition == 1'b1) ? i_input_data[422 % IN_WIDTH] : ping_storage_data_252 ^ i_input_data[422 % IN_WIDTH];
                555 / IN_WIDTH: ping_storage_data_252 <= (fillup_transition == 1'b1) ? i_input_data[555 % IN_WIDTH] : ping_storage_data_252 ^ i_input_data[555 % IN_WIDTH];
                699 / IN_WIDTH: ping_storage_data_252 <= (fillup_transition == 1'b1) ? i_input_data[699 % IN_WIDTH] : ping_storage_data_252 ^ i_input_data[699 % IN_WIDTH];
                1116 / IN_WIDTH: ping_storage_data_252 <= (fillup_transition == 1'b1) ? i_input_data[1116 % IN_WIDTH] : ping_storage_data_252 ^ i_input_data[1116 % IN_WIDTH];
                default: ping_storage_data_252 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_252;
                endcase
            end else begin
                case (input_count)
                324 / IN_WIDTH: pong_storage_data_252 <= (fillup_transition == 1'b1) ? i_input_data[324 % IN_WIDTH] : pong_storage_data_252 ^ i_input_data[324 % IN_WIDTH];
                422 / IN_WIDTH: pong_storage_data_252 <= (fillup_transition == 1'b1) ? i_input_data[422 % IN_WIDTH] : pong_storage_data_252 ^ i_input_data[422 % IN_WIDTH];
                555 / IN_WIDTH: pong_storage_data_252 <= (fillup_transition == 1'b1) ? i_input_data[555 % IN_WIDTH] : pong_storage_data_252 ^ i_input_data[555 % IN_WIDTH];
                699 / IN_WIDTH: pong_storage_data_252 <= (fillup_transition == 1'b1) ? i_input_data[699 % IN_WIDTH] : pong_storage_data_252 ^ i_input_data[699 % IN_WIDTH];
                1116 / IN_WIDTH: pong_storage_data_252 <= (fillup_transition == 1'b1) ? i_input_data[1116 % IN_WIDTH] : pong_storage_data_252 ^ i_input_data[1116 % IN_WIDTH];
                default: pong_storage_data_252 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_252;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_252 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_252;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_252 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_252;
            end
        end
    end
end

logic ping_storage_data_253;
logic pong_storage_data_253;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_253 <= 1'b0;
        pong_storage_data_253 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                325 / IN_WIDTH: ping_storage_data_253 <= (fillup_transition == 1'b1) ? i_input_data[325 % IN_WIDTH] : ping_storage_data_253 ^ i_input_data[325 % IN_WIDTH];
                423 / IN_WIDTH: ping_storage_data_253 <= (fillup_transition == 1'b1) ? i_input_data[423 % IN_WIDTH] : ping_storage_data_253 ^ i_input_data[423 % IN_WIDTH];
                556 / IN_WIDTH: ping_storage_data_253 <= (fillup_transition == 1'b1) ? i_input_data[556 % IN_WIDTH] : ping_storage_data_253 ^ i_input_data[556 % IN_WIDTH];
                700 / IN_WIDTH: ping_storage_data_253 <= (fillup_transition == 1'b1) ? i_input_data[700 % IN_WIDTH] : ping_storage_data_253 ^ i_input_data[700 % IN_WIDTH];
                1117 / IN_WIDTH: ping_storage_data_253 <= (fillup_transition == 1'b1) ? i_input_data[1117 % IN_WIDTH] : ping_storage_data_253 ^ i_input_data[1117 % IN_WIDTH];
                default: ping_storage_data_253 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_253;
                endcase
            end else begin
                case (input_count)
                325 / IN_WIDTH: pong_storage_data_253 <= (fillup_transition == 1'b1) ? i_input_data[325 % IN_WIDTH] : pong_storage_data_253 ^ i_input_data[325 % IN_WIDTH];
                423 / IN_WIDTH: pong_storage_data_253 <= (fillup_transition == 1'b1) ? i_input_data[423 % IN_WIDTH] : pong_storage_data_253 ^ i_input_data[423 % IN_WIDTH];
                556 / IN_WIDTH: pong_storage_data_253 <= (fillup_transition == 1'b1) ? i_input_data[556 % IN_WIDTH] : pong_storage_data_253 ^ i_input_data[556 % IN_WIDTH];
                700 / IN_WIDTH: pong_storage_data_253 <= (fillup_transition == 1'b1) ? i_input_data[700 % IN_WIDTH] : pong_storage_data_253 ^ i_input_data[700 % IN_WIDTH];
                1117 / IN_WIDTH: pong_storage_data_253 <= (fillup_transition == 1'b1) ? i_input_data[1117 % IN_WIDTH] : pong_storage_data_253 ^ i_input_data[1117 % IN_WIDTH];
                default: pong_storage_data_253 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_253;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_253 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_253;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_253 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_253;
            end
        end
    end
end

logic ping_storage_data_254;
logic pong_storage_data_254;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_254 <= 1'b0;
        pong_storage_data_254 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                326 / IN_WIDTH: ping_storage_data_254 <= (fillup_transition == 1'b1) ? i_input_data[326 % IN_WIDTH] : ping_storage_data_254 ^ i_input_data[326 % IN_WIDTH];
                424 / IN_WIDTH: ping_storage_data_254 <= (fillup_transition == 1'b1) ? i_input_data[424 % IN_WIDTH] : ping_storage_data_254 ^ i_input_data[424 % IN_WIDTH];
                557 / IN_WIDTH: ping_storage_data_254 <= (fillup_transition == 1'b1) ? i_input_data[557 % IN_WIDTH] : ping_storage_data_254 ^ i_input_data[557 % IN_WIDTH];
                701 / IN_WIDTH: ping_storage_data_254 <= (fillup_transition == 1'b1) ? i_input_data[701 % IN_WIDTH] : ping_storage_data_254 ^ i_input_data[701 % IN_WIDTH];
                1118 / IN_WIDTH: ping_storage_data_254 <= (fillup_transition == 1'b1) ? i_input_data[1118 % IN_WIDTH] : ping_storage_data_254 ^ i_input_data[1118 % IN_WIDTH];
                default: ping_storage_data_254 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_254;
                endcase
            end else begin
                case (input_count)
                326 / IN_WIDTH: pong_storage_data_254 <= (fillup_transition == 1'b1) ? i_input_data[326 % IN_WIDTH] : pong_storage_data_254 ^ i_input_data[326 % IN_WIDTH];
                424 / IN_WIDTH: pong_storage_data_254 <= (fillup_transition == 1'b1) ? i_input_data[424 % IN_WIDTH] : pong_storage_data_254 ^ i_input_data[424 % IN_WIDTH];
                557 / IN_WIDTH: pong_storage_data_254 <= (fillup_transition == 1'b1) ? i_input_data[557 % IN_WIDTH] : pong_storage_data_254 ^ i_input_data[557 % IN_WIDTH];
                701 / IN_WIDTH: pong_storage_data_254 <= (fillup_transition == 1'b1) ? i_input_data[701 % IN_WIDTH] : pong_storage_data_254 ^ i_input_data[701 % IN_WIDTH];
                1118 / IN_WIDTH: pong_storage_data_254 <= (fillup_transition == 1'b1) ? i_input_data[1118 % IN_WIDTH] : pong_storage_data_254 ^ i_input_data[1118 % IN_WIDTH];
                default: pong_storage_data_254 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_254;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_254 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_254;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_254 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_254;
            end
        end
    end
end

logic ping_storage_data_255;
logic pong_storage_data_255;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_255 <= 1'b0;
        pong_storage_data_255 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                327 / IN_WIDTH: ping_storage_data_255 <= (fillup_transition == 1'b1) ? i_input_data[327 % IN_WIDTH] : ping_storage_data_255 ^ i_input_data[327 % IN_WIDTH];
                425 / IN_WIDTH: ping_storage_data_255 <= (fillup_transition == 1'b1) ? i_input_data[425 % IN_WIDTH] : ping_storage_data_255 ^ i_input_data[425 % IN_WIDTH];
                558 / IN_WIDTH: ping_storage_data_255 <= (fillup_transition == 1'b1) ? i_input_data[558 % IN_WIDTH] : ping_storage_data_255 ^ i_input_data[558 % IN_WIDTH];
                702 / IN_WIDTH: ping_storage_data_255 <= (fillup_transition == 1'b1) ? i_input_data[702 % IN_WIDTH] : ping_storage_data_255 ^ i_input_data[702 % IN_WIDTH];
                1119 / IN_WIDTH: ping_storage_data_255 <= (fillup_transition == 1'b1) ? i_input_data[1119 % IN_WIDTH] : ping_storage_data_255 ^ i_input_data[1119 % IN_WIDTH];
                default: ping_storage_data_255 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_255;
                endcase
            end else begin
                case (input_count)
                327 / IN_WIDTH: pong_storage_data_255 <= (fillup_transition == 1'b1) ? i_input_data[327 % IN_WIDTH] : pong_storage_data_255 ^ i_input_data[327 % IN_WIDTH];
                425 / IN_WIDTH: pong_storage_data_255 <= (fillup_transition == 1'b1) ? i_input_data[425 % IN_WIDTH] : pong_storage_data_255 ^ i_input_data[425 % IN_WIDTH];
                558 / IN_WIDTH: pong_storage_data_255 <= (fillup_transition == 1'b1) ? i_input_data[558 % IN_WIDTH] : pong_storage_data_255 ^ i_input_data[558 % IN_WIDTH];
                702 / IN_WIDTH: pong_storage_data_255 <= (fillup_transition == 1'b1) ? i_input_data[702 % IN_WIDTH] : pong_storage_data_255 ^ i_input_data[702 % IN_WIDTH];
                1119 / IN_WIDTH: pong_storage_data_255 <= (fillup_transition == 1'b1) ? i_input_data[1119 % IN_WIDTH] : pong_storage_data_255 ^ i_input_data[1119 % IN_WIDTH];
                default: pong_storage_data_255 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_255;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_255 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_255;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_255 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_255;
            end
        end
    end
end

logic ping_storage_data_256;
logic pong_storage_data_256;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_256 <= 1'b0;
        pong_storage_data_256 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                328 / IN_WIDTH: ping_storage_data_256 <= (fillup_transition == 1'b1) ? i_input_data[328 % IN_WIDTH] : ping_storage_data_256 ^ i_input_data[328 % IN_WIDTH];
                426 / IN_WIDTH: ping_storage_data_256 <= (fillup_transition == 1'b1) ? i_input_data[426 % IN_WIDTH] : ping_storage_data_256 ^ i_input_data[426 % IN_WIDTH];
                559 / IN_WIDTH: ping_storage_data_256 <= (fillup_transition == 1'b1) ? i_input_data[559 % IN_WIDTH] : ping_storage_data_256 ^ i_input_data[559 % IN_WIDTH];
                703 / IN_WIDTH: ping_storage_data_256 <= (fillup_transition == 1'b1) ? i_input_data[703 % IN_WIDTH] : ping_storage_data_256 ^ i_input_data[703 % IN_WIDTH];
                1120 / IN_WIDTH: ping_storage_data_256 <= (fillup_transition == 1'b1) ? i_input_data[1120 % IN_WIDTH] : ping_storage_data_256 ^ i_input_data[1120 % IN_WIDTH];
                default: ping_storage_data_256 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_256;
                endcase
            end else begin
                case (input_count)
                328 / IN_WIDTH: pong_storage_data_256 <= (fillup_transition == 1'b1) ? i_input_data[328 % IN_WIDTH] : pong_storage_data_256 ^ i_input_data[328 % IN_WIDTH];
                426 / IN_WIDTH: pong_storage_data_256 <= (fillup_transition == 1'b1) ? i_input_data[426 % IN_WIDTH] : pong_storage_data_256 ^ i_input_data[426 % IN_WIDTH];
                559 / IN_WIDTH: pong_storage_data_256 <= (fillup_transition == 1'b1) ? i_input_data[559 % IN_WIDTH] : pong_storage_data_256 ^ i_input_data[559 % IN_WIDTH];
                703 / IN_WIDTH: pong_storage_data_256 <= (fillup_transition == 1'b1) ? i_input_data[703 % IN_WIDTH] : pong_storage_data_256 ^ i_input_data[703 % IN_WIDTH];
                1120 / IN_WIDTH: pong_storage_data_256 <= (fillup_transition == 1'b1) ? i_input_data[1120 % IN_WIDTH] : pong_storage_data_256 ^ i_input_data[1120 % IN_WIDTH];
                default: pong_storage_data_256 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_256;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_256 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_256;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_256 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_256;
            end
        end
    end
end

logic ping_storage_data_257;
logic pong_storage_data_257;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_257 <= 1'b0;
        pong_storage_data_257 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                329 / IN_WIDTH: ping_storage_data_257 <= (fillup_transition == 1'b1) ? i_input_data[329 % IN_WIDTH] : ping_storage_data_257 ^ i_input_data[329 % IN_WIDTH];
                427 / IN_WIDTH: ping_storage_data_257 <= (fillup_transition == 1'b1) ? i_input_data[427 % IN_WIDTH] : ping_storage_data_257 ^ i_input_data[427 % IN_WIDTH];
                560 / IN_WIDTH: ping_storage_data_257 <= (fillup_transition == 1'b1) ? i_input_data[560 % IN_WIDTH] : ping_storage_data_257 ^ i_input_data[560 % IN_WIDTH];
                704 / IN_WIDTH: ping_storage_data_257 <= (fillup_transition == 1'b1) ? i_input_data[704 % IN_WIDTH] : ping_storage_data_257 ^ i_input_data[704 % IN_WIDTH];
                1121 / IN_WIDTH: ping_storage_data_257 <= (fillup_transition == 1'b1) ? i_input_data[1121 % IN_WIDTH] : ping_storage_data_257 ^ i_input_data[1121 % IN_WIDTH];
                default: ping_storage_data_257 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_257;
                endcase
            end else begin
                case (input_count)
                329 / IN_WIDTH: pong_storage_data_257 <= (fillup_transition == 1'b1) ? i_input_data[329 % IN_WIDTH] : pong_storage_data_257 ^ i_input_data[329 % IN_WIDTH];
                427 / IN_WIDTH: pong_storage_data_257 <= (fillup_transition == 1'b1) ? i_input_data[427 % IN_WIDTH] : pong_storage_data_257 ^ i_input_data[427 % IN_WIDTH];
                560 / IN_WIDTH: pong_storage_data_257 <= (fillup_transition == 1'b1) ? i_input_data[560 % IN_WIDTH] : pong_storage_data_257 ^ i_input_data[560 % IN_WIDTH];
                704 / IN_WIDTH: pong_storage_data_257 <= (fillup_transition == 1'b1) ? i_input_data[704 % IN_WIDTH] : pong_storage_data_257 ^ i_input_data[704 % IN_WIDTH];
                1121 / IN_WIDTH: pong_storage_data_257 <= (fillup_transition == 1'b1) ? i_input_data[1121 % IN_WIDTH] : pong_storage_data_257 ^ i_input_data[1121 % IN_WIDTH];
                default: pong_storage_data_257 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_257;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_257 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_257;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_257 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_257;
            end
        end
    end
end

logic ping_storage_data_258;
logic pong_storage_data_258;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_258 <= 1'b0;
        pong_storage_data_258 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                330 / IN_WIDTH: ping_storage_data_258 <= (fillup_transition == 1'b1) ? i_input_data[330 % IN_WIDTH] : ping_storage_data_258 ^ i_input_data[330 % IN_WIDTH];
                428 / IN_WIDTH: ping_storage_data_258 <= (fillup_transition == 1'b1) ? i_input_data[428 % IN_WIDTH] : ping_storage_data_258 ^ i_input_data[428 % IN_WIDTH];
                561 / IN_WIDTH: ping_storage_data_258 <= (fillup_transition == 1'b1) ? i_input_data[561 % IN_WIDTH] : ping_storage_data_258 ^ i_input_data[561 % IN_WIDTH];
                705 / IN_WIDTH: ping_storage_data_258 <= (fillup_transition == 1'b1) ? i_input_data[705 % IN_WIDTH] : ping_storage_data_258 ^ i_input_data[705 % IN_WIDTH];
                1122 / IN_WIDTH: ping_storage_data_258 <= (fillup_transition == 1'b1) ? i_input_data[1122 % IN_WIDTH] : ping_storage_data_258 ^ i_input_data[1122 % IN_WIDTH];
                default: ping_storage_data_258 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_258;
                endcase
            end else begin
                case (input_count)
                330 / IN_WIDTH: pong_storage_data_258 <= (fillup_transition == 1'b1) ? i_input_data[330 % IN_WIDTH] : pong_storage_data_258 ^ i_input_data[330 % IN_WIDTH];
                428 / IN_WIDTH: pong_storage_data_258 <= (fillup_transition == 1'b1) ? i_input_data[428 % IN_WIDTH] : pong_storage_data_258 ^ i_input_data[428 % IN_WIDTH];
                561 / IN_WIDTH: pong_storage_data_258 <= (fillup_transition == 1'b1) ? i_input_data[561 % IN_WIDTH] : pong_storage_data_258 ^ i_input_data[561 % IN_WIDTH];
                705 / IN_WIDTH: pong_storage_data_258 <= (fillup_transition == 1'b1) ? i_input_data[705 % IN_WIDTH] : pong_storage_data_258 ^ i_input_data[705 % IN_WIDTH];
                1122 / IN_WIDTH: pong_storage_data_258 <= (fillup_transition == 1'b1) ? i_input_data[1122 % IN_WIDTH] : pong_storage_data_258 ^ i_input_data[1122 % IN_WIDTH];
                default: pong_storage_data_258 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_258;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_258 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_258;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_258 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_258;
            end
        end
    end
end

logic ping_storage_data_259;
logic pong_storage_data_259;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_259 <= 1'b0;
        pong_storage_data_259 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                331 / IN_WIDTH: ping_storage_data_259 <= (fillup_transition == 1'b1) ? i_input_data[331 % IN_WIDTH] : ping_storage_data_259 ^ i_input_data[331 % IN_WIDTH];
                429 / IN_WIDTH: ping_storage_data_259 <= (fillup_transition == 1'b1) ? i_input_data[429 % IN_WIDTH] : ping_storage_data_259 ^ i_input_data[429 % IN_WIDTH];
                562 / IN_WIDTH: ping_storage_data_259 <= (fillup_transition == 1'b1) ? i_input_data[562 % IN_WIDTH] : ping_storage_data_259 ^ i_input_data[562 % IN_WIDTH];
                706 / IN_WIDTH: ping_storage_data_259 <= (fillup_transition == 1'b1) ? i_input_data[706 % IN_WIDTH] : ping_storage_data_259 ^ i_input_data[706 % IN_WIDTH];
                1123 / IN_WIDTH: ping_storage_data_259 <= (fillup_transition == 1'b1) ? i_input_data[1123 % IN_WIDTH] : ping_storage_data_259 ^ i_input_data[1123 % IN_WIDTH];
                default: ping_storage_data_259 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_259;
                endcase
            end else begin
                case (input_count)
                331 / IN_WIDTH: pong_storage_data_259 <= (fillup_transition == 1'b1) ? i_input_data[331 % IN_WIDTH] : pong_storage_data_259 ^ i_input_data[331 % IN_WIDTH];
                429 / IN_WIDTH: pong_storage_data_259 <= (fillup_transition == 1'b1) ? i_input_data[429 % IN_WIDTH] : pong_storage_data_259 ^ i_input_data[429 % IN_WIDTH];
                562 / IN_WIDTH: pong_storage_data_259 <= (fillup_transition == 1'b1) ? i_input_data[562 % IN_WIDTH] : pong_storage_data_259 ^ i_input_data[562 % IN_WIDTH];
                706 / IN_WIDTH: pong_storage_data_259 <= (fillup_transition == 1'b1) ? i_input_data[706 % IN_WIDTH] : pong_storage_data_259 ^ i_input_data[706 % IN_WIDTH];
                1123 / IN_WIDTH: pong_storage_data_259 <= (fillup_transition == 1'b1) ? i_input_data[1123 % IN_WIDTH] : pong_storage_data_259 ^ i_input_data[1123 % IN_WIDTH];
                default: pong_storage_data_259 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_259;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_259 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_259;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_259 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_259;
            end
        end
    end
end

logic ping_storage_data_260;
logic pong_storage_data_260;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_260 <= 1'b0;
        pong_storage_data_260 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                332 / IN_WIDTH: ping_storage_data_260 <= (fillup_transition == 1'b1) ? i_input_data[332 % IN_WIDTH] : ping_storage_data_260 ^ i_input_data[332 % IN_WIDTH];
                430 / IN_WIDTH: ping_storage_data_260 <= (fillup_transition == 1'b1) ? i_input_data[430 % IN_WIDTH] : ping_storage_data_260 ^ i_input_data[430 % IN_WIDTH];
                563 / IN_WIDTH: ping_storage_data_260 <= (fillup_transition == 1'b1) ? i_input_data[563 % IN_WIDTH] : ping_storage_data_260 ^ i_input_data[563 % IN_WIDTH];
                707 / IN_WIDTH: ping_storage_data_260 <= (fillup_transition == 1'b1) ? i_input_data[707 % IN_WIDTH] : ping_storage_data_260 ^ i_input_data[707 % IN_WIDTH];
                1124 / IN_WIDTH: ping_storage_data_260 <= (fillup_transition == 1'b1) ? i_input_data[1124 % IN_WIDTH] : ping_storage_data_260 ^ i_input_data[1124 % IN_WIDTH];
                default: ping_storage_data_260 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_260;
                endcase
            end else begin
                case (input_count)
                332 / IN_WIDTH: pong_storage_data_260 <= (fillup_transition == 1'b1) ? i_input_data[332 % IN_WIDTH] : pong_storage_data_260 ^ i_input_data[332 % IN_WIDTH];
                430 / IN_WIDTH: pong_storage_data_260 <= (fillup_transition == 1'b1) ? i_input_data[430 % IN_WIDTH] : pong_storage_data_260 ^ i_input_data[430 % IN_WIDTH];
                563 / IN_WIDTH: pong_storage_data_260 <= (fillup_transition == 1'b1) ? i_input_data[563 % IN_WIDTH] : pong_storage_data_260 ^ i_input_data[563 % IN_WIDTH];
                707 / IN_WIDTH: pong_storage_data_260 <= (fillup_transition == 1'b1) ? i_input_data[707 % IN_WIDTH] : pong_storage_data_260 ^ i_input_data[707 % IN_WIDTH];
                1124 / IN_WIDTH: pong_storage_data_260 <= (fillup_transition == 1'b1) ? i_input_data[1124 % IN_WIDTH] : pong_storage_data_260 ^ i_input_data[1124 % IN_WIDTH];
                default: pong_storage_data_260 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_260;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_260 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_260;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_260 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_260;
            end
        end
    end
end

logic ping_storage_data_261;
logic pong_storage_data_261;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_261 <= 1'b0;
        pong_storage_data_261 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                333 / IN_WIDTH: ping_storage_data_261 <= (fillup_transition == 1'b1) ? i_input_data[333 % IN_WIDTH] : ping_storage_data_261 ^ i_input_data[333 % IN_WIDTH];
                431 / IN_WIDTH: ping_storage_data_261 <= (fillup_transition == 1'b1) ? i_input_data[431 % IN_WIDTH] : ping_storage_data_261 ^ i_input_data[431 % IN_WIDTH];
                564 / IN_WIDTH: ping_storage_data_261 <= (fillup_transition == 1'b1) ? i_input_data[564 % IN_WIDTH] : ping_storage_data_261 ^ i_input_data[564 % IN_WIDTH];
                708 / IN_WIDTH: ping_storage_data_261 <= (fillup_transition == 1'b1) ? i_input_data[708 % IN_WIDTH] : ping_storage_data_261 ^ i_input_data[708 % IN_WIDTH];
                1125 / IN_WIDTH: ping_storage_data_261 <= (fillup_transition == 1'b1) ? i_input_data[1125 % IN_WIDTH] : ping_storage_data_261 ^ i_input_data[1125 % IN_WIDTH];
                default: ping_storage_data_261 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_261;
                endcase
            end else begin
                case (input_count)
                333 / IN_WIDTH: pong_storage_data_261 <= (fillup_transition == 1'b1) ? i_input_data[333 % IN_WIDTH] : pong_storage_data_261 ^ i_input_data[333 % IN_WIDTH];
                431 / IN_WIDTH: pong_storage_data_261 <= (fillup_transition == 1'b1) ? i_input_data[431 % IN_WIDTH] : pong_storage_data_261 ^ i_input_data[431 % IN_WIDTH];
                564 / IN_WIDTH: pong_storage_data_261 <= (fillup_transition == 1'b1) ? i_input_data[564 % IN_WIDTH] : pong_storage_data_261 ^ i_input_data[564 % IN_WIDTH];
                708 / IN_WIDTH: pong_storage_data_261 <= (fillup_transition == 1'b1) ? i_input_data[708 % IN_WIDTH] : pong_storage_data_261 ^ i_input_data[708 % IN_WIDTH];
                1125 / IN_WIDTH: pong_storage_data_261 <= (fillup_transition == 1'b1) ? i_input_data[1125 % IN_WIDTH] : pong_storage_data_261 ^ i_input_data[1125 % IN_WIDTH];
                default: pong_storage_data_261 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_261;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_261 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_261;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_261 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_261;
            end
        end
    end
end

logic ping_storage_data_262;
logic pong_storage_data_262;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_262 <= 1'b0;
        pong_storage_data_262 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                334 / IN_WIDTH: ping_storage_data_262 <= (fillup_transition == 1'b1) ? i_input_data[334 % IN_WIDTH] : ping_storage_data_262 ^ i_input_data[334 % IN_WIDTH];
                432 / IN_WIDTH: ping_storage_data_262 <= (fillup_transition == 1'b1) ? i_input_data[432 % IN_WIDTH] : ping_storage_data_262 ^ i_input_data[432 % IN_WIDTH];
                565 / IN_WIDTH: ping_storage_data_262 <= (fillup_transition == 1'b1) ? i_input_data[565 % IN_WIDTH] : ping_storage_data_262 ^ i_input_data[565 % IN_WIDTH];
                709 / IN_WIDTH: ping_storage_data_262 <= (fillup_transition == 1'b1) ? i_input_data[709 % IN_WIDTH] : ping_storage_data_262 ^ i_input_data[709 % IN_WIDTH];
                1126 / IN_WIDTH: ping_storage_data_262 <= (fillup_transition == 1'b1) ? i_input_data[1126 % IN_WIDTH] : ping_storage_data_262 ^ i_input_data[1126 % IN_WIDTH];
                default: ping_storage_data_262 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_262;
                endcase
            end else begin
                case (input_count)
                334 / IN_WIDTH: pong_storage_data_262 <= (fillup_transition == 1'b1) ? i_input_data[334 % IN_WIDTH] : pong_storage_data_262 ^ i_input_data[334 % IN_WIDTH];
                432 / IN_WIDTH: pong_storage_data_262 <= (fillup_transition == 1'b1) ? i_input_data[432 % IN_WIDTH] : pong_storage_data_262 ^ i_input_data[432 % IN_WIDTH];
                565 / IN_WIDTH: pong_storage_data_262 <= (fillup_transition == 1'b1) ? i_input_data[565 % IN_WIDTH] : pong_storage_data_262 ^ i_input_data[565 % IN_WIDTH];
                709 / IN_WIDTH: pong_storage_data_262 <= (fillup_transition == 1'b1) ? i_input_data[709 % IN_WIDTH] : pong_storage_data_262 ^ i_input_data[709 % IN_WIDTH];
                1126 / IN_WIDTH: pong_storage_data_262 <= (fillup_transition == 1'b1) ? i_input_data[1126 % IN_WIDTH] : pong_storage_data_262 ^ i_input_data[1126 % IN_WIDTH];
                default: pong_storage_data_262 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_262;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_262 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_262;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_262 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_262;
            end
        end
    end
end

logic ping_storage_data_263;
logic pong_storage_data_263;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_263 <= 1'b0;
        pong_storage_data_263 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                335 / IN_WIDTH: ping_storage_data_263 <= (fillup_transition == 1'b1) ? i_input_data[335 % IN_WIDTH] : ping_storage_data_263 ^ i_input_data[335 % IN_WIDTH];
                433 / IN_WIDTH: ping_storage_data_263 <= (fillup_transition == 1'b1) ? i_input_data[433 % IN_WIDTH] : ping_storage_data_263 ^ i_input_data[433 % IN_WIDTH];
                566 / IN_WIDTH: ping_storage_data_263 <= (fillup_transition == 1'b1) ? i_input_data[566 % IN_WIDTH] : ping_storage_data_263 ^ i_input_data[566 % IN_WIDTH];
                710 / IN_WIDTH: ping_storage_data_263 <= (fillup_transition == 1'b1) ? i_input_data[710 % IN_WIDTH] : ping_storage_data_263 ^ i_input_data[710 % IN_WIDTH];
                1127 / IN_WIDTH: ping_storage_data_263 <= (fillup_transition == 1'b1) ? i_input_data[1127 % IN_WIDTH] : ping_storage_data_263 ^ i_input_data[1127 % IN_WIDTH];
                default: ping_storage_data_263 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_263;
                endcase
            end else begin
                case (input_count)
                335 / IN_WIDTH: pong_storage_data_263 <= (fillup_transition == 1'b1) ? i_input_data[335 % IN_WIDTH] : pong_storage_data_263 ^ i_input_data[335 % IN_WIDTH];
                433 / IN_WIDTH: pong_storage_data_263 <= (fillup_transition == 1'b1) ? i_input_data[433 % IN_WIDTH] : pong_storage_data_263 ^ i_input_data[433 % IN_WIDTH];
                566 / IN_WIDTH: pong_storage_data_263 <= (fillup_transition == 1'b1) ? i_input_data[566 % IN_WIDTH] : pong_storage_data_263 ^ i_input_data[566 % IN_WIDTH];
                710 / IN_WIDTH: pong_storage_data_263 <= (fillup_transition == 1'b1) ? i_input_data[710 % IN_WIDTH] : pong_storage_data_263 ^ i_input_data[710 % IN_WIDTH];
                1127 / IN_WIDTH: pong_storage_data_263 <= (fillup_transition == 1'b1) ? i_input_data[1127 % IN_WIDTH] : pong_storage_data_263 ^ i_input_data[1127 % IN_WIDTH];
                default: pong_storage_data_263 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_263;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_263 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_263;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_263 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_263;
            end
        end
    end
end

logic ping_storage_data_264;
logic pong_storage_data_264;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_264 <= 1'b0;
        pong_storage_data_264 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                336 / IN_WIDTH: ping_storage_data_264 <= (fillup_transition == 1'b1) ? i_input_data[336 % IN_WIDTH] : ping_storage_data_264 ^ i_input_data[336 % IN_WIDTH];
                434 / IN_WIDTH: ping_storage_data_264 <= (fillup_transition == 1'b1) ? i_input_data[434 % IN_WIDTH] : ping_storage_data_264 ^ i_input_data[434 % IN_WIDTH];
                567 / IN_WIDTH: ping_storage_data_264 <= (fillup_transition == 1'b1) ? i_input_data[567 % IN_WIDTH] : ping_storage_data_264 ^ i_input_data[567 % IN_WIDTH];
                711 / IN_WIDTH: ping_storage_data_264 <= (fillup_transition == 1'b1) ? i_input_data[711 % IN_WIDTH] : ping_storage_data_264 ^ i_input_data[711 % IN_WIDTH];
                1128 / IN_WIDTH: ping_storage_data_264 <= (fillup_transition == 1'b1) ? i_input_data[1128 % IN_WIDTH] : ping_storage_data_264 ^ i_input_data[1128 % IN_WIDTH];
                default: ping_storage_data_264 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_264;
                endcase
            end else begin
                case (input_count)
                336 / IN_WIDTH: pong_storage_data_264 <= (fillup_transition == 1'b1) ? i_input_data[336 % IN_WIDTH] : pong_storage_data_264 ^ i_input_data[336 % IN_WIDTH];
                434 / IN_WIDTH: pong_storage_data_264 <= (fillup_transition == 1'b1) ? i_input_data[434 % IN_WIDTH] : pong_storage_data_264 ^ i_input_data[434 % IN_WIDTH];
                567 / IN_WIDTH: pong_storage_data_264 <= (fillup_transition == 1'b1) ? i_input_data[567 % IN_WIDTH] : pong_storage_data_264 ^ i_input_data[567 % IN_WIDTH];
                711 / IN_WIDTH: pong_storage_data_264 <= (fillup_transition == 1'b1) ? i_input_data[711 % IN_WIDTH] : pong_storage_data_264 ^ i_input_data[711 % IN_WIDTH];
                1128 / IN_WIDTH: pong_storage_data_264 <= (fillup_transition == 1'b1) ? i_input_data[1128 % IN_WIDTH] : pong_storage_data_264 ^ i_input_data[1128 % IN_WIDTH];
                default: pong_storage_data_264 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_264;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_264 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_264;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_264 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_264;
            end
        end
    end
end

logic ping_storage_data_265;
logic pong_storage_data_265;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_265 <= 1'b0;
        pong_storage_data_265 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                337 / IN_WIDTH: ping_storage_data_265 <= (fillup_transition == 1'b1) ? i_input_data[337 % IN_WIDTH] : ping_storage_data_265 ^ i_input_data[337 % IN_WIDTH];
                435 / IN_WIDTH: ping_storage_data_265 <= (fillup_transition == 1'b1) ? i_input_data[435 % IN_WIDTH] : ping_storage_data_265 ^ i_input_data[435 % IN_WIDTH];
                568 / IN_WIDTH: ping_storage_data_265 <= (fillup_transition == 1'b1) ? i_input_data[568 % IN_WIDTH] : ping_storage_data_265 ^ i_input_data[568 % IN_WIDTH];
                712 / IN_WIDTH: ping_storage_data_265 <= (fillup_transition == 1'b1) ? i_input_data[712 % IN_WIDTH] : ping_storage_data_265 ^ i_input_data[712 % IN_WIDTH];
                1129 / IN_WIDTH: ping_storage_data_265 <= (fillup_transition == 1'b1) ? i_input_data[1129 % IN_WIDTH] : ping_storage_data_265 ^ i_input_data[1129 % IN_WIDTH];
                default: ping_storage_data_265 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_265;
                endcase
            end else begin
                case (input_count)
                337 / IN_WIDTH: pong_storage_data_265 <= (fillup_transition == 1'b1) ? i_input_data[337 % IN_WIDTH] : pong_storage_data_265 ^ i_input_data[337 % IN_WIDTH];
                435 / IN_WIDTH: pong_storage_data_265 <= (fillup_transition == 1'b1) ? i_input_data[435 % IN_WIDTH] : pong_storage_data_265 ^ i_input_data[435 % IN_WIDTH];
                568 / IN_WIDTH: pong_storage_data_265 <= (fillup_transition == 1'b1) ? i_input_data[568 % IN_WIDTH] : pong_storage_data_265 ^ i_input_data[568 % IN_WIDTH];
                712 / IN_WIDTH: pong_storage_data_265 <= (fillup_transition == 1'b1) ? i_input_data[712 % IN_WIDTH] : pong_storage_data_265 ^ i_input_data[712 % IN_WIDTH];
                1129 / IN_WIDTH: pong_storage_data_265 <= (fillup_transition == 1'b1) ? i_input_data[1129 % IN_WIDTH] : pong_storage_data_265 ^ i_input_data[1129 % IN_WIDTH];
                default: pong_storage_data_265 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_265;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_265 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_265;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_265 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_265;
            end
        end
    end
end

logic ping_storage_data_266;
logic pong_storage_data_266;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_266 <= 1'b0;
        pong_storage_data_266 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                338 / IN_WIDTH: ping_storage_data_266 <= (fillup_transition == 1'b1) ? i_input_data[338 % IN_WIDTH] : ping_storage_data_266 ^ i_input_data[338 % IN_WIDTH];
                436 / IN_WIDTH: ping_storage_data_266 <= (fillup_transition == 1'b1) ? i_input_data[436 % IN_WIDTH] : ping_storage_data_266 ^ i_input_data[436 % IN_WIDTH];
                569 / IN_WIDTH: ping_storage_data_266 <= (fillup_transition == 1'b1) ? i_input_data[569 % IN_WIDTH] : ping_storage_data_266 ^ i_input_data[569 % IN_WIDTH];
                713 / IN_WIDTH: ping_storage_data_266 <= (fillup_transition == 1'b1) ? i_input_data[713 % IN_WIDTH] : ping_storage_data_266 ^ i_input_data[713 % IN_WIDTH];
                1130 / IN_WIDTH: ping_storage_data_266 <= (fillup_transition == 1'b1) ? i_input_data[1130 % IN_WIDTH] : ping_storage_data_266 ^ i_input_data[1130 % IN_WIDTH];
                default: ping_storage_data_266 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_266;
                endcase
            end else begin
                case (input_count)
                338 / IN_WIDTH: pong_storage_data_266 <= (fillup_transition == 1'b1) ? i_input_data[338 % IN_WIDTH] : pong_storage_data_266 ^ i_input_data[338 % IN_WIDTH];
                436 / IN_WIDTH: pong_storage_data_266 <= (fillup_transition == 1'b1) ? i_input_data[436 % IN_WIDTH] : pong_storage_data_266 ^ i_input_data[436 % IN_WIDTH];
                569 / IN_WIDTH: pong_storage_data_266 <= (fillup_transition == 1'b1) ? i_input_data[569 % IN_WIDTH] : pong_storage_data_266 ^ i_input_data[569 % IN_WIDTH];
                713 / IN_WIDTH: pong_storage_data_266 <= (fillup_transition == 1'b1) ? i_input_data[713 % IN_WIDTH] : pong_storage_data_266 ^ i_input_data[713 % IN_WIDTH];
                1130 / IN_WIDTH: pong_storage_data_266 <= (fillup_transition == 1'b1) ? i_input_data[1130 % IN_WIDTH] : pong_storage_data_266 ^ i_input_data[1130 % IN_WIDTH];
                default: pong_storage_data_266 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_266;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_266 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_266;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_266 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_266;
            end
        end
    end
end

logic ping_storage_data_267;
logic pong_storage_data_267;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_267 <= 1'b0;
        pong_storage_data_267 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                339 / IN_WIDTH: ping_storage_data_267 <= (fillup_transition == 1'b1) ? i_input_data[339 % IN_WIDTH] : ping_storage_data_267 ^ i_input_data[339 % IN_WIDTH];
                437 / IN_WIDTH: ping_storage_data_267 <= (fillup_transition == 1'b1) ? i_input_data[437 % IN_WIDTH] : ping_storage_data_267 ^ i_input_data[437 % IN_WIDTH];
                570 / IN_WIDTH: ping_storage_data_267 <= (fillup_transition == 1'b1) ? i_input_data[570 % IN_WIDTH] : ping_storage_data_267 ^ i_input_data[570 % IN_WIDTH];
                714 / IN_WIDTH: ping_storage_data_267 <= (fillup_transition == 1'b1) ? i_input_data[714 % IN_WIDTH] : ping_storage_data_267 ^ i_input_data[714 % IN_WIDTH];
                1131 / IN_WIDTH: ping_storage_data_267 <= (fillup_transition == 1'b1) ? i_input_data[1131 % IN_WIDTH] : ping_storage_data_267 ^ i_input_data[1131 % IN_WIDTH];
                default: ping_storage_data_267 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_267;
                endcase
            end else begin
                case (input_count)
                339 / IN_WIDTH: pong_storage_data_267 <= (fillup_transition == 1'b1) ? i_input_data[339 % IN_WIDTH] : pong_storage_data_267 ^ i_input_data[339 % IN_WIDTH];
                437 / IN_WIDTH: pong_storage_data_267 <= (fillup_transition == 1'b1) ? i_input_data[437 % IN_WIDTH] : pong_storage_data_267 ^ i_input_data[437 % IN_WIDTH];
                570 / IN_WIDTH: pong_storage_data_267 <= (fillup_transition == 1'b1) ? i_input_data[570 % IN_WIDTH] : pong_storage_data_267 ^ i_input_data[570 % IN_WIDTH];
                714 / IN_WIDTH: pong_storage_data_267 <= (fillup_transition == 1'b1) ? i_input_data[714 % IN_WIDTH] : pong_storage_data_267 ^ i_input_data[714 % IN_WIDTH];
                1131 / IN_WIDTH: pong_storage_data_267 <= (fillup_transition == 1'b1) ? i_input_data[1131 % IN_WIDTH] : pong_storage_data_267 ^ i_input_data[1131 % IN_WIDTH];
                default: pong_storage_data_267 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_267;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_267 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_267;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_267 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_267;
            end
        end
    end
end

logic ping_storage_data_268;
logic pong_storage_data_268;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_268 <= 1'b0;
        pong_storage_data_268 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                340 / IN_WIDTH: ping_storage_data_268 <= (fillup_transition == 1'b1) ? i_input_data[340 % IN_WIDTH] : ping_storage_data_268 ^ i_input_data[340 % IN_WIDTH];
                438 / IN_WIDTH: ping_storage_data_268 <= (fillup_transition == 1'b1) ? i_input_data[438 % IN_WIDTH] : ping_storage_data_268 ^ i_input_data[438 % IN_WIDTH];
                571 / IN_WIDTH: ping_storage_data_268 <= (fillup_transition == 1'b1) ? i_input_data[571 % IN_WIDTH] : ping_storage_data_268 ^ i_input_data[571 % IN_WIDTH];
                715 / IN_WIDTH: ping_storage_data_268 <= (fillup_transition == 1'b1) ? i_input_data[715 % IN_WIDTH] : ping_storage_data_268 ^ i_input_data[715 % IN_WIDTH];
                1132 / IN_WIDTH: ping_storage_data_268 <= (fillup_transition == 1'b1) ? i_input_data[1132 % IN_WIDTH] : ping_storage_data_268 ^ i_input_data[1132 % IN_WIDTH];
                default: ping_storage_data_268 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_268;
                endcase
            end else begin
                case (input_count)
                340 / IN_WIDTH: pong_storage_data_268 <= (fillup_transition == 1'b1) ? i_input_data[340 % IN_WIDTH] : pong_storage_data_268 ^ i_input_data[340 % IN_WIDTH];
                438 / IN_WIDTH: pong_storage_data_268 <= (fillup_transition == 1'b1) ? i_input_data[438 % IN_WIDTH] : pong_storage_data_268 ^ i_input_data[438 % IN_WIDTH];
                571 / IN_WIDTH: pong_storage_data_268 <= (fillup_transition == 1'b1) ? i_input_data[571 % IN_WIDTH] : pong_storage_data_268 ^ i_input_data[571 % IN_WIDTH];
                715 / IN_WIDTH: pong_storage_data_268 <= (fillup_transition == 1'b1) ? i_input_data[715 % IN_WIDTH] : pong_storage_data_268 ^ i_input_data[715 % IN_WIDTH];
                1132 / IN_WIDTH: pong_storage_data_268 <= (fillup_transition == 1'b1) ? i_input_data[1132 % IN_WIDTH] : pong_storage_data_268 ^ i_input_data[1132 % IN_WIDTH];
                default: pong_storage_data_268 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_268;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_268 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_268;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_268 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_268;
            end
        end
    end
end

logic ping_storage_data_269;
logic pong_storage_data_269;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_269 <= 1'b0;
        pong_storage_data_269 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                341 / IN_WIDTH: ping_storage_data_269 <= (fillup_transition == 1'b1) ? i_input_data[341 % IN_WIDTH] : ping_storage_data_269 ^ i_input_data[341 % IN_WIDTH];
                439 / IN_WIDTH: ping_storage_data_269 <= (fillup_transition == 1'b1) ? i_input_data[439 % IN_WIDTH] : ping_storage_data_269 ^ i_input_data[439 % IN_WIDTH];
                572 / IN_WIDTH: ping_storage_data_269 <= (fillup_transition == 1'b1) ? i_input_data[572 % IN_WIDTH] : ping_storage_data_269 ^ i_input_data[572 % IN_WIDTH];
                716 / IN_WIDTH: ping_storage_data_269 <= (fillup_transition == 1'b1) ? i_input_data[716 % IN_WIDTH] : ping_storage_data_269 ^ i_input_data[716 % IN_WIDTH];
                1133 / IN_WIDTH: ping_storage_data_269 <= (fillup_transition == 1'b1) ? i_input_data[1133 % IN_WIDTH] : ping_storage_data_269 ^ i_input_data[1133 % IN_WIDTH];
                default: ping_storage_data_269 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_269;
                endcase
            end else begin
                case (input_count)
                341 / IN_WIDTH: pong_storage_data_269 <= (fillup_transition == 1'b1) ? i_input_data[341 % IN_WIDTH] : pong_storage_data_269 ^ i_input_data[341 % IN_WIDTH];
                439 / IN_WIDTH: pong_storage_data_269 <= (fillup_transition == 1'b1) ? i_input_data[439 % IN_WIDTH] : pong_storage_data_269 ^ i_input_data[439 % IN_WIDTH];
                572 / IN_WIDTH: pong_storage_data_269 <= (fillup_transition == 1'b1) ? i_input_data[572 % IN_WIDTH] : pong_storage_data_269 ^ i_input_data[572 % IN_WIDTH];
                716 / IN_WIDTH: pong_storage_data_269 <= (fillup_transition == 1'b1) ? i_input_data[716 % IN_WIDTH] : pong_storage_data_269 ^ i_input_data[716 % IN_WIDTH];
                1133 / IN_WIDTH: pong_storage_data_269 <= (fillup_transition == 1'b1) ? i_input_data[1133 % IN_WIDTH] : pong_storage_data_269 ^ i_input_data[1133 % IN_WIDTH];
                default: pong_storage_data_269 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_269;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_269 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_269;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_269 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_269;
            end
        end
    end
end

logic ping_storage_data_270;
logic pong_storage_data_270;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_270 <= 1'b0;
        pong_storage_data_270 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                342 / IN_WIDTH: ping_storage_data_270 <= (fillup_transition == 1'b1) ? i_input_data[342 % IN_WIDTH] : ping_storage_data_270 ^ i_input_data[342 % IN_WIDTH];
                440 / IN_WIDTH: ping_storage_data_270 <= (fillup_transition == 1'b1) ? i_input_data[440 % IN_WIDTH] : ping_storage_data_270 ^ i_input_data[440 % IN_WIDTH];
                573 / IN_WIDTH: ping_storage_data_270 <= (fillup_transition == 1'b1) ? i_input_data[573 % IN_WIDTH] : ping_storage_data_270 ^ i_input_data[573 % IN_WIDTH];
                717 / IN_WIDTH: ping_storage_data_270 <= (fillup_transition == 1'b1) ? i_input_data[717 % IN_WIDTH] : ping_storage_data_270 ^ i_input_data[717 % IN_WIDTH];
                1134 / IN_WIDTH: ping_storage_data_270 <= (fillup_transition == 1'b1) ? i_input_data[1134 % IN_WIDTH] : ping_storage_data_270 ^ i_input_data[1134 % IN_WIDTH];
                default: ping_storage_data_270 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_270;
                endcase
            end else begin
                case (input_count)
                342 / IN_WIDTH: pong_storage_data_270 <= (fillup_transition == 1'b1) ? i_input_data[342 % IN_WIDTH] : pong_storage_data_270 ^ i_input_data[342 % IN_WIDTH];
                440 / IN_WIDTH: pong_storage_data_270 <= (fillup_transition == 1'b1) ? i_input_data[440 % IN_WIDTH] : pong_storage_data_270 ^ i_input_data[440 % IN_WIDTH];
                573 / IN_WIDTH: pong_storage_data_270 <= (fillup_transition == 1'b1) ? i_input_data[573 % IN_WIDTH] : pong_storage_data_270 ^ i_input_data[573 % IN_WIDTH];
                717 / IN_WIDTH: pong_storage_data_270 <= (fillup_transition == 1'b1) ? i_input_data[717 % IN_WIDTH] : pong_storage_data_270 ^ i_input_data[717 % IN_WIDTH];
                1134 / IN_WIDTH: pong_storage_data_270 <= (fillup_transition == 1'b1) ? i_input_data[1134 % IN_WIDTH] : pong_storage_data_270 ^ i_input_data[1134 % IN_WIDTH];
                default: pong_storage_data_270 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_270;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_270 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_270;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_270 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_270;
            end
        end
    end
end

logic ping_storage_data_271;
logic pong_storage_data_271;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_271 <= 1'b0;
        pong_storage_data_271 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                343 / IN_WIDTH: ping_storage_data_271 <= (fillup_transition == 1'b1) ? i_input_data[343 % IN_WIDTH] : ping_storage_data_271 ^ i_input_data[343 % IN_WIDTH];
                441 / IN_WIDTH: ping_storage_data_271 <= (fillup_transition == 1'b1) ? i_input_data[441 % IN_WIDTH] : ping_storage_data_271 ^ i_input_data[441 % IN_WIDTH];
                574 / IN_WIDTH: ping_storage_data_271 <= (fillup_transition == 1'b1) ? i_input_data[574 % IN_WIDTH] : ping_storage_data_271 ^ i_input_data[574 % IN_WIDTH];
                718 / IN_WIDTH: ping_storage_data_271 <= (fillup_transition == 1'b1) ? i_input_data[718 % IN_WIDTH] : ping_storage_data_271 ^ i_input_data[718 % IN_WIDTH];
                1135 / IN_WIDTH: ping_storage_data_271 <= (fillup_transition == 1'b1) ? i_input_data[1135 % IN_WIDTH] : ping_storage_data_271 ^ i_input_data[1135 % IN_WIDTH];
                default: ping_storage_data_271 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_271;
                endcase
            end else begin
                case (input_count)
                343 / IN_WIDTH: pong_storage_data_271 <= (fillup_transition == 1'b1) ? i_input_data[343 % IN_WIDTH] : pong_storage_data_271 ^ i_input_data[343 % IN_WIDTH];
                441 / IN_WIDTH: pong_storage_data_271 <= (fillup_transition == 1'b1) ? i_input_data[441 % IN_WIDTH] : pong_storage_data_271 ^ i_input_data[441 % IN_WIDTH];
                574 / IN_WIDTH: pong_storage_data_271 <= (fillup_transition == 1'b1) ? i_input_data[574 % IN_WIDTH] : pong_storage_data_271 ^ i_input_data[574 % IN_WIDTH];
                718 / IN_WIDTH: pong_storage_data_271 <= (fillup_transition == 1'b1) ? i_input_data[718 % IN_WIDTH] : pong_storage_data_271 ^ i_input_data[718 % IN_WIDTH];
                1135 / IN_WIDTH: pong_storage_data_271 <= (fillup_transition == 1'b1) ? i_input_data[1135 % IN_WIDTH] : pong_storage_data_271 ^ i_input_data[1135 % IN_WIDTH];
                default: pong_storage_data_271 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_271;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_271 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_271;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_271 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_271;
            end
        end
    end
end

logic ping_storage_data_272;
logic pong_storage_data_272;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_272 <= 1'b0;
        pong_storage_data_272 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                344 / IN_WIDTH: ping_storage_data_272 <= (fillup_transition == 1'b1) ? i_input_data[344 % IN_WIDTH] : ping_storage_data_272 ^ i_input_data[344 % IN_WIDTH];
                442 / IN_WIDTH: ping_storage_data_272 <= (fillup_transition == 1'b1) ? i_input_data[442 % IN_WIDTH] : ping_storage_data_272 ^ i_input_data[442 % IN_WIDTH];
                575 / IN_WIDTH: ping_storage_data_272 <= (fillup_transition == 1'b1) ? i_input_data[575 % IN_WIDTH] : ping_storage_data_272 ^ i_input_data[575 % IN_WIDTH];
                719 / IN_WIDTH: ping_storage_data_272 <= (fillup_transition == 1'b1) ? i_input_data[719 % IN_WIDTH] : ping_storage_data_272 ^ i_input_data[719 % IN_WIDTH];
                1136 / IN_WIDTH: ping_storage_data_272 <= (fillup_transition == 1'b1) ? i_input_data[1136 % IN_WIDTH] : ping_storage_data_272 ^ i_input_data[1136 % IN_WIDTH];
                default: ping_storage_data_272 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_272;
                endcase
            end else begin
                case (input_count)
                344 / IN_WIDTH: pong_storage_data_272 <= (fillup_transition == 1'b1) ? i_input_data[344 % IN_WIDTH] : pong_storage_data_272 ^ i_input_data[344 % IN_WIDTH];
                442 / IN_WIDTH: pong_storage_data_272 <= (fillup_transition == 1'b1) ? i_input_data[442 % IN_WIDTH] : pong_storage_data_272 ^ i_input_data[442 % IN_WIDTH];
                575 / IN_WIDTH: pong_storage_data_272 <= (fillup_transition == 1'b1) ? i_input_data[575 % IN_WIDTH] : pong_storage_data_272 ^ i_input_data[575 % IN_WIDTH];
                719 / IN_WIDTH: pong_storage_data_272 <= (fillup_transition == 1'b1) ? i_input_data[719 % IN_WIDTH] : pong_storage_data_272 ^ i_input_data[719 % IN_WIDTH];
                1136 / IN_WIDTH: pong_storage_data_272 <= (fillup_transition == 1'b1) ? i_input_data[1136 % IN_WIDTH] : pong_storage_data_272 ^ i_input_data[1136 % IN_WIDTH];
                default: pong_storage_data_272 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_272;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_272 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_272;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_272 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_272;
            end
        end
    end
end

logic ping_storage_data_273;
logic pong_storage_data_273;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_273 <= 1'b0;
        pong_storage_data_273 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                345 / IN_WIDTH: ping_storage_data_273 <= (fillup_transition == 1'b1) ? i_input_data[345 % IN_WIDTH] : ping_storage_data_273 ^ i_input_data[345 % IN_WIDTH];
                443 / IN_WIDTH: ping_storage_data_273 <= (fillup_transition == 1'b1) ? i_input_data[443 % IN_WIDTH] : ping_storage_data_273 ^ i_input_data[443 % IN_WIDTH];
                480 / IN_WIDTH: ping_storage_data_273 <= (fillup_transition == 1'b1) ? i_input_data[480 % IN_WIDTH] : ping_storage_data_273 ^ i_input_data[480 % IN_WIDTH];
                720 / IN_WIDTH: ping_storage_data_273 <= (fillup_transition == 1'b1) ? i_input_data[720 % IN_WIDTH] : ping_storage_data_273 ^ i_input_data[720 % IN_WIDTH];
                1137 / IN_WIDTH: ping_storage_data_273 <= (fillup_transition == 1'b1) ? i_input_data[1137 % IN_WIDTH] : ping_storage_data_273 ^ i_input_data[1137 % IN_WIDTH];
                default: ping_storage_data_273 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_273;
                endcase
            end else begin
                case (input_count)
                345 / IN_WIDTH: pong_storage_data_273 <= (fillup_transition == 1'b1) ? i_input_data[345 % IN_WIDTH] : pong_storage_data_273 ^ i_input_data[345 % IN_WIDTH];
                443 / IN_WIDTH: pong_storage_data_273 <= (fillup_transition == 1'b1) ? i_input_data[443 % IN_WIDTH] : pong_storage_data_273 ^ i_input_data[443 % IN_WIDTH];
                480 / IN_WIDTH: pong_storage_data_273 <= (fillup_transition == 1'b1) ? i_input_data[480 % IN_WIDTH] : pong_storage_data_273 ^ i_input_data[480 % IN_WIDTH];
                720 / IN_WIDTH: pong_storage_data_273 <= (fillup_transition == 1'b1) ? i_input_data[720 % IN_WIDTH] : pong_storage_data_273 ^ i_input_data[720 % IN_WIDTH];
                1137 / IN_WIDTH: pong_storage_data_273 <= (fillup_transition == 1'b1) ? i_input_data[1137 % IN_WIDTH] : pong_storage_data_273 ^ i_input_data[1137 % IN_WIDTH];
                default: pong_storage_data_273 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_273;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_273 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_273;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_273 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_273;
            end
        end
    end
end

logic ping_storage_data_274;
logic pong_storage_data_274;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_274 <= 1'b0;
        pong_storage_data_274 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                346 / IN_WIDTH: ping_storage_data_274 <= (fillup_transition == 1'b1) ? i_input_data[346 % IN_WIDTH] : ping_storage_data_274 ^ i_input_data[346 % IN_WIDTH];
                444 / IN_WIDTH: ping_storage_data_274 <= (fillup_transition == 1'b1) ? i_input_data[444 % IN_WIDTH] : ping_storage_data_274 ^ i_input_data[444 % IN_WIDTH];
                481 / IN_WIDTH: ping_storage_data_274 <= (fillup_transition == 1'b1) ? i_input_data[481 % IN_WIDTH] : ping_storage_data_274 ^ i_input_data[481 % IN_WIDTH];
                721 / IN_WIDTH: ping_storage_data_274 <= (fillup_transition == 1'b1) ? i_input_data[721 % IN_WIDTH] : ping_storage_data_274 ^ i_input_data[721 % IN_WIDTH];
                1138 / IN_WIDTH: ping_storage_data_274 <= (fillup_transition == 1'b1) ? i_input_data[1138 % IN_WIDTH] : ping_storage_data_274 ^ i_input_data[1138 % IN_WIDTH];
                default: ping_storage_data_274 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_274;
                endcase
            end else begin
                case (input_count)
                346 / IN_WIDTH: pong_storage_data_274 <= (fillup_transition == 1'b1) ? i_input_data[346 % IN_WIDTH] : pong_storage_data_274 ^ i_input_data[346 % IN_WIDTH];
                444 / IN_WIDTH: pong_storage_data_274 <= (fillup_transition == 1'b1) ? i_input_data[444 % IN_WIDTH] : pong_storage_data_274 ^ i_input_data[444 % IN_WIDTH];
                481 / IN_WIDTH: pong_storage_data_274 <= (fillup_transition == 1'b1) ? i_input_data[481 % IN_WIDTH] : pong_storage_data_274 ^ i_input_data[481 % IN_WIDTH];
                721 / IN_WIDTH: pong_storage_data_274 <= (fillup_transition == 1'b1) ? i_input_data[721 % IN_WIDTH] : pong_storage_data_274 ^ i_input_data[721 % IN_WIDTH];
                1138 / IN_WIDTH: pong_storage_data_274 <= (fillup_transition == 1'b1) ? i_input_data[1138 % IN_WIDTH] : pong_storage_data_274 ^ i_input_data[1138 % IN_WIDTH];
                default: pong_storage_data_274 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_274;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_274 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_274;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_274 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_274;
            end
        end
    end
end

logic ping_storage_data_275;
logic pong_storage_data_275;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_275 <= 1'b0;
        pong_storage_data_275 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                347 / IN_WIDTH: ping_storage_data_275 <= (fillup_transition == 1'b1) ? i_input_data[347 % IN_WIDTH] : ping_storage_data_275 ^ i_input_data[347 % IN_WIDTH];
                445 / IN_WIDTH: ping_storage_data_275 <= (fillup_transition == 1'b1) ? i_input_data[445 % IN_WIDTH] : ping_storage_data_275 ^ i_input_data[445 % IN_WIDTH];
                482 / IN_WIDTH: ping_storage_data_275 <= (fillup_transition == 1'b1) ? i_input_data[482 % IN_WIDTH] : ping_storage_data_275 ^ i_input_data[482 % IN_WIDTH];
                722 / IN_WIDTH: ping_storage_data_275 <= (fillup_transition == 1'b1) ? i_input_data[722 % IN_WIDTH] : ping_storage_data_275 ^ i_input_data[722 % IN_WIDTH];
                1139 / IN_WIDTH: ping_storage_data_275 <= (fillup_transition == 1'b1) ? i_input_data[1139 % IN_WIDTH] : ping_storage_data_275 ^ i_input_data[1139 % IN_WIDTH];
                default: ping_storage_data_275 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_275;
                endcase
            end else begin
                case (input_count)
                347 / IN_WIDTH: pong_storage_data_275 <= (fillup_transition == 1'b1) ? i_input_data[347 % IN_WIDTH] : pong_storage_data_275 ^ i_input_data[347 % IN_WIDTH];
                445 / IN_WIDTH: pong_storage_data_275 <= (fillup_transition == 1'b1) ? i_input_data[445 % IN_WIDTH] : pong_storage_data_275 ^ i_input_data[445 % IN_WIDTH];
                482 / IN_WIDTH: pong_storage_data_275 <= (fillup_transition == 1'b1) ? i_input_data[482 % IN_WIDTH] : pong_storage_data_275 ^ i_input_data[482 % IN_WIDTH];
                722 / IN_WIDTH: pong_storage_data_275 <= (fillup_transition == 1'b1) ? i_input_data[722 % IN_WIDTH] : pong_storage_data_275 ^ i_input_data[722 % IN_WIDTH];
                1139 / IN_WIDTH: pong_storage_data_275 <= (fillup_transition == 1'b1) ? i_input_data[1139 % IN_WIDTH] : pong_storage_data_275 ^ i_input_data[1139 % IN_WIDTH];
                default: pong_storage_data_275 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_275;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_275 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_275;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_275 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_275;
            end
        end
    end
end

logic ping_storage_data_276;
logic pong_storage_data_276;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_276 <= 1'b0;
        pong_storage_data_276 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                348 / IN_WIDTH: ping_storage_data_276 <= (fillup_transition == 1'b1) ? i_input_data[348 % IN_WIDTH] : ping_storage_data_276 ^ i_input_data[348 % IN_WIDTH];
                446 / IN_WIDTH: ping_storage_data_276 <= (fillup_transition == 1'b1) ? i_input_data[446 % IN_WIDTH] : ping_storage_data_276 ^ i_input_data[446 % IN_WIDTH];
                483 / IN_WIDTH: ping_storage_data_276 <= (fillup_transition == 1'b1) ? i_input_data[483 % IN_WIDTH] : ping_storage_data_276 ^ i_input_data[483 % IN_WIDTH];
                723 / IN_WIDTH: ping_storage_data_276 <= (fillup_transition == 1'b1) ? i_input_data[723 % IN_WIDTH] : ping_storage_data_276 ^ i_input_data[723 % IN_WIDTH];
                1140 / IN_WIDTH: ping_storage_data_276 <= (fillup_transition == 1'b1) ? i_input_data[1140 % IN_WIDTH] : ping_storage_data_276 ^ i_input_data[1140 % IN_WIDTH];
                default: ping_storage_data_276 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_276;
                endcase
            end else begin
                case (input_count)
                348 / IN_WIDTH: pong_storage_data_276 <= (fillup_transition == 1'b1) ? i_input_data[348 % IN_WIDTH] : pong_storage_data_276 ^ i_input_data[348 % IN_WIDTH];
                446 / IN_WIDTH: pong_storage_data_276 <= (fillup_transition == 1'b1) ? i_input_data[446 % IN_WIDTH] : pong_storage_data_276 ^ i_input_data[446 % IN_WIDTH];
                483 / IN_WIDTH: pong_storage_data_276 <= (fillup_transition == 1'b1) ? i_input_data[483 % IN_WIDTH] : pong_storage_data_276 ^ i_input_data[483 % IN_WIDTH];
                723 / IN_WIDTH: pong_storage_data_276 <= (fillup_transition == 1'b1) ? i_input_data[723 % IN_WIDTH] : pong_storage_data_276 ^ i_input_data[723 % IN_WIDTH];
                1140 / IN_WIDTH: pong_storage_data_276 <= (fillup_transition == 1'b1) ? i_input_data[1140 % IN_WIDTH] : pong_storage_data_276 ^ i_input_data[1140 % IN_WIDTH];
                default: pong_storage_data_276 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_276;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_276 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_276;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_276 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_276;
            end
        end
    end
end

logic ping_storage_data_277;
logic pong_storage_data_277;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_277 <= 1'b0;
        pong_storage_data_277 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                349 / IN_WIDTH: ping_storage_data_277 <= (fillup_transition == 1'b1) ? i_input_data[349 % IN_WIDTH] : ping_storage_data_277 ^ i_input_data[349 % IN_WIDTH];
                447 / IN_WIDTH: ping_storage_data_277 <= (fillup_transition == 1'b1) ? i_input_data[447 % IN_WIDTH] : ping_storage_data_277 ^ i_input_data[447 % IN_WIDTH];
                484 / IN_WIDTH: ping_storage_data_277 <= (fillup_transition == 1'b1) ? i_input_data[484 % IN_WIDTH] : ping_storage_data_277 ^ i_input_data[484 % IN_WIDTH];
                724 / IN_WIDTH: ping_storage_data_277 <= (fillup_transition == 1'b1) ? i_input_data[724 % IN_WIDTH] : ping_storage_data_277 ^ i_input_data[724 % IN_WIDTH];
                1141 / IN_WIDTH: ping_storage_data_277 <= (fillup_transition == 1'b1) ? i_input_data[1141 % IN_WIDTH] : ping_storage_data_277 ^ i_input_data[1141 % IN_WIDTH];
                default: ping_storage_data_277 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_277;
                endcase
            end else begin
                case (input_count)
                349 / IN_WIDTH: pong_storage_data_277 <= (fillup_transition == 1'b1) ? i_input_data[349 % IN_WIDTH] : pong_storage_data_277 ^ i_input_data[349 % IN_WIDTH];
                447 / IN_WIDTH: pong_storage_data_277 <= (fillup_transition == 1'b1) ? i_input_data[447 % IN_WIDTH] : pong_storage_data_277 ^ i_input_data[447 % IN_WIDTH];
                484 / IN_WIDTH: pong_storage_data_277 <= (fillup_transition == 1'b1) ? i_input_data[484 % IN_WIDTH] : pong_storage_data_277 ^ i_input_data[484 % IN_WIDTH];
                724 / IN_WIDTH: pong_storage_data_277 <= (fillup_transition == 1'b1) ? i_input_data[724 % IN_WIDTH] : pong_storage_data_277 ^ i_input_data[724 % IN_WIDTH];
                1141 / IN_WIDTH: pong_storage_data_277 <= (fillup_transition == 1'b1) ? i_input_data[1141 % IN_WIDTH] : pong_storage_data_277 ^ i_input_data[1141 % IN_WIDTH];
                default: pong_storage_data_277 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_277;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_277 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_277;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_277 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_277;
            end
        end
    end
end

logic ping_storage_data_278;
logic pong_storage_data_278;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_278 <= 1'b0;
        pong_storage_data_278 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                350 / IN_WIDTH: ping_storage_data_278 <= (fillup_transition == 1'b1) ? i_input_data[350 % IN_WIDTH] : ping_storage_data_278 ^ i_input_data[350 % IN_WIDTH];
                448 / IN_WIDTH: ping_storage_data_278 <= (fillup_transition == 1'b1) ? i_input_data[448 % IN_WIDTH] : ping_storage_data_278 ^ i_input_data[448 % IN_WIDTH];
                485 / IN_WIDTH: ping_storage_data_278 <= (fillup_transition == 1'b1) ? i_input_data[485 % IN_WIDTH] : ping_storage_data_278 ^ i_input_data[485 % IN_WIDTH];
                725 / IN_WIDTH: ping_storage_data_278 <= (fillup_transition == 1'b1) ? i_input_data[725 % IN_WIDTH] : ping_storage_data_278 ^ i_input_data[725 % IN_WIDTH];
                1142 / IN_WIDTH: ping_storage_data_278 <= (fillup_transition == 1'b1) ? i_input_data[1142 % IN_WIDTH] : ping_storage_data_278 ^ i_input_data[1142 % IN_WIDTH];
                default: ping_storage_data_278 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_278;
                endcase
            end else begin
                case (input_count)
                350 / IN_WIDTH: pong_storage_data_278 <= (fillup_transition == 1'b1) ? i_input_data[350 % IN_WIDTH] : pong_storage_data_278 ^ i_input_data[350 % IN_WIDTH];
                448 / IN_WIDTH: pong_storage_data_278 <= (fillup_transition == 1'b1) ? i_input_data[448 % IN_WIDTH] : pong_storage_data_278 ^ i_input_data[448 % IN_WIDTH];
                485 / IN_WIDTH: pong_storage_data_278 <= (fillup_transition == 1'b1) ? i_input_data[485 % IN_WIDTH] : pong_storage_data_278 ^ i_input_data[485 % IN_WIDTH];
                725 / IN_WIDTH: pong_storage_data_278 <= (fillup_transition == 1'b1) ? i_input_data[725 % IN_WIDTH] : pong_storage_data_278 ^ i_input_data[725 % IN_WIDTH];
                1142 / IN_WIDTH: pong_storage_data_278 <= (fillup_transition == 1'b1) ? i_input_data[1142 % IN_WIDTH] : pong_storage_data_278 ^ i_input_data[1142 % IN_WIDTH];
                default: pong_storage_data_278 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_278;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_278 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_278;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_278 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_278;
            end
        end
    end
end

logic ping_storage_data_279;
logic pong_storage_data_279;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_279 <= 1'b0;
        pong_storage_data_279 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                351 / IN_WIDTH: ping_storage_data_279 <= (fillup_transition == 1'b1) ? i_input_data[351 % IN_WIDTH] : ping_storage_data_279 ^ i_input_data[351 % IN_WIDTH];
                449 / IN_WIDTH: ping_storage_data_279 <= (fillup_transition == 1'b1) ? i_input_data[449 % IN_WIDTH] : ping_storage_data_279 ^ i_input_data[449 % IN_WIDTH];
                486 / IN_WIDTH: ping_storage_data_279 <= (fillup_transition == 1'b1) ? i_input_data[486 % IN_WIDTH] : ping_storage_data_279 ^ i_input_data[486 % IN_WIDTH];
                726 / IN_WIDTH: ping_storage_data_279 <= (fillup_transition == 1'b1) ? i_input_data[726 % IN_WIDTH] : ping_storage_data_279 ^ i_input_data[726 % IN_WIDTH];
                1143 / IN_WIDTH: ping_storage_data_279 <= (fillup_transition == 1'b1) ? i_input_data[1143 % IN_WIDTH] : ping_storage_data_279 ^ i_input_data[1143 % IN_WIDTH];
                default: ping_storage_data_279 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_279;
                endcase
            end else begin
                case (input_count)
                351 / IN_WIDTH: pong_storage_data_279 <= (fillup_transition == 1'b1) ? i_input_data[351 % IN_WIDTH] : pong_storage_data_279 ^ i_input_data[351 % IN_WIDTH];
                449 / IN_WIDTH: pong_storage_data_279 <= (fillup_transition == 1'b1) ? i_input_data[449 % IN_WIDTH] : pong_storage_data_279 ^ i_input_data[449 % IN_WIDTH];
                486 / IN_WIDTH: pong_storage_data_279 <= (fillup_transition == 1'b1) ? i_input_data[486 % IN_WIDTH] : pong_storage_data_279 ^ i_input_data[486 % IN_WIDTH];
                726 / IN_WIDTH: pong_storage_data_279 <= (fillup_transition == 1'b1) ? i_input_data[726 % IN_WIDTH] : pong_storage_data_279 ^ i_input_data[726 % IN_WIDTH];
                1143 / IN_WIDTH: pong_storage_data_279 <= (fillup_transition == 1'b1) ? i_input_data[1143 % IN_WIDTH] : pong_storage_data_279 ^ i_input_data[1143 % IN_WIDTH];
                default: pong_storage_data_279 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_279;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_279 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_279;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_279 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_279;
            end
        end
    end
end

logic ping_storage_data_280;
logic pong_storage_data_280;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_280 <= 1'b0;
        pong_storage_data_280 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                352 / IN_WIDTH: ping_storage_data_280 <= (fillup_transition == 1'b1) ? i_input_data[352 % IN_WIDTH] : ping_storage_data_280 ^ i_input_data[352 % IN_WIDTH];
                450 / IN_WIDTH: ping_storage_data_280 <= (fillup_transition == 1'b1) ? i_input_data[450 % IN_WIDTH] : ping_storage_data_280 ^ i_input_data[450 % IN_WIDTH];
                487 / IN_WIDTH: ping_storage_data_280 <= (fillup_transition == 1'b1) ? i_input_data[487 % IN_WIDTH] : ping_storage_data_280 ^ i_input_data[487 % IN_WIDTH];
                727 / IN_WIDTH: ping_storage_data_280 <= (fillup_transition == 1'b1) ? i_input_data[727 % IN_WIDTH] : ping_storage_data_280 ^ i_input_data[727 % IN_WIDTH];
                1144 / IN_WIDTH: ping_storage_data_280 <= (fillup_transition == 1'b1) ? i_input_data[1144 % IN_WIDTH] : ping_storage_data_280 ^ i_input_data[1144 % IN_WIDTH];
                default: ping_storage_data_280 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_280;
                endcase
            end else begin
                case (input_count)
                352 / IN_WIDTH: pong_storage_data_280 <= (fillup_transition == 1'b1) ? i_input_data[352 % IN_WIDTH] : pong_storage_data_280 ^ i_input_data[352 % IN_WIDTH];
                450 / IN_WIDTH: pong_storage_data_280 <= (fillup_transition == 1'b1) ? i_input_data[450 % IN_WIDTH] : pong_storage_data_280 ^ i_input_data[450 % IN_WIDTH];
                487 / IN_WIDTH: pong_storage_data_280 <= (fillup_transition == 1'b1) ? i_input_data[487 % IN_WIDTH] : pong_storage_data_280 ^ i_input_data[487 % IN_WIDTH];
                727 / IN_WIDTH: pong_storage_data_280 <= (fillup_transition == 1'b1) ? i_input_data[727 % IN_WIDTH] : pong_storage_data_280 ^ i_input_data[727 % IN_WIDTH];
                1144 / IN_WIDTH: pong_storage_data_280 <= (fillup_transition == 1'b1) ? i_input_data[1144 % IN_WIDTH] : pong_storage_data_280 ^ i_input_data[1144 % IN_WIDTH];
                default: pong_storage_data_280 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_280;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_280 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_280;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_280 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_280;
            end
        end
    end
end

logic ping_storage_data_281;
logic pong_storage_data_281;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_281 <= 1'b0;
        pong_storage_data_281 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                353 / IN_WIDTH: ping_storage_data_281 <= (fillup_transition == 1'b1) ? i_input_data[353 % IN_WIDTH] : ping_storage_data_281 ^ i_input_data[353 % IN_WIDTH];
                451 / IN_WIDTH: ping_storage_data_281 <= (fillup_transition == 1'b1) ? i_input_data[451 % IN_WIDTH] : ping_storage_data_281 ^ i_input_data[451 % IN_WIDTH];
                488 / IN_WIDTH: ping_storage_data_281 <= (fillup_transition == 1'b1) ? i_input_data[488 % IN_WIDTH] : ping_storage_data_281 ^ i_input_data[488 % IN_WIDTH];
                728 / IN_WIDTH: ping_storage_data_281 <= (fillup_transition == 1'b1) ? i_input_data[728 % IN_WIDTH] : ping_storage_data_281 ^ i_input_data[728 % IN_WIDTH];
                1145 / IN_WIDTH: ping_storage_data_281 <= (fillup_transition == 1'b1) ? i_input_data[1145 % IN_WIDTH] : ping_storage_data_281 ^ i_input_data[1145 % IN_WIDTH];
                default: ping_storage_data_281 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_281;
                endcase
            end else begin
                case (input_count)
                353 / IN_WIDTH: pong_storage_data_281 <= (fillup_transition == 1'b1) ? i_input_data[353 % IN_WIDTH] : pong_storage_data_281 ^ i_input_data[353 % IN_WIDTH];
                451 / IN_WIDTH: pong_storage_data_281 <= (fillup_transition == 1'b1) ? i_input_data[451 % IN_WIDTH] : pong_storage_data_281 ^ i_input_data[451 % IN_WIDTH];
                488 / IN_WIDTH: pong_storage_data_281 <= (fillup_transition == 1'b1) ? i_input_data[488 % IN_WIDTH] : pong_storage_data_281 ^ i_input_data[488 % IN_WIDTH];
                728 / IN_WIDTH: pong_storage_data_281 <= (fillup_transition == 1'b1) ? i_input_data[728 % IN_WIDTH] : pong_storage_data_281 ^ i_input_data[728 % IN_WIDTH];
                1145 / IN_WIDTH: pong_storage_data_281 <= (fillup_transition == 1'b1) ? i_input_data[1145 % IN_WIDTH] : pong_storage_data_281 ^ i_input_data[1145 % IN_WIDTH];
                default: pong_storage_data_281 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_281;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_281 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_281;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_281 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_281;
            end
        end
    end
end

logic ping_storage_data_282;
logic pong_storage_data_282;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_282 <= 1'b0;
        pong_storage_data_282 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                354 / IN_WIDTH: ping_storage_data_282 <= (fillup_transition == 1'b1) ? i_input_data[354 % IN_WIDTH] : ping_storage_data_282 ^ i_input_data[354 % IN_WIDTH];
                452 / IN_WIDTH: ping_storage_data_282 <= (fillup_transition == 1'b1) ? i_input_data[452 % IN_WIDTH] : ping_storage_data_282 ^ i_input_data[452 % IN_WIDTH];
                489 / IN_WIDTH: ping_storage_data_282 <= (fillup_transition == 1'b1) ? i_input_data[489 % IN_WIDTH] : ping_storage_data_282 ^ i_input_data[489 % IN_WIDTH];
                729 / IN_WIDTH: ping_storage_data_282 <= (fillup_transition == 1'b1) ? i_input_data[729 % IN_WIDTH] : ping_storage_data_282 ^ i_input_data[729 % IN_WIDTH];
                1146 / IN_WIDTH: ping_storage_data_282 <= (fillup_transition == 1'b1) ? i_input_data[1146 % IN_WIDTH] : ping_storage_data_282 ^ i_input_data[1146 % IN_WIDTH];
                default: ping_storage_data_282 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_282;
                endcase
            end else begin
                case (input_count)
                354 / IN_WIDTH: pong_storage_data_282 <= (fillup_transition == 1'b1) ? i_input_data[354 % IN_WIDTH] : pong_storage_data_282 ^ i_input_data[354 % IN_WIDTH];
                452 / IN_WIDTH: pong_storage_data_282 <= (fillup_transition == 1'b1) ? i_input_data[452 % IN_WIDTH] : pong_storage_data_282 ^ i_input_data[452 % IN_WIDTH];
                489 / IN_WIDTH: pong_storage_data_282 <= (fillup_transition == 1'b1) ? i_input_data[489 % IN_WIDTH] : pong_storage_data_282 ^ i_input_data[489 % IN_WIDTH];
                729 / IN_WIDTH: pong_storage_data_282 <= (fillup_transition == 1'b1) ? i_input_data[729 % IN_WIDTH] : pong_storage_data_282 ^ i_input_data[729 % IN_WIDTH];
                1146 / IN_WIDTH: pong_storage_data_282 <= (fillup_transition == 1'b1) ? i_input_data[1146 % IN_WIDTH] : pong_storage_data_282 ^ i_input_data[1146 % IN_WIDTH];
                default: pong_storage_data_282 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_282;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_282 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_282;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_282 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_282;
            end
        end
    end
end

logic ping_storage_data_283;
logic pong_storage_data_283;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_283 <= 1'b0;
        pong_storage_data_283 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                355 / IN_WIDTH: ping_storage_data_283 <= (fillup_transition == 1'b1) ? i_input_data[355 % IN_WIDTH] : ping_storage_data_283 ^ i_input_data[355 % IN_WIDTH];
                453 / IN_WIDTH: ping_storage_data_283 <= (fillup_transition == 1'b1) ? i_input_data[453 % IN_WIDTH] : ping_storage_data_283 ^ i_input_data[453 % IN_WIDTH];
                490 / IN_WIDTH: ping_storage_data_283 <= (fillup_transition == 1'b1) ? i_input_data[490 % IN_WIDTH] : ping_storage_data_283 ^ i_input_data[490 % IN_WIDTH];
                730 / IN_WIDTH: ping_storage_data_283 <= (fillup_transition == 1'b1) ? i_input_data[730 % IN_WIDTH] : ping_storage_data_283 ^ i_input_data[730 % IN_WIDTH];
                1147 / IN_WIDTH: ping_storage_data_283 <= (fillup_transition == 1'b1) ? i_input_data[1147 % IN_WIDTH] : ping_storage_data_283 ^ i_input_data[1147 % IN_WIDTH];
                default: ping_storage_data_283 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_283;
                endcase
            end else begin
                case (input_count)
                355 / IN_WIDTH: pong_storage_data_283 <= (fillup_transition == 1'b1) ? i_input_data[355 % IN_WIDTH] : pong_storage_data_283 ^ i_input_data[355 % IN_WIDTH];
                453 / IN_WIDTH: pong_storage_data_283 <= (fillup_transition == 1'b1) ? i_input_data[453 % IN_WIDTH] : pong_storage_data_283 ^ i_input_data[453 % IN_WIDTH];
                490 / IN_WIDTH: pong_storage_data_283 <= (fillup_transition == 1'b1) ? i_input_data[490 % IN_WIDTH] : pong_storage_data_283 ^ i_input_data[490 % IN_WIDTH];
                730 / IN_WIDTH: pong_storage_data_283 <= (fillup_transition == 1'b1) ? i_input_data[730 % IN_WIDTH] : pong_storage_data_283 ^ i_input_data[730 % IN_WIDTH];
                1147 / IN_WIDTH: pong_storage_data_283 <= (fillup_transition == 1'b1) ? i_input_data[1147 % IN_WIDTH] : pong_storage_data_283 ^ i_input_data[1147 % IN_WIDTH];
                default: pong_storage_data_283 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_283;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_283 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_283;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_283 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_283;
            end
        end
    end
end

logic ping_storage_data_284;
logic pong_storage_data_284;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_284 <= 1'b0;
        pong_storage_data_284 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                356 / IN_WIDTH: ping_storage_data_284 <= (fillup_transition == 1'b1) ? i_input_data[356 % IN_WIDTH] : ping_storage_data_284 ^ i_input_data[356 % IN_WIDTH];
                454 / IN_WIDTH: ping_storage_data_284 <= (fillup_transition == 1'b1) ? i_input_data[454 % IN_WIDTH] : ping_storage_data_284 ^ i_input_data[454 % IN_WIDTH];
                491 / IN_WIDTH: ping_storage_data_284 <= (fillup_transition == 1'b1) ? i_input_data[491 % IN_WIDTH] : ping_storage_data_284 ^ i_input_data[491 % IN_WIDTH];
                731 / IN_WIDTH: ping_storage_data_284 <= (fillup_transition == 1'b1) ? i_input_data[731 % IN_WIDTH] : ping_storage_data_284 ^ i_input_data[731 % IN_WIDTH];
                1148 / IN_WIDTH: ping_storage_data_284 <= (fillup_transition == 1'b1) ? i_input_data[1148 % IN_WIDTH] : ping_storage_data_284 ^ i_input_data[1148 % IN_WIDTH];
                default: ping_storage_data_284 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_284;
                endcase
            end else begin
                case (input_count)
                356 / IN_WIDTH: pong_storage_data_284 <= (fillup_transition == 1'b1) ? i_input_data[356 % IN_WIDTH] : pong_storage_data_284 ^ i_input_data[356 % IN_WIDTH];
                454 / IN_WIDTH: pong_storage_data_284 <= (fillup_transition == 1'b1) ? i_input_data[454 % IN_WIDTH] : pong_storage_data_284 ^ i_input_data[454 % IN_WIDTH];
                491 / IN_WIDTH: pong_storage_data_284 <= (fillup_transition == 1'b1) ? i_input_data[491 % IN_WIDTH] : pong_storage_data_284 ^ i_input_data[491 % IN_WIDTH];
                731 / IN_WIDTH: pong_storage_data_284 <= (fillup_transition == 1'b1) ? i_input_data[731 % IN_WIDTH] : pong_storage_data_284 ^ i_input_data[731 % IN_WIDTH];
                1148 / IN_WIDTH: pong_storage_data_284 <= (fillup_transition == 1'b1) ? i_input_data[1148 % IN_WIDTH] : pong_storage_data_284 ^ i_input_data[1148 % IN_WIDTH];
                default: pong_storage_data_284 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_284;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_284 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_284;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_284 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_284;
            end
        end
    end
end

logic ping_storage_data_285;
logic pong_storage_data_285;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_285 <= 1'b0;
        pong_storage_data_285 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                357 / IN_WIDTH: ping_storage_data_285 <= (fillup_transition == 1'b1) ? i_input_data[357 % IN_WIDTH] : ping_storage_data_285 ^ i_input_data[357 % IN_WIDTH];
                455 / IN_WIDTH: ping_storage_data_285 <= (fillup_transition == 1'b1) ? i_input_data[455 % IN_WIDTH] : ping_storage_data_285 ^ i_input_data[455 % IN_WIDTH];
                492 / IN_WIDTH: ping_storage_data_285 <= (fillup_transition == 1'b1) ? i_input_data[492 % IN_WIDTH] : ping_storage_data_285 ^ i_input_data[492 % IN_WIDTH];
                732 / IN_WIDTH: ping_storage_data_285 <= (fillup_transition == 1'b1) ? i_input_data[732 % IN_WIDTH] : ping_storage_data_285 ^ i_input_data[732 % IN_WIDTH];
                1149 / IN_WIDTH: ping_storage_data_285 <= (fillup_transition == 1'b1) ? i_input_data[1149 % IN_WIDTH] : ping_storage_data_285 ^ i_input_data[1149 % IN_WIDTH];
                default: ping_storage_data_285 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_285;
                endcase
            end else begin
                case (input_count)
                357 / IN_WIDTH: pong_storage_data_285 <= (fillup_transition == 1'b1) ? i_input_data[357 % IN_WIDTH] : pong_storage_data_285 ^ i_input_data[357 % IN_WIDTH];
                455 / IN_WIDTH: pong_storage_data_285 <= (fillup_transition == 1'b1) ? i_input_data[455 % IN_WIDTH] : pong_storage_data_285 ^ i_input_data[455 % IN_WIDTH];
                492 / IN_WIDTH: pong_storage_data_285 <= (fillup_transition == 1'b1) ? i_input_data[492 % IN_WIDTH] : pong_storage_data_285 ^ i_input_data[492 % IN_WIDTH];
                732 / IN_WIDTH: pong_storage_data_285 <= (fillup_transition == 1'b1) ? i_input_data[732 % IN_WIDTH] : pong_storage_data_285 ^ i_input_data[732 % IN_WIDTH];
                1149 / IN_WIDTH: pong_storage_data_285 <= (fillup_transition == 1'b1) ? i_input_data[1149 % IN_WIDTH] : pong_storage_data_285 ^ i_input_data[1149 % IN_WIDTH];
                default: pong_storage_data_285 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_285;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_285 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_285;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_285 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_285;
            end
        end
    end
end

logic ping_storage_data_286;
logic pong_storage_data_286;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_286 <= 1'b0;
        pong_storage_data_286 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                358 / IN_WIDTH: ping_storage_data_286 <= (fillup_transition == 1'b1) ? i_input_data[358 % IN_WIDTH] : ping_storage_data_286 ^ i_input_data[358 % IN_WIDTH];
                456 / IN_WIDTH: ping_storage_data_286 <= (fillup_transition == 1'b1) ? i_input_data[456 % IN_WIDTH] : ping_storage_data_286 ^ i_input_data[456 % IN_WIDTH];
                493 / IN_WIDTH: ping_storage_data_286 <= (fillup_transition == 1'b1) ? i_input_data[493 % IN_WIDTH] : ping_storage_data_286 ^ i_input_data[493 % IN_WIDTH];
                733 / IN_WIDTH: ping_storage_data_286 <= (fillup_transition == 1'b1) ? i_input_data[733 % IN_WIDTH] : ping_storage_data_286 ^ i_input_data[733 % IN_WIDTH];
                1150 / IN_WIDTH: ping_storage_data_286 <= (fillup_transition == 1'b1) ? i_input_data[1150 % IN_WIDTH] : ping_storage_data_286 ^ i_input_data[1150 % IN_WIDTH];
                default: ping_storage_data_286 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_286;
                endcase
            end else begin
                case (input_count)
                358 / IN_WIDTH: pong_storage_data_286 <= (fillup_transition == 1'b1) ? i_input_data[358 % IN_WIDTH] : pong_storage_data_286 ^ i_input_data[358 % IN_WIDTH];
                456 / IN_WIDTH: pong_storage_data_286 <= (fillup_transition == 1'b1) ? i_input_data[456 % IN_WIDTH] : pong_storage_data_286 ^ i_input_data[456 % IN_WIDTH];
                493 / IN_WIDTH: pong_storage_data_286 <= (fillup_transition == 1'b1) ? i_input_data[493 % IN_WIDTH] : pong_storage_data_286 ^ i_input_data[493 % IN_WIDTH];
                733 / IN_WIDTH: pong_storage_data_286 <= (fillup_transition == 1'b1) ? i_input_data[733 % IN_WIDTH] : pong_storage_data_286 ^ i_input_data[733 % IN_WIDTH];
                1150 / IN_WIDTH: pong_storage_data_286 <= (fillup_transition == 1'b1) ? i_input_data[1150 % IN_WIDTH] : pong_storage_data_286 ^ i_input_data[1150 % IN_WIDTH];
                default: pong_storage_data_286 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_286;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_286 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_286;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_286 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_286;
            end
        end
    end
end

logic ping_storage_data_287;
logic pong_storage_data_287;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_287 <= 1'b0;
        pong_storage_data_287 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                359 / IN_WIDTH: ping_storage_data_287 <= (fillup_transition == 1'b1) ? i_input_data[359 % IN_WIDTH] : ping_storage_data_287 ^ i_input_data[359 % IN_WIDTH];
                457 / IN_WIDTH: ping_storage_data_287 <= (fillup_transition == 1'b1) ? i_input_data[457 % IN_WIDTH] : ping_storage_data_287 ^ i_input_data[457 % IN_WIDTH];
                494 / IN_WIDTH: ping_storage_data_287 <= (fillup_transition == 1'b1) ? i_input_data[494 % IN_WIDTH] : ping_storage_data_287 ^ i_input_data[494 % IN_WIDTH];
                734 / IN_WIDTH: ping_storage_data_287 <= (fillup_transition == 1'b1) ? i_input_data[734 % IN_WIDTH] : ping_storage_data_287 ^ i_input_data[734 % IN_WIDTH];
                1151 / IN_WIDTH: ping_storage_data_287 <= (fillup_transition == 1'b1) ? i_input_data[1151 % IN_WIDTH] : ping_storage_data_287 ^ i_input_data[1151 % IN_WIDTH];
                default: ping_storage_data_287 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_287;
                endcase
            end else begin
                case (input_count)
                359 / IN_WIDTH: pong_storage_data_287 <= (fillup_transition == 1'b1) ? i_input_data[359 % IN_WIDTH] : pong_storage_data_287 ^ i_input_data[359 % IN_WIDTH];
                457 / IN_WIDTH: pong_storage_data_287 <= (fillup_transition == 1'b1) ? i_input_data[457 % IN_WIDTH] : pong_storage_data_287 ^ i_input_data[457 % IN_WIDTH];
                494 / IN_WIDTH: pong_storage_data_287 <= (fillup_transition == 1'b1) ? i_input_data[494 % IN_WIDTH] : pong_storage_data_287 ^ i_input_data[494 % IN_WIDTH];
                734 / IN_WIDTH: pong_storage_data_287 <= (fillup_transition == 1'b1) ? i_input_data[734 % IN_WIDTH] : pong_storage_data_287 ^ i_input_data[734 % IN_WIDTH];
                1151 / IN_WIDTH: pong_storage_data_287 <= (fillup_transition == 1'b1) ? i_input_data[1151 % IN_WIDTH] : pong_storage_data_287 ^ i_input_data[1151 % IN_WIDTH];
                default: pong_storage_data_287 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_287;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_287 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_287;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_287 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_287;
            end
        end
    end
end

logic ping_storage_data_288;
logic pong_storage_data_288;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_288 <= 1'b0;
        pong_storage_data_288 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                35 / IN_WIDTH: ping_storage_data_288 <= (fillup_transition == 1'b1) ? i_input_data[35 % IN_WIDTH] : ping_storage_data_288 ^ i_input_data[35 % IN_WIDTH];
                241 / IN_WIDTH: ping_storage_data_288 <= (fillup_transition == 1'b1) ? i_input_data[241 % IN_WIDTH] : ping_storage_data_288 ^ i_input_data[241 % IN_WIDTH];
                799 / IN_WIDTH: ping_storage_data_288 <= (fillup_transition == 1'b1) ? i_input_data[799 % IN_WIDTH] : ping_storage_data_288 ^ i_input_data[799 % IN_WIDTH];
                935 / IN_WIDTH: ping_storage_data_288 <= (fillup_transition == 1'b1) ? i_input_data[935 % IN_WIDTH] : ping_storage_data_288 ^ i_input_data[935 % IN_WIDTH];
                default: ping_storage_data_288 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_288;
                endcase
            end else begin
                case (input_count)
                35 / IN_WIDTH: pong_storage_data_288 <= (fillup_transition == 1'b1) ? i_input_data[35 % IN_WIDTH] : pong_storage_data_288 ^ i_input_data[35 % IN_WIDTH];
                241 / IN_WIDTH: pong_storage_data_288 <= (fillup_transition == 1'b1) ? i_input_data[241 % IN_WIDTH] : pong_storage_data_288 ^ i_input_data[241 % IN_WIDTH];
                799 / IN_WIDTH: pong_storage_data_288 <= (fillup_transition == 1'b1) ? i_input_data[799 % IN_WIDTH] : pong_storage_data_288 ^ i_input_data[799 % IN_WIDTH];
                935 / IN_WIDTH: pong_storage_data_288 <= (fillup_transition == 1'b1) ? i_input_data[935 % IN_WIDTH] : pong_storage_data_288 ^ i_input_data[935 % IN_WIDTH];
                default: pong_storage_data_288 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_288;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_288 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_288;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_288 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_288;
            end
        end
    end
end

logic ping_storage_data_289;
logic pong_storage_data_289;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_289 <= 1'b0;
        pong_storage_data_289 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                36 / IN_WIDTH: ping_storage_data_289 <= (fillup_transition == 1'b1) ? i_input_data[36 % IN_WIDTH] : ping_storage_data_289 ^ i_input_data[36 % IN_WIDTH];
                242 / IN_WIDTH: ping_storage_data_289 <= (fillup_transition == 1'b1) ? i_input_data[242 % IN_WIDTH] : ping_storage_data_289 ^ i_input_data[242 % IN_WIDTH];
                800 / IN_WIDTH: ping_storage_data_289 <= (fillup_transition == 1'b1) ? i_input_data[800 % IN_WIDTH] : ping_storage_data_289 ^ i_input_data[800 % IN_WIDTH];
                936 / IN_WIDTH: ping_storage_data_289 <= (fillup_transition == 1'b1) ? i_input_data[936 % IN_WIDTH] : ping_storage_data_289 ^ i_input_data[936 % IN_WIDTH];
                default: ping_storage_data_289 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_289;
                endcase
            end else begin
                case (input_count)
                36 / IN_WIDTH: pong_storage_data_289 <= (fillup_transition == 1'b1) ? i_input_data[36 % IN_WIDTH] : pong_storage_data_289 ^ i_input_data[36 % IN_WIDTH];
                242 / IN_WIDTH: pong_storage_data_289 <= (fillup_transition == 1'b1) ? i_input_data[242 % IN_WIDTH] : pong_storage_data_289 ^ i_input_data[242 % IN_WIDTH];
                800 / IN_WIDTH: pong_storage_data_289 <= (fillup_transition == 1'b1) ? i_input_data[800 % IN_WIDTH] : pong_storage_data_289 ^ i_input_data[800 % IN_WIDTH];
                936 / IN_WIDTH: pong_storage_data_289 <= (fillup_transition == 1'b1) ? i_input_data[936 % IN_WIDTH] : pong_storage_data_289 ^ i_input_data[936 % IN_WIDTH];
                default: pong_storage_data_289 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_289;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_289 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_289;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_289 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_289;
            end
        end
    end
end

logic ping_storage_data_290;
logic pong_storage_data_290;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_290 <= 1'b0;
        pong_storage_data_290 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                37 / IN_WIDTH: ping_storage_data_290 <= (fillup_transition == 1'b1) ? i_input_data[37 % IN_WIDTH] : ping_storage_data_290 ^ i_input_data[37 % IN_WIDTH];
                243 / IN_WIDTH: ping_storage_data_290 <= (fillup_transition == 1'b1) ? i_input_data[243 % IN_WIDTH] : ping_storage_data_290 ^ i_input_data[243 % IN_WIDTH];
                801 / IN_WIDTH: ping_storage_data_290 <= (fillup_transition == 1'b1) ? i_input_data[801 % IN_WIDTH] : ping_storage_data_290 ^ i_input_data[801 % IN_WIDTH];
                937 / IN_WIDTH: ping_storage_data_290 <= (fillup_transition == 1'b1) ? i_input_data[937 % IN_WIDTH] : ping_storage_data_290 ^ i_input_data[937 % IN_WIDTH];
                default: ping_storage_data_290 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_290;
                endcase
            end else begin
                case (input_count)
                37 / IN_WIDTH: pong_storage_data_290 <= (fillup_transition == 1'b1) ? i_input_data[37 % IN_WIDTH] : pong_storage_data_290 ^ i_input_data[37 % IN_WIDTH];
                243 / IN_WIDTH: pong_storage_data_290 <= (fillup_transition == 1'b1) ? i_input_data[243 % IN_WIDTH] : pong_storage_data_290 ^ i_input_data[243 % IN_WIDTH];
                801 / IN_WIDTH: pong_storage_data_290 <= (fillup_transition == 1'b1) ? i_input_data[801 % IN_WIDTH] : pong_storage_data_290 ^ i_input_data[801 % IN_WIDTH];
                937 / IN_WIDTH: pong_storage_data_290 <= (fillup_transition == 1'b1) ? i_input_data[937 % IN_WIDTH] : pong_storage_data_290 ^ i_input_data[937 % IN_WIDTH];
                default: pong_storage_data_290 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_290;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_290 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_290;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_290 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_290;
            end
        end
    end
end

logic ping_storage_data_291;
logic pong_storage_data_291;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_291 <= 1'b0;
        pong_storage_data_291 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                38 / IN_WIDTH: ping_storage_data_291 <= (fillup_transition == 1'b1) ? i_input_data[38 % IN_WIDTH] : ping_storage_data_291 ^ i_input_data[38 % IN_WIDTH];
                244 / IN_WIDTH: ping_storage_data_291 <= (fillup_transition == 1'b1) ? i_input_data[244 % IN_WIDTH] : ping_storage_data_291 ^ i_input_data[244 % IN_WIDTH];
                802 / IN_WIDTH: ping_storage_data_291 <= (fillup_transition == 1'b1) ? i_input_data[802 % IN_WIDTH] : ping_storage_data_291 ^ i_input_data[802 % IN_WIDTH];
                938 / IN_WIDTH: ping_storage_data_291 <= (fillup_transition == 1'b1) ? i_input_data[938 % IN_WIDTH] : ping_storage_data_291 ^ i_input_data[938 % IN_WIDTH];
                default: ping_storage_data_291 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_291;
                endcase
            end else begin
                case (input_count)
                38 / IN_WIDTH: pong_storage_data_291 <= (fillup_transition == 1'b1) ? i_input_data[38 % IN_WIDTH] : pong_storage_data_291 ^ i_input_data[38 % IN_WIDTH];
                244 / IN_WIDTH: pong_storage_data_291 <= (fillup_transition == 1'b1) ? i_input_data[244 % IN_WIDTH] : pong_storage_data_291 ^ i_input_data[244 % IN_WIDTH];
                802 / IN_WIDTH: pong_storage_data_291 <= (fillup_transition == 1'b1) ? i_input_data[802 % IN_WIDTH] : pong_storage_data_291 ^ i_input_data[802 % IN_WIDTH];
                938 / IN_WIDTH: pong_storage_data_291 <= (fillup_transition == 1'b1) ? i_input_data[938 % IN_WIDTH] : pong_storage_data_291 ^ i_input_data[938 % IN_WIDTH];
                default: pong_storage_data_291 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_291;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_291 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_291;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_291 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_291;
            end
        end
    end
end

logic ping_storage_data_292;
logic pong_storage_data_292;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_292 <= 1'b0;
        pong_storage_data_292 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                39 / IN_WIDTH: ping_storage_data_292 <= (fillup_transition == 1'b1) ? i_input_data[39 % IN_WIDTH] : ping_storage_data_292 ^ i_input_data[39 % IN_WIDTH];
                245 / IN_WIDTH: ping_storage_data_292 <= (fillup_transition == 1'b1) ? i_input_data[245 % IN_WIDTH] : ping_storage_data_292 ^ i_input_data[245 % IN_WIDTH];
                803 / IN_WIDTH: ping_storage_data_292 <= (fillup_transition == 1'b1) ? i_input_data[803 % IN_WIDTH] : ping_storage_data_292 ^ i_input_data[803 % IN_WIDTH];
                939 / IN_WIDTH: ping_storage_data_292 <= (fillup_transition == 1'b1) ? i_input_data[939 % IN_WIDTH] : ping_storage_data_292 ^ i_input_data[939 % IN_WIDTH];
                default: ping_storage_data_292 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_292;
                endcase
            end else begin
                case (input_count)
                39 / IN_WIDTH: pong_storage_data_292 <= (fillup_transition == 1'b1) ? i_input_data[39 % IN_WIDTH] : pong_storage_data_292 ^ i_input_data[39 % IN_WIDTH];
                245 / IN_WIDTH: pong_storage_data_292 <= (fillup_transition == 1'b1) ? i_input_data[245 % IN_WIDTH] : pong_storage_data_292 ^ i_input_data[245 % IN_WIDTH];
                803 / IN_WIDTH: pong_storage_data_292 <= (fillup_transition == 1'b1) ? i_input_data[803 % IN_WIDTH] : pong_storage_data_292 ^ i_input_data[803 % IN_WIDTH];
                939 / IN_WIDTH: pong_storage_data_292 <= (fillup_transition == 1'b1) ? i_input_data[939 % IN_WIDTH] : pong_storage_data_292 ^ i_input_data[939 % IN_WIDTH];
                default: pong_storage_data_292 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_292;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_292 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_292;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_292 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_292;
            end
        end
    end
end

logic ping_storage_data_293;
logic pong_storage_data_293;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_293 <= 1'b0;
        pong_storage_data_293 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                40 / IN_WIDTH: ping_storage_data_293 <= (fillup_transition == 1'b1) ? i_input_data[40 % IN_WIDTH] : ping_storage_data_293 ^ i_input_data[40 % IN_WIDTH];
                246 / IN_WIDTH: ping_storage_data_293 <= (fillup_transition == 1'b1) ? i_input_data[246 % IN_WIDTH] : ping_storage_data_293 ^ i_input_data[246 % IN_WIDTH];
                804 / IN_WIDTH: ping_storage_data_293 <= (fillup_transition == 1'b1) ? i_input_data[804 % IN_WIDTH] : ping_storage_data_293 ^ i_input_data[804 % IN_WIDTH];
                940 / IN_WIDTH: ping_storage_data_293 <= (fillup_transition == 1'b1) ? i_input_data[940 % IN_WIDTH] : ping_storage_data_293 ^ i_input_data[940 % IN_WIDTH];
                default: ping_storage_data_293 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_293;
                endcase
            end else begin
                case (input_count)
                40 / IN_WIDTH: pong_storage_data_293 <= (fillup_transition == 1'b1) ? i_input_data[40 % IN_WIDTH] : pong_storage_data_293 ^ i_input_data[40 % IN_WIDTH];
                246 / IN_WIDTH: pong_storage_data_293 <= (fillup_transition == 1'b1) ? i_input_data[246 % IN_WIDTH] : pong_storage_data_293 ^ i_input_data[246 % IN_WIDTH];
                804 / IN_WIDTH: pong_storage_data_293 <= (fillup_transition == 1'b1) ? i_input_data[804 % IN_WIDTH] : pong_storage_data_293 ^ i_input_data[804 % IN_WIDTH];
                940 / IN_WIDTH: pong_storage_data_293 <= (fillup_transition == 1'b1) ? i_input_data[940 % IN_WIDTH] : pong_storage_data_293 ^ i_input_data[940 % IN_WIDTH];
                default: pong_storage_data_293 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_293;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_293 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_293;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_293 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_293;
            end
        end
    end
end

logic ping_storage_data_294;
logic pong_storage_data_294;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_294 <= 1'b0;
        pong_storage_data_294 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                41 / IN_WIDTH: ping_storage_data_294 <= (fillup_transition == 1'b1) ? i_input_data[41 % IN_WIDTH] : ping_storage_data_294 ^ i_input_data[41 % IN_WIDTH];
                247 / IN_WIDTH: ping_storage_data_294 <= (fillup_transition == 1'b1) ? i_input_data[247 % IN_WIDTH] : ping_storage_data_294 ^ i_input_data[247 % IN_WIDTH];
                805 / IN_WIDTH: ping_storage_data_294 <= (fillup_transition == 1'b1) ? i_input_data[805 % IN_WIDTH] : ping_storage_data_294 ^ i_input_data[805 % IN_WIDTH];
                941 / IN_WIDTH: ping_storage_data_294 <= (fillup_transition == 1'b1) ? i_input_data[941 % IN_WIDTH] : ping_storage_data_294 ^ i_input_data[941 % IN_WIDTH];
                default: ping_storage_data_294 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_294;
                endcase
            end else begin
                case (input_count)
                41 / IN_WIDTH: pong_storage_data_294 <= (fillup_transition == 1'b1) ? i_input_data[41 % IN_WIDTH] : pong_storage_data_294 ^ i_input_data[41 % IN_WIDTH];
                247 / IN_WIDTH: pong_storage_data_294 <= (fillup_transition == 1'b1) ? i_input_data[247 % IN_WIDTH] : pong_storage_data_294 ^ i_input_data[247 % IN_WIDTH];
                805 / IN_WIDTH: pong_storage_data_294 <= (fillup_transition == 1'b1) ? i_input_data[805 % IN_WIDTH] : pong_storage_data_294 ^ i_input_data[805 % IN_WIDTH];
                941 / IN_WIDTH: pong_storage_data_294 <= (fillup_transition == 1'b1) ? i_input_data[941 % IN_WIDTH] : pong_storage_data_294 ^ i_input_data[941 % IN_WIDTH];
                default: pong_storage_data_294 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_294;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_294 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_294;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_294 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_294;
            end
        end
    end
end

logic ping_storage_data_295;
logic pong_storage_data_295;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_295 <= 1'b0;
        pong_storage_data_295 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                42 / IN_WIDTH: ping_storage_data_295 <= (fillup_transition == 1'b1) ? i_input_data[42 % IN_WIDTH] : ping_storage_data_295 ^ i_input_data[42 % IN_WIDTH];
                248 / IN_WIDTH: ping_storage_data_295 <= (fillup_transition == 1'b1) ? i_input_data[248 % IN_WIDTH] : ping_storage_data_295 ^ i_input_data[248 % IN_WIDTH];
                806 / IN_WIDTH: ping_storage_data_295 <= (fillup_transition == 1'b1) ? i_input_data[806 % IN_WIDTH] : ping_storage_data_295 ^ i_input_data[806 % IN_WIDTH];
                942 / IN_WIDTH: ping_storage_data_295 <= (fillup_transition == 1'b1) ? i_input_data[942 % IN_WIDTH] : ping_storage_data_295 ^ i_input_data[942 % IN_WIDTH];
                default: ping_storage_data_295 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_295;
                endcase
            end else begin
                case (input_count)
                42 / IN_WIDTH: pong_storage_data_295 <= (fillup_transition == 1'b1) ? i_input_data[42 % IN_WIDTH] : pong_storage_data_295 ^ i_input_data[42 % IN_WIDTH];
                248 / IN_WIDTH: pong_storage_data_295 <= (fillup_transition == 1'b1) ? i_input_data[248 % IN_WIDTH] : pong_storage_data_295 ^ i_input_data[248 % IN_WIDTH];
                806 / IN_WIDTH: pong_storage_data_295 <= (fillup_transition == 1'b1) ? i_input_data[806 % IN_WIDTH] : pong_storage_data_295 ^ i_input_data[806 % IN_WIDTH];
                942 / IN_WIDTH: pong_storage_data_295 <= (fillup_transition == 1'b1) ? i_input_data[942 % IN_WIDTH] : pong_storage_data_295 ^ i_input_data[942 % IN_WIDTH];
                default: pong_storage_data_295 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_295;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_295 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_295;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_295 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_295;
            end
        end
    end
end

logic ping_storage_data_296;
logic pong_storage_data_296;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_296 <= 1'b0;
        pong_storage_data_296 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                43 / IN_WIDTH: ping_storage_data_296 <= (fillup_transition == 1'b1) ? i_input_data[43 % IN_WIDTH] : ping_storage_data_296 ^ i_input_data[43 % IN_WIDTH];
                249 / IN_WIDTH: ping_storage_data_296 <= (fillup_transition == 1'b1) ? i_input_data[249 % IN_WIDTH] : ping_storage_data_296 ^ i_input_data[249 % IN_WIDTH];
                807 / IN_WIDTH: ping_storage_data_296 <= (fillup_transition == 1'b1) ? i_input_data[807 % IN_WIDTH] : ping_storage_data_296 ^ i_input_data[807 % IN_WIDTH];
                943 / IN_WIDTH: ping_storage_data_296 <= (fillup_transition == 1'b1) ? i_input_data[943 % IN_WIDTH] : ping_storage_data_296 ^ i_input_data[943 % IN_WIDTH];
                default: ping_storage_data_296 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_296;
                endcase
            end else begin
                case (input_count)
                43 / IN_WIDTH: pong_storage_data_296 <= (fillup_transition == 1'b1) ? i_input_data[43 % IN_WIDTH] : pong_storage_data_296 ^ i_input_data[43 % IN_WIDTH];
                249 / IN_WIDTH: pong_storage_data_296 <= (fillup_transition == 1'b1) ? i_input_data[249 % IN_WIDTH] : pong_storage_data_296 ^ i_input_data[249 % IN_WIDTH];
                807 / IN_WIDTH: pong_storage_data_296 <= (fillup_transition == 1'b1) ? i_input_data[807 % IN_WIDTH] : pong_storage_data_296 ^ i_input_data[807 % IN_WIDTH];
                943 / IN_WIDTH: pong_storage_data_296 <= (fillup_transition == 1'b1) ? i_input_data[943 % IN_WIDTH] : pong_storage_data_296 ^ i_input_data[943 % IN_WIDTH];
                default: pong_storage_data_296 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_296;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_296 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_296;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_296 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_296;
            end
        end
    end
end

logic ping_storage_data_297;
logic pong_storage_data_297;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_297 <= 1'b0;
        pong_storage_data_297 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                44 / IN_WIDTH: ping_storage_data_297 <= (fillup_transition == 1'b1) ? i_input_data[44 % IN_WIDTH] : ping_storage_data_297 ^ i_input_data[44 % IN_WIDTH];
                250 / IN_WIDTH: ping_storage_data_297 <= (fillup_transition == 1'b1) ? i_input_data[250 % IN_WIDTH] : ping_storage_data_297 ^ i_input_data[250 % IN_WIDTH];
                808 / IN_WIDTH: ping_storage_data_297 <= (fillup_transition == 1'b1) ? i_input_data[808 % IN_WIDTH] : ping_storage_data_297 ^ i_input_data[808 % IN_WIDTH];
                944 / IN_WIDTH: ping_storage_data_297 <= (fillup_transition == 1'b1) ? i_input_data[944 % IN_WIDTH] : ping_storage_data_297 ^ i_input_data[944 % IN_WIDTH];
                default: ping_storage_data_297 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_297;
                endcase
            end else begin
                case (input_count)
                44 / IN_WIDTH: pong_storage_data_297 <= (fillup_transition == 1'b1) ? i_input_data[44 % IN_WIDTH] : pong_storage_data_297 ^ i_input_data[44 % IN_WIDTH];
                250 / IN_WIDTH: pong_storage_data_297 <= (fillup_transition == 1'b1) ? i_input_data[250 % IN_WIDTH] : pong_storage_data_297 ^ i_input_data[250 % IN_WIDTH];
                808 / IN_WIDTH: pong_storage_data_297 <= (fillup_transition == 1'b1) ? i_input_data[808 % IN_WIDTH] : pong_storage_data_297 ^ i_input_data[808 % IN_WIDTH];
                944 / IN_WIDTH: pong_storage_data_297 <= (fillup_transition == 1'b1) ? i_input_data[944 % IN_WIDTH] : pong_storage_data_297 ^ i_input_data[944 % IN_WIDTH];
                default: pong_storage_data_297 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_297;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_297 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_297;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_297 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_297;
            end
        end
    end
end

logic ping_storage_data_298;
logic pong_storage_data_298;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_298 <= 1'b0;
        pong_storage_data_298 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                45 / IN_WIDTH: ping_storage_data_298 <= (fillup_transition == 1'b1) ? i_input_data[45 % IN_WIDTH] : ping_storage_data_298 ^ i_input_data[45 % IN_WIDTH];
                251 / IN_WIDTH: ping_storage_data_298 <= (fillup_transition == 1'b1) ? i_input_data[251 % IN_WIDTH] : ping_storage_data_298 ^ i_input_data[251 % IN_WIDTH];
                809 / IN_WIDTH: ping_storage_data_298 <= (fillup_transition == 1'b1) ? i_input_data[809 % IN_WIDTH] : ping_storage_data_298 ^ i_input_data[809 % IN_WIDTH];
                945 / IN_WIDTH: ping_storage_data_298 <= (fillup_transition == 1'b1) ? i_input_data[945 % IN_WIDTH] : ping_storage_data_298 ^ i_input_data[945 % IN_WIDTH];
                default: ping_storage_data_298 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_298;
                endcase
            end else begin
                case (input_count)
                45 / IN_WIDTH: pong_storage_data_298 <= (fillup_transition == 1'b1) ? i_input_data[45 % IN_WIDTH] : pong_storage_data_298 ^ i_input_data[45 % IN_WIDTH];
                251 / IN_WIDTH: pong_storage_data_298 <= (fillup_transition == 1'b1) ? i_input_data[251 % IN_WIDTH] : pong_storage_data_298 ^ i_input_data[251 % IN_WIDTH];
                809 / IN_WIDTH: pong_storage_data_298 <= (fillup_transition == 1'b1) ? i_input_data[809 % IN_WIDTH] : pong_storage_data_298 ^ i_input_data[809 % IN_WIDTH];
                945 / IN_WIDTH: pong_storage_data_298 <= (fillup_transition == 1'b1) ? i_input_data[945 % IN_WIDTH] : pong_storage_data_298 ^ i_input_data[945 % IN_WIDTH];
                default: pong_storage_data_298 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_298;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_298 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_298;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_298 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_298;
            end
        end
    end
end

logic ping_storage_data_299;
logic pong_storage_data_299;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_299 <= 1'b0;
        pong_storage_data_299 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                46 / IN_WIDTH: ping_storage_data_299 <= (fillup_transition == 1'b1) ? i_input_data[46 % IN_WIDTH] : ping_storage_data_299 ^ i_input_data[46 % IN_WIDTH];
                252 / IN_WIDTH: ping_storage_data_299 <= (fillup_transition == 1'b1) ? i_input_data[252 % IN_WIDTH] : ping_storage_data_299 ^ i_input_data[252 % IN_WIDTH];
                810 / IN_WIDTH: ping_storage_data_299 <= (fillup_transition == 1'b1) ? i_input_data[810 % IN_WIDTH] : ping_storage_data_299 ^ i_input_data[810 % IN_WIDTH];
                946 / IN_WIDTH: ping_storage_data_299 <= (fillup_transition == 1'b1) ? i_input_data[946 % IN_WIDTH] : ping_storage_data_299 ^ i_input_data[946 % IN_WIDTH];
                default: ping_storage_data_299 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_299;
                endcase
            end else begin
                case (input_count)
                46 / IN_WIDTH: pong_storage_data_299 <= (fillup_transition == 1'b1) ? i_input_data[46 % IN_WIDTH] : pong_storage_data_299 ^ i_input_data[46 % IN_WIDTH];
                252 / IN_WIDTH: pong_storage_data_299 <= (fillup_transition == 1'b1) ? i_input_data[252 % IN_WIDTH] : pong_storage_data_299 ^ i_input_data[252 % IN_WIDTH];
                810 / IN_WIDTH: pong_storage_data_299 <= (fillup_transition == 1'b1) ? i_input_data[810 % IN_WIDTH] : pong_storage_data_299 ^ i_input_data[810 % IN_WIDTH];
                946 / IN_WIDTH: pong_storage_data_299 <= (fillup_transition == 1'b1) ? i_input_data[946 % IN_WIDTH] : pong_storage_data_299 ^ i_input_data[946 % IN_WIDTH];
                default: pong_storage_data_299 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_299;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_299 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_299;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_299 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_299;
            end
        end
    end
end

logic ping_storage_data_300;
logic pong_storage_data_300;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_300 <= 1'b0;
        pong_storage_data_300 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                47 / IN_WIDTH: ping_storage_data_300 <= (fillup_transition == 1'b1) ? i_input_data[47 % IN_WIDTH] : ping_storage_data_300 ^ i_input_data[47 % IN_WIDTH];
                253 / IN_WIDTH: ping_storage_data_300 <= (fillup_transition == 1'b1) ? i_input_data[253 % IN_WIDTH] : ping_storage_data_300 ^ i_input_data[253 % IN_WIDTH];
                811 / IN_WIDTH: ping_storage_data_300 <= (fillup_transition == 1'b1) ? i_input_data[811 % IN_WIDTH] : ping_storage_data_300 ^ i_input_data[811 % IN_WIDTH];
                947 / IN_WIDTH: ping_storage_data_300 <= (fillup_transition == 1'b1) ? i_input_data[947 % IN_WIDTH] : ping_storage_data_300 ^ i_input_data[947 % IN_WIDTH];
                default: ping_storage_data_300 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_300;
                endcase
            end else begin
                case (input_count)
                47 / IN_WIDTH: pong_storage_data_300 <= (fillup_transition == 1'b1) ? i_input_data[47 % IN_WIDTH] : pong_storage_data_300 ^ i_input_data[47 % IN_WIDTH];
                253 / IN_WIDTH: pong_storage_data_300 <= (fillup_transition == 1'b1) ? i_input_data[253 % IN_WIDTH] : pong_storage_data_300 ^ i_input_data[253 % IN_WIDTH];
                811 / IN_WIDTH: pong_storage_data_300 <= (fillup_transition == 1'b1) ? i_input_data[811 % IN_WIDTH] : pong_storage_data_300 ^ i_input_data[811 % IN_WIDTH];
                947 / IN_WIDTH: pong_storage_data_300 <= (fillup_transition == 1'b1) ? i_input_data[947 % IN_WIDTH] : pong_storage_data_300 ^ i_input_data[947 % IN_WIDTH];
                default: pong_storage_data_300 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_300;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_300 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_300;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_300 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_300;
            end
        end
    end
end

logic ping_storage_data_301;
logic pong_storage_data_301;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_301 <= 1'b0;
        pong_storage_data_301 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                48 / IN_WIDTH: ping_storage_data_301 <= (fillup_transition == 1'b1) ? i_input_data[48 % IN_WIDTH] : ping_storage_data_301 ^ i_input_data[48 % IN_WIDTH];
                254 / IN_WIDTH: ping_storage_data_301 <= (fillup_transition == 1'b1) ? i_input_data[254 % IN_WIDTH] : ping_storage_data_301 ^ i_input_data[254 % IN_WIDTH];
                812 / IN_WIDTH: ping_storage_data_301 <= (fillup_transition == 1'b1) ? i_input_data[812 % IN_WIDTH] : ping_storage_data_301 ^ i_input_data[812 % IN_WIDTH];
                948 / IN_WIDTH: ping_storage_data_301 <= (fillup_transition == 1'b1) ? i_input_data[948 % IN_WIDTH] : ping_storage_data_301 ^ i_input_data[948 % IN_WIDTH];
                default: ping_storage_data_301 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_301;
                endcase
            end else begin
                case (input_count)
                48 / IN_WIDTH: pong_storage_data_301 <= (fillup_transition == 1'b1) ? i_input_data[48 % IN_WIDTH] : pong_storage_data_301 ^ i_input_data[48 % IN_WIDTH];
                254 / IN_WIDTH: pong_storage_data_301 <= (fillup_transition == 1'b1) ? i_input_data[254 % IN_WIDTH] : pong_storage_data_301 ^ i_input_data[254 % IN_WIDTH];
                812 / IN_WIDTH: pong_storage_data_301 <= (fillup_transition == 1'b1) ? i_input_data[812 % IN_WIDTH] : pong_storage_data_301 ^ i_input_data[812 % IN_WIDTH];
                948 / IN_WIDTH: pong_storage_data_301 <= (fillup_transition == 1'b1) ? i_input_data[948 % IN_WIDTH] : pong_storage_data_301 ^ i_input_data[948 % IN_WIDTH];
                default: pong_storage_data_301 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_301;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_301 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_301;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_301 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_301;
            end
        end
    end
end

logic ping_storage_data_302;
logic pong_storage_data_302;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_302 <= 1'b0;
        pong_storage_data_302 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                49 / IN_WIDTH: ping_storage_data_302 <= (fillup_transition == 1'b1) ? i_input_data[49 % IN_WIDTH] : ping_storage_data_302 ^ i_input_data[49 % IN_WIDTH];
                255 / IN_WIDTH: ping_storage_data_302 <= (fillup_transition == 1'b1) ? i_input_data[255 % IN_WIDTH] : ping_storage_data_302 ^ i_input_data[255 % IN_WIDTH];
                813 / IN_WIDTH: ping_storage_data_302 <= (fillup_transition == 1'b1) ? i_input_data[813 % IN_WIDTH] : ping_storage_data_302 ^ i_input_data[813 % IN_WIDTH];
                949 / IN_WIDTH: ping_storage_data_302 <= (fillup_transition == 1'b1) ? i_input_data[949 % IN_WIDTH] : ping_storage_data_302 ^ i_input_data[949 % IN_WIDTH];
                default: ping_storage_data_302 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_302;
                endcase
            end else begin
                case (input_count)
                49 / IN_WIDTH: pong_storage_data_302 <= (fillup_transition == 1'b1) ? i_input_data[49 % IN_WIDTH] : pong_storage_data_302 ^ i_input_data[49 % IN_WIDTH];
                255 / IN_WIDTH: pong_storage_data_302 <= (fillup_transition == 1'b1) ? i_input_data[255 % IN_WIDTH] : pong_storage_data_302 ^ i_input_data[255 % IN_WIDTH];
                813 / IN_WIDTH: pong_storage_data_302 <= (fillup_transition == 1'b1) ? i_input_data[813 % IN_WIDTH] : pong_storage_data_302 ^ i_input_data[813 % IN_WIDTH];
                949 / IN_WIDTH: pong_storage_data_302 <= (fillup_transition == 1'b1) ? i_input_data[949 % IN_WIDTH] : pong_storage_data_302 ^ i_input_data[949 % IN_WIDTH];
                default: pong_storage_data_302 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_302;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_302 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_302;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_302 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_302;
            end
        end
    end
end

logic ping_storage_data_303;
logic pong_storage_data_303;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_303 <= 1'b0;
        pong_storage_data_303 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                50 / IN_WIDTH: ping_storage_data_303 <= (fillup_transition == 1'b1) ? i_input_data[50 % IN_WIDTH] : ping_storage_data_303 ^ i_input_data[50 % IN_WIDTH];
                256 / IN_WIDTH: ping_storage_data_303 <= (fillup_transition == 1'b1) ? i_input_data[256 % IN_WIDTH] : ping_storage_data_303 ^ i_input_data[256 % IN_WIDTH];
                814 / IN_WIDTH: ping_storage_data_303 <= (fillup_transition == 1'b1) ? i_input_data[814 % IN_WIDTH] : ping_storage_data_303 ^ i_input_data[814 % IN_WIDTH];
                950 / IN_WIDTH: ping_storage_data_303 <= (fillup_transition == 1'b1) ? i_input_data[950 % IN_WIDTH] : ping_storage_data_303 ^ i_input_data[950 % IN_WIDTH];
                default: ping_storage_data_303 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_303;
                endcase
            end else begin
                case (input_count)
                50 / IN_WIDTH: pong_storage_data_303 <= (fillup_transition == 1'b1) ? i_input_data[50 % IN_WIDTH] : pong_storage_data_303 ^ i_input_data[50 % IN_WIDTH];
                256 / IN_WIDTH: pong_storage_data_303 <= (fillup_transition == 1'b1) ? i_input_data[256 % IN_WIDTH] : pong_storage_data_303 ^ i_input_data[256 % IN_WIDTH];
                814 / IN_WIDTH: pong_storage_data_303 <= (fillup_transition == 1'b1) ? i_input_data[814 % IN_WIDTH] : pong_storage_data_303 ^ i_input_data[814 % IN_WIDTH];
                950 / IN_WIDTH: pong_storage_data_303 <= (fillup_transition == 1'b1) ? i_input_data[950 % IN_WIDTH] : pong_storage_data_303 ^ i_input_data[950 % IN_WIDTH];
                default: pong_storage_data_303 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_303;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_303 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_303;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_303 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_303;
            end
        end
    end
end

logic ping_storage_data_304;
logic pong_storage_data_304;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_304 <= 1'b0;
        pong_storage_data_304 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                51 / IN_WIDTH: ping_storage_data_304 <= (fillup_transition == 1'b1) ? i_input_data[51 % IN_WIDTH] : ping_storage_data_304 ^ i_input_data[51 % IN_WIDTH];
                257 / IN_WIDTH: ping_storage_data_304 <= (fillup_transition == 1'b1) ? i_input_data[257 % IN_WIDTH] : ping_storage_data_304 ^ i_input_data[257 % IN_WIDTH];
                815 / IN_WIDTH: ping_storage_data_304 <= (fillup_transition == 1'b1) ? i_input_data[815 % IN_WIDTH] : ping_storage_data_304 ^ i_input_data[815 % IN_WIDTH];
                951 / IN_WIDTH: ping_storage_data_304 <= (fillup_transition == 1'b1) ? i_input_data[951 % IN_WIDTH] : ping_storage_data_304 ^ i_input_data[951 % IN_WIDTH];
                default: ping_storage_data_304 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_304;
                endcase
            end else begin
                case (input_count)
                51 / IN_WIDTH: pong_storage_data_304 <= (fillup_transition == 1'b1) ? i_input_data[51 % IN_WIDTH] : pong_storage_data_304 ^ i_input_data[51 % IN_WIDTH];
                257 / IN_WIDTH: pong_storage_data_304 <= (fillup_transition == 1'b1) ? i_input_data[257 % IN_WIDTH] : pong_storage_data_304 ^ i_input_data[257 % IN_WIDTH];
                815 / IN_WIDTH: pong_storage_data_304 <= (fillup_transition == 1'b1) ? i_input_data[815 % IN_WIDTH] : pong_storage_data_304 ^ i_input_data[815 % IN_WIDTH];
                951 / IN_WIDTH: pong_storage_data_304 <= (fillup_transition == 1'b1) ? i_input_data[951 % IN_WIDTH] : pong_storage_data_304 ^ i_input_data[951 % IN_WIDTH];
                default: pong_storage_data_304 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_304;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_304 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_304;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_304 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_304;
            end
        end
    end
end

logic ping_storage_data_305;
logic pong_storage_data_305;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_305 <= 1'b0;
        pong_storage_data_305 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                52 / IN_WIDTH: ping_storage_data_305 <= (fillup_transition == 1'b1) ? i_input_data[52 % IN_WIDTH] : ping_storage_data_305 ^ i_input_data[52 % IN_WIDTH];
                258 / IN_WIDTH: ping_storage_data_305 <= (fillup_transition == 1'b1) ? i_input_data[258 % IN_WIDTH] : ping_storage_data_305 ^ i_input_data[258 % IN_WIDTH];
                816 / IN_WIDTH: ping_storage_data_305 <= (fillup_transition == 1'b1) ? i_input_data[816 % IN_WIDTH] : ping_storage_data_305 ^ i_input_data[816 % IN_WIDTH];
                952 / IN_WIDTH: ping_storage_data_305 <= (fillup_transition == 1'b1) ? i_input_data[952 % IN_WIDTH] : ping_storage_data_305 ^ i_input_data[952 % IN_WIDTH];
                default: ping_storage_data_305 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_305;
                endcase
            end else begin
                case (input_count)
                52 / IN_WIDTH: pong_storage_data_305 <= (fillup_transition == 1'b1) ? i_input_data[52 % IN_WIDTH] : pong_storage_data_305 ^ i_input_data[52 % IN_WIDTH];
                258 / IN_WIDTH: pong_storage_data_305 <= (fillup_transition == 1'b1) ? i_input_data[258 % IN_WIDTH] : pong_storage_data_305 ^ i_input_data[258 % IN_WIDTH];
                816 / IN_WIDTH: pong_storage_data_305 <= (fillup_transition == 1'b1) ? i_input_data[816 % IN_WIDTH] : pong_storage_data_305 ^ i_input_data[816 % IN_WIDTH];
                952 / IN_WIDTH: pong_storage_data_305 <= (fillup_transition == 1'b1) ? i_input_data[952 % IN_WIDTH] : pong_storage_data_305 ^ i_input_data[952 % IN_WIDTH];
                default: pong_storage_data_305 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_305;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_305 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_305;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_305 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_305;
            end
        end
    end
end

logic ping_storage_data_306;
logic pong_storage_data_306;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_306 <= 1'b0;
        pong_storage_data_306 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                53 / IN_WIDTH: ping_storage_data_306 <= (fillup_transition == 1'b1) ? i_input_data[53 % IN_WIDTH] : ping_storage_data_306 ^ i_input_data[53 % IN_WIDTH];
                259 / IN_WIDTH: ping_storage_data_306 <= (fillup_transition == 1'b1) ? i_input_data[259 % IN_WIDTH] : ping_storage_data_306 ^ i_input_data[259 % IN_WIDTH];
                817 / IN_WIDTH: ping_storage_data_306 <= (fillup_transition == 1'b1) ? i_input_data[817 % IN_WIDTH] : ping_storage_data_306 ^ i_input_data[817 % IN_WIDTH];
                953 / IN_WIDTH: ping_storage_data_306 <= (fillup_transition == 1'b1) ? i_input_data[953 % IN_WIDTH] : ping_storage_data_306 ^ i_input_data[953 % IN_WIDTH];
                default: ping_storage_data_306 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_306;
                endcase
            end else begin
                case (input_count)
                53 / IN_WIDTH: pong_storage_data_306 <= (fillup_transition == 1'b1) ? i_input_data[53 % IN_WIDTH] : pong_storage_data_306 ^ i_input_data[53 % IN_WIDTH];
                259 / IN_WIDTH: pong_storage_data_306 <= (fillup_transition == 1'b1) ? i_input_data[259 % IN_WIDTH] : pong_storage_data_306 ^ i_input_data[259 % IN_WIDTH];
                817 / IN_WIDTH: pong_storage_data_306 <= (fillup_transition == 1'b1) ? i_input_data[817 % IN_WIDTH] : pong_storage_data_306 ^ i_input_data[817 % IN_WIDTH];
                953 / IN_WIDTH: pong_storage_data_306 <= (fillup_transition == 1'b1) ? i_input_data[953 % IN_WIDTH] : pong_storage_data_306 ^ i_input_data[953 % IN_WIDTH];
                default: pong_storage_data_306 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_306;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_306 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_306;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_306 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_306;
            end
        end
    end
end

logic ping_storage_data_307;
logic pong_storage_data_307;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_307 <= 1'b0;
        pong_storage_data_307 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                54 / IN_WIDTH: ping_storage_data_307 <= (fillup_transition == 1'b1) ? i_input_data[54 % IN_WIDTH] : ping_storage_data_307 ^ i_input_data[54 % IN_WIDTH];
                260 / IN_WIDTH: ping_storage_data_307 <= (fillup_transition == 1'b1) ? i_input_data[260 % IN_WIDTH] : ping_storage_data_307 ^ i_input_data[260 % IN_WIDTH];
                818 / IN_WIDTH: ping_storage_data_307 <= (fillup_transition == 1'b1) ? i_input_data[818 % IN_WIDTH] : ping_storage_data_307 ^ i_input_data[818 % IN_WIDTH];
                954 / IN_WIDTH: ping_storage_data_307 <= (fillup_transition == 1'b1) ? i_input_data[954 % IN_WIDTH] : ping_storage_data_307 ^ i_input_data[954 % IN_WIDTH];
                default: ping_storage_data_307 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_307;
                endcase
            end else begin
                case (input_count)
                54 / IN_WIDTH: pong_storage_data_307 <= (fillup_transition == 1'b1) ? i_input_data[54 % IN_WIDTH] : pong_storage_data_307 ^ i_input_data[54 % IN_WIDTH];
                260 / IN_WIDTH: pong_storage_data_307 <= (fillup_transition == 1'b1) ? i_input_data[260 % IN_WIDTH] : pong_storage_data_307 ^ i_input_data[260 % IN_WIDTH];
                818 / IN_WIDTH: pong_storage_data_307 <= (fillup_transition == 1'b1) ? i_input_data[818 % IN_WIDTH] : pong_storage_data_307 ^ i_input_data[818 % IN_WIDTH];
                954 / IN_WIDTH: pong_storage_data_307 <= (fillup_transition == 1'b1) ? i_input_data[954 % IN_WIDTH] : pong_storage_data_307 ^ i_input_data[954 % IN_WIDTH];
                default: pong_storage_data_307 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_307;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_307 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_307;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_307 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_307;
            end
        end
    end
end

logic ping_storage_data_308;
logic pong_storage_data_308;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_308 <= 1'b0;
        pong_storage_data_308 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                55 / IN_WIDTH: ping_storage_data_308 <= (fillup_transition == 1'b1) ? i_input_data[55 % IN_WIDTH] : ping_storage_data_308 ^ i_input_data[55 % IN_WIDTH];
                261 / IN_WIDTH: ping_storage_data_308 <= (fillup_transition == 1'b1) ? i_input_data[261 % IN_WIDTH] : ping_storage_data_308 ^ i_input_data[261 % IN_WIDTH];
                819 / IN_WIDTH: ping_storage_data_308 <= (fillup_transition == 1'b1) ? i_input_data[819 % IN_WIDTH] : ping_storage_data_308 ^ i_input_data[819 % IN_WIDTH];
                955 / IN_WIDTH: ping_storage_data_308 <= (fillup_transition == 1'b1) ? i_input_data[955 % IN_WIDTH] : ping_storage_data_308 ^ i_input_data[955 % IN_WIDTH];
                default: ping_storage_data_308 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_308;
                endcase
            end else begin
                case (input_count)
                55 / IN_WIDTH: pong_storage_data_308 <= (fillup_transition == 1'b1) ? i_input_data[55 % IN_WIDTH] : pong_storage_data_308 ^ i_input_data[55 % IN_WIDTH];
                261 / IN_WIDTH: pong_storage_data_308 <= (fillup_transition == 1'b1) ? i_input_data[261 % IN_WIDTH] : pong_storage_data_308 ^ i_input_data[261 % IN_WIDTH];
                819 / IN_WIDTH: pong_storage_data_308 <= (fillup_transition == 1'b1) ? i_input_data[819 % IN_WIDTH] : pong_storage_data_308 ^ i_input_data[819 % IN_WIDTH];
                955 / IN_WIDTH: pong_storage_data_308 <= (fillup_transition == 1'b1) ? i_input_data[955 % IN_WIDTH] : pong_storage_data_308 ^ i_input_data[955 % IN_WIDTH];
                default: pong_storage_data_308 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_308;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_308 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_308;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_308 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_308;
            end
        end
    end
end

logic ping_storage_data_309;
logic pong_storage_data_309;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_309 <= 1'b0;
        pong_storage_data_309 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                56 / IN_WIDTH: ping_storage_data_309 <= (fillup_transition == 1'b1) ? i_input_data[56 % IN_WIDTH] : ping_storage_data_309 ^ i_input_data[56 % IN_WIDTH];
                262 / IN_WIDTH: ping_storage_data_309 <= (fillup_transition == 1'b1) ? i_input_data[262 % IN_WIDTH] : ping_storage_data_309 ^ i_input_data[262 % IN_WIDTH];
                820 / IN_WIDTH: ping_storage_data_309 <= (fillup_transition == 1'b1) ? i_input_data[820 % IN_WIDTH] : ping_storage_data_309 ^ i_input_data[820 % IN_WIDTH];
                956 / IN_WIDTH: ping_storage_data_309 <= (fillup_transition == 1'b1) ? i_input_data[956 % IN_WIDTH] : ping_storage_data_309 ^ i_input_data[956 % IN_WIDTH];
                default: ping_storage_data_309 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_309;
                endcase
            end else begin
                case (input_count)
                56 / IN_WIDTH: pong_storage_data_309 <= (fillup_transition == 1'b1) ? i_input_data[56 % IN_WIDTH] : pong_storage_data_309 ^ i_input_data[56 % IN_WIDTH];
                262 / IN_WIDTH: pong_storage_data_309 <= (fillup_transition == 1'b1) ? i_input_data[262 % IN_WIDTH] : pong_storage_data_309 ^ i_input_data[262 % IN_WIDTH];
                820 / IN_WIDTH: pong_storage_data_309 <= (fillup_transition == 1'b1) ? i_input_data[820 % IN_WIDTH] : pong_storage_data_309 ^ i_input_data[820 % IN_WIDTH];
                956 / IN_WIDTH: pong_storage_data_309 <= (fillup_transition == 1'b1) ? i_input_data[956 % IN_WIDTH] : pong_storage_data_309 ^ i_input_data[956 % IN_WIDTH];
                default: pong_storage_data_309 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_309;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_309 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_309;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_309 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_309;
            end
        end
    end
end

logic ping_storage_data_310;
logic pong_storage_data_310;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_310 <= 1'b0;
        pong_storage_data_310 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                57 / IN_WIDTH: ping_storage_data_310 <= (fillup_transition == 1'b1) ? i_input_data[57 % IN_WIDTH] : ping_storage_data_310 ^ i_input_data[57 % IN_WIDTH];
                263 / IN_WIDTH: ping_storage_data_310 <= (fillup_transition == 1'b1) ? i_input_data[263 % IN_WIDTH] : ping_storage_data_310 ^ i_input_data[263 % IN_WIDTH];
                821 / IN_WIDTH: ping_storage_data_310 <= (fillup_transition == 1'b1) ? i_input_data[821 % IN_WIDTH] : ping_storage_data_310 ^ i_input_data[821 % IN_WIDTH];
                957 / IN_WIDTH: ping_storage_data_310 <= (fillup_transition == 1'b1) ? i_input_data[957 % IN_WIDTH] : ping_storage_data_310 ^ i_input_data[957 % IN_WIDTH];
                default: ping_storage_data_310 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_310;
                endcase
            end else begin
                case (input_count)
                57 / IN_WIDTH: pong_storage_data_310 <= (fillup_transition == 1'b1) ? i_input_data[57 % IN_WIDTH] : pong_storage_data_310 ^ i_input_data[57 % IN_WIDTH];
                263 / IN_WIDTH: pong_storage_data_310 <= (fillup_transition == 1'b1) ? i_input_data[263 % IN_WIDTH] : pong_storage_data_310 ^ i_input_data[263 % IN_WIDTH];
                821 / IN_WIDTH: pong_storage_data_310 <= (fillup_transition == 1'b1) ? i_input_data[821 % IN_WIDTH] : pong_storage_data_310 ^ i_input_data[821 % IN_WIDTH];
                957 / IN_WIDTH: pong_storage_data_310 <= (fillup_transition == 1'b1) ? i_input_data[957 % IN_WIDTH] : pong_storage_data_310 ^ i_input_data[957 % IN_WIDTH];
                default: pong_storage_data_310 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_310;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_310 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_310;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_310 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_310;
            end
        end
    end
end

logic ping_storage_data_311;
logic pong_storage_data_311;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_311 <= 1'b0;
        pong_storage_data_311 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                58 / IN_WIDTH: ping_storage_data_311 <= (fillup_transition == 1'b1) ? i_input_data[58 % IN_WIDTH] : ping_storage_data_311 ^ i_input_data[58 % IN_WIDTH];
                264 / IN_WIDTH: ping_storage_data_311 <= (fillup_transition == 1'b1) ? i_input_data[264 % IN_WIDTH] : ping_storage_data_311 ^ i_input_data[264 % IN_WIDTH];
                822 / IN_WIDTH: ping_storage_data_311 <= (fillup_transition == 1'b1) ? i_input_data[822 % IN_WIDTH] : ping_storage_data_311 ^ i_input_data[822 % IN_WIDTH];
                958 / IN_WIDTH: ping_storage_data_311 <= (fillup_transition == 1'b1) ? i_input_data[958 % IN_WIDTH] : ping_storage_data_311 ^ i_input_data[958 % IN_WIDTH];
                default: ping_storage_data_311 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_311;
                endcase
            end else begin
                case (input_count)
                58 / IN_WIDTH: pong_storage_data_311 <= (fillup_transition == 1'b1) ? i_input_data[58 % IN_WIDTH] : pong_storage_data_311 ^ i_input_data[58 % IN_WIDTH];
                264 / IN_WIDTH: pong_storage_data_311 <= (fillup_transition == 1'b1) ? i_input_data[264 % IN_WIDTH] : pong_storage_data_311 ^ i_input_data[264 % IN_WIDTH];
                822 / IN_WIDTH: pong_storage_data_311 <= (fillup_transition == 1'b1) ? i_input_data[822 % IN_WIDTH] : pong_storage_data_311 ^ i_input_data[822 % IN_WIDTH];
                958 / IN_WIDTH: pong_storage_data_311 <= (fillup_transition == 1'b1) ? i_input_data[958 % IN_WIDTH] : pong_storage_data_311 ^ i_input_data[958 % IN_WIDTH];
                default: pong_storage_data_311 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_311;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_311 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_311;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_311 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_311;
            end
        end
    end
end

logic ping_storage_data_312;
logic pong_storage_data_312;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_312 <= 1'b0;
        pong_storage_data_312 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                59 / IN_WIDTH: ping_storage_data_312 <= (fillup_transition == 1'b1) ? i_input_data[59 % IN_WIDTH] : ping_storage_data_312 ^ i_input_data[59 % IN_WIDTH];
                265 / IN_WIDTH: ping_storage_data_312 <= (fillup_transition == 1'b1) ? i_input_data[265 % IN_WIDTH] : ping_storage_data_312 ^ i_input_data[265 % IN_WIDTH];
                823 / IN_WIDTH: ping_storage_data_312 <= (fillup_transition == 1'b1) ? i_input_data[823 % IN_WIDTH] : ping_storage_data_312 ^ i_input_data[823 % IN_WIDTH];
                959 / IN_WIDTH: ping_storage_data_312 <= (fillup_transition == 1'b1) ? i_input_data[959 % IN_WIDTH] : ping_storage_data_312 ^ i_input_data[959 % IN_WIDTH];
                default: ping_storage_data_312 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_312;
                endcase
            end else begin
                case (input_count)
                59 / IN_WIDTH: pong_storage_data_312 <= (fillup_transition == 1'b1) ? i_input_data[59 % IN_WIDTH] : pong_storage_data_312 ^ i_input_data[59 % IN_WIDTH];
                265 / IN_WIDTH: pong_storage_data_312 <= (fillup_transition == 1'b1) ? i_input_data[265 % IN_WIDTH] : pong_storage_data_312 ^ i_input_data[265 % IN_WIDTH];
                823 / IN_WIDTH: pong_storage_data_312 <= (fillup_transition == 1'b1) ? i_input_data[823 % IN_WIDTH] : pong_storage_data_312 ^ i_input_data[823 % IN_WIDTH];
                959 / IN_WIDTH: pong_storage_data_312 <= (fillup_transition == 1'b1) ? i_input_data[959 % IN_WIDTH] : pong_storage_data_312 ^ i_input_data[959 % IN_WIDTH];
                default: pong_storage_data_312 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_312;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_312 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_312;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_312 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_312;
            end
        end
    end
end

logic ping_storage_data_313;
logic pong_storage_data_313;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_313 <= 1'b0;
        pong_storage_data_313 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                60 / IN_WIDTH: ping_storage_data_313 <= (fillup_transition == 1'b1) ? i_input_data[60 % IN_WIDTH] : ping_storage_data_313 ^ i_input_data[60 % IN_WIDTH];
                266 / IN_WIDTH: ping_storage_data_313 <= (fillup_transition == 1'b1) ? i_input_data[266 % IN_WIDTH] : ping_storage_data_313 ^ i_input_data[266 % IN_WIDTH];
                824 / IN_WIDTH: ping_storage_data_313 <= (fillup_transition == 1'b1) ? i_input_data[824 % IN_WIDTH] : ping_storage_data_313 ^ i_input_data[824 % IN_WIDTH];
                864 / IN_WIDTH: ping_storage_data_313 <= (fillup_transition == 1'b1) ? i_input_data[864 % IN_WIDTH] : ping_storage_data_313 ^ i_input_data[864 % IN_WIDTH];
                default: ping_storage_data_313 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_313;
                endcase
            end else begin
                case (input_count)
                60 / IN_WIDTH: pong_storage_data_313 <= (fillup_transition == 1'b1) ? i_input_data[60 % IN_WIDTH] : pong_storage_data_313 ^ i_input_data[60 % IN_WIDTH];
                266 / IN_WIDTH: pong_storage_data_313 <= (fillup_transition == 1'b1) ? i_input_data[266 % IN_WIDTH] : pong_storage_data_313 ^ i_input_data[266 % IN_WIDTH];
                824 / IN_WIDTH: pong_storage_data_313 <= (fillup_transition == 1'b1) ? i_input_data[824 % IN_WIDTH] : pong_storage_data_313 ^ i_input_data[824 % IN_WIDTH];
                864 / IN_WIDTH: pong_storage_data_313 <= (fillup_transition == 1'b1) ? i_input_data[864 % IN_WIDTH] : pong_storage_data_313 ^ i_input_data[864 % IN_WIDTH];
                default: pong_storage_data_313 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_313;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_313 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_313;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_313 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_313;
            end
        end
    end
end

logic ping_storage_data_314;
logic pong_storage_data_314;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_314 <= 1'b0;
        pong_storage_data_314 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                61 / IN_WIDTH: ping_storage_data_314 <= (fillup_transition == 1'b1) ? i_input_data[61 % IN_WIDTH] : ping_storage_data_314 ^ i_input_data[61 % IN_WIDTH];
                267 / IN_WIDTH: ping_storage_data_314 <= (fillup_transition == 1'b1) ? i_input_data[267 % IN_WIDTH] : ping_storage_data_314 ^ i_input_data[267 % IN_WIDTH];
                825 / IN_WIDTH: ping_storage_data_314 <= (fillup_transition == 1'b1) ? i_input_data[825 % IN_WIDTH] : ping_storage_data_314 ^ i_input_data[825 % IN_WIDTH];
                865 / IN_WIDTH: ping_storage_data_314 <= (fillup_transition == 1'b1) ? i_input_data[865 % IN_WIDTH] : ping_storage_data_314 ^ i_input_data[865 % IN_WIDTH];
                default: ping_storage_data_314 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_314;
                endcase
            end else begin
                case (input_count)
                61 / IN_WIDTH: pong_storage_data_314 <= (fillup_transition == 1'b1) ? i_input_data[61 % IN_WIDTH] : pong_storage_data_314 ^ i_input_data[61 % IN_WIDTH];
                267 / IN_WIDTH: pong_storage_data_314 <= (fillup_transition == 1'b1) ? i_input_data[267 % IN_WIDTH] : pong_storage_data_314 ^ i_input_data[267 % IN_WIDTH];
                825 / IN_WIDTH: pong_storage_data_314 <= (fillup_transition == 1'b1) ? i_input_data[825 % IN_WIDTH] : pong_storage_data_314 ^ i_input_data[825 % IN_WIDTH];
                865 / IN_WIDTH: pong_storage_data_314 <= (fillup_transition == 1'b1) ? i_input_data[865 % IN_WIDTH] : pong_storage_data_314 ^ i_input_data[865 % IN_WIDTH];
                default: pong_storage_data_314 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_314;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_314 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_314;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_314 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_314;
            end
        end
    end
end

logic ping_storage_data_315;
logic pong_storage_data_315;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_315 <= 1'b0;
        pong_storage_data_315 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                62 / IN_WIDTH: ping_storage_data_315 <= (fillup_transition == 1'b1) ? i_input_data[62 % IN_WIDTH] : ping_storage_data_315 ^ i_input_data[62 % IN_WIDTH];
                268 / IN_WIDTH: ping_storage_data_315 <= (fillup_transition == 1'b1) ? i_input_data[268 % IN_WIDTH] : ping_storage_data_315 ^ i_input_data[268 % IN_WIDTH];
                826 / IN_WIDTH: ping_storage_data_315 <= (fillup_transition == 1'b1) ? i_input_data[826 % IN_WIDTH] : ping_storage_data_315 ^ i_input_data[826 % IN_WIDTH];
                866 / IN_WIDTH: ping_storage_data_315 <= (fillup_transition == 1'b1) ? i_input_data[866 % IN_WIDTH] : ping_storage_data_315 ^ i_input_data[866 % IN_WIDTH];
                default: ping_storage_data_315 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_315;
                endcase
            end else begin
                case (input_count)
                62 / IN_WIDTH: pong_storage_data_315 <= (fillup_transition == 1'b1) ? i_input_data[62 % IN_WIDTH] : pong_storage_data_315 ^ i_input_data[62 % IN_WIDTH];
                268 / IN_WIDTH: pong_storage_data_315 <= (fillup_transition == 1'b1) ? i_input_data[268 % IN_WIDTH] : pong_storage_data_315 ^ i_input_data[268 % IN_WIDTH];
                826 / IN_WIDTH: pong_storage_data_315 <= (fillup_transition == 1'b1) ? i_input_data[826 % IN_WIDTH] : pong_storage_data_315 ^ i_input_data[826 % IN_WIDTH];
                866 / IN_WIDTH: pong_storage_data_315 <= (fillup_transition == 1'b1) ? i_input_data[866 % IN_WIDTH] : pong_storage_data_315 ^ i_input_data[866 % IN_WIDTH];
                default: pong_storage_data_315 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_315;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_315 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_315;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_315 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_315;
            end
        end
    end
end

logic ping_storage_data_316;
logic pong_storage_data_316;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_316 <= 1'b0;
        pong_storage_data_316 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                63 / IN_WIDTH: ping_storage_data_316 <= (fillup_transition == 1'b1) ? i_input_data[63 % IN_WIDTH] : ping_storage_data_316 ^ i_input_data[63 % IN_WIDTH];
                269 / IN_WIDTH: ping_storage_data_316 <= (fillup_transition == 1'b1) ? i_input_data[269 % IN_WIDTH] : ping_storage_data_316 ^ i_input_data[269 % IN_WIDTH];
                827 / IN_WIDTH: ping_storage_data_316 <= (fillup_transition == 1'b1) ? i_input_data[827 % IN_WIDTH] : ping_storage_data_316 ^ i_input_data[827 % IN_WIDTH];
                867 / IN_WIDTH: ping_storage_data_316 <= (fillup_transition == 1'b1) ? i_input_data[867 % IN_WIDTH] : ping_storage_data_316 ^ i_input_data[867 % IN_WIDTH];
                default: ping_storage_data_316 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_316;
                endcase
            end else begin
                case (input_count)
                63 / IN_WIDTH: pong_storage_data_316 <= (fillup_transition == 1'b1) ? i_input_data[63 % IN_WIDTH] : pong_storage_data_316 ^ i_input_data[63 % IN_WIDTH];
                269 / IN_WIDTH: pong_storage_data_316 <= (fillup_transition == 1'b1) ? i_input_data[269 % IN_WIDTH] : pong_storage_data_316 ^ i_input_data[269 % IN_WIDTH];
                827 / IN_WIDTH: pong_storage_data_316 <= (fillup_transition == 1'b1) ? i_input_data[827 % IN_WIDTH] : pong_storage_data_316 ^ i_input_data[827 % IN_WIDTH];
                867 / IN_WIDTH: pong_storage_data_316 <= (fillup_transition == 1'b1) ? i_input_data[867 % IN_WIDTH] : pong_storage_data_316 ^ i_input_data[867 % IN_WIDTH];
                default: pong_storage_data_316 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_316;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_316 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_316;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_316 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_316;
            end
        end
    end
end

logic ping_storage_data_317;
logic pong_storage_data_317;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_317 <= 1'b0;
        pong_storage_data_317 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                64 / IN_WIDTH: ping_storage_data_317 <= (fillup_transition == 1'b1) ? i_input_data[64 % IN_WIDTH] : ping_storage_data_317 ^ i_input_data[64 % IN_WIDTH];
                270 / IN_WIDTH: ping_storage_data_317 <= (fillup_transition == 1'b1) ? i_input_data[270 % IN_WIDTH] : ping_storage_data_317 ^ i_input_data[270 % IN_WIDTH];
                828 / IN_WIDTH: ping_storage_data_317 <= (fillup_transition == 1'b1) ? i_input_data[828 % IN_WIDTH] : ping_storage_data_317 ^ i_input_data[828 % IN_WIDTH];
                868 / IN_WIDTH: ping_storage_data_317 <= (fillup_transition == 1'b1) ? i_input_data[868 % IN_WIDTH] : ping_storage_data_317 ^ i_input_data[868 % IN_WIDTH];
                default: ping_storage_data_317 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_317;
                endcase
            end else begin
                case (input_count)
                64 / IN_WIDTH: pong_storage_data_317 <= (fillup_transition == 1'b1) ? i_input_data[64 % IN_WIDTH] : pong_storage_data_317 ^ i_input_data[64 % IN_WIDTH];
                270 / IN_WIDTH: pong_storage_data_317 <= (fillup_transition == 1'b1) ? i_input_data[270 % IN_WIDTH] : pong_storage_data_317 ^ i_input_data[270 % IN_WIDTH];
                828 / IN_WIDTH: pong_storage_data_317 <= (fillup_transition == 1'b1) ? i_input_data[828 % IN_WIDTH] : pong_storage_data_317 ^ i_input_data[828 % IN_WIDTH];
                868 / IN_WIDTH: pong_storage_data_317 <= (fillup_transition == 1'b1) ? i_input_data[868 % IN_WIDTH] : pong_storage_data_317 ^ i_input_data[868 % IN_WIDTH];
                default: pong_storage_data_317 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_317;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_317 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_317;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_317 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_317;
            end
        end
    end
end

logic ping_storage_data_318;
logic pong_storage_data_318;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_318 <= 1'b0;
        pong_storage_data_318 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                65 / IN_WIDTH: ping_storage_data_318 <= (fillup_transition == 1'b1) ? i_input_data[65 % IN_WIDTH] : ping_storage_data_318 ^ i_input_data[65 % IN_WIDTH];
                271 / IN_WIDTH: ping_storage_data_318 <= (fillup_transition == 1'b1) ? i_input_data[271 % IN_WIDTH] : ping_storage_data_318 ^ i_input_data[271 % IN_WIDTH];
                829 / IN_WIDTH: ping_storage_data_318 <= (fillup_transition == 1'b1) ? i_input_data[829 % IN_WIDTH] : ping_storage_data_318 ^ i_input_data[829 % IN_WIDTH];
                869 / IN_WIDTH: ping_storage_data_318 <= (fillup_transition == 1'b1) ? i_input_data[869 % IN_WIDTH] : ping_storage_data_318 ^ i_input_data[869 % IN_WIDTH];
                default: ping_storage_data_318 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_318;
                endcase
            end else begin
                case (input_count)
                65 / IN_WIDTH: pong_storage_data_318 <= (fillup_transition == 1'b1) ? i_input_data[65 % IN_WIDTH] : pong_storage_data_318 ^ i_input_data[65 % IN_WIDTH];
                271 / IN_WIDTH: pong_storage_data_318 <= (fillup_transition == 1'b1) ? i_input_data[271 % IN_WIDTH] : pong_storage_data_318 ^ i_input_data[271 % IN_WIDTH];
                829 / IN_WIDTH: pong_storage_data_318 <= (fillup_transition == 1'b1) ? i_input_data[829 % IN_WIDTH] : pong_storage_data_318 ^ i_input_data[829 % IN_WIDTH];
                869 / IN_WIDTH: pong_storage_data_318 <= (fillup_transition == 1'b1) ? i_input_data[869 % IN_WIDTH] : pong_storage_data_318 ^ i_input_data[869 % IN_WIDTH];
                default: pong_storage_data_318 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_318;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_318 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_318;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_318 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_318;
            end
        end
    end
end

logic ping_storage_data_319;
logic pong_storage_data_319;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_319 <= 1'b0;
        pong_storage_data_319 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                66 / IN_WIDTH: ping_storage_data_319 <= (fillup_transition == 1'b1) ? i_input_data[66 % IN_WIDTH] : ping_storage_data_319 ^ i_input_data[66 % IN_WIDTH];
                272 / IN_WIDTH: ping_storage_data_319 <= (fillup_transition == 1'b1) ? i_input_data[272 % IN_WIDTH] : ping_storage_data_319 ^ i_input_data[272 % IN_WIDTH];
                830 / IN_WIDTH: ping_storage_data_319 <= (fillup_transition == 1'b1) ? i_input_data[830 % IN_WIDTH] : ping_storage_data_319 ^ i_input_data[830 % IN_WIDTH];
                870 / IN_WIDTH: ping_storage_data_319 <= (fillup_transition == 1'b1) ? i_input_data[870 % IN_WIDTH] : ping_storage_data_319 ^ i_input_data[870 % IN_WIDTH];
                default: ping_storage_data_319 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_319;
                endcase
            end else begin
                case (input_count)
                66 / IN_WIDTH: pong_storage_data_319 <= (fillup_transition == 1'b1) ? i_input_data[66 % IN_WIDTH] : pong_storage_data_319 ^ i_input_data[66 % IN_WIDTH];
                272 / IN_WIDTH: pong_storage_data_319 <= (fillup_transition == 1'b1) ? i_input_data[272 % IN_WIDTH] : pong_storage_data_319 ^ i_input_data[272 % IN_WIDTH];
                830 / IN_WIDTH: pong_storage_data_319 <= (fillup_transition == 1'b1) ? i_input_data[830 % IN_WIDTH] : pong_storage_data_319 ^ i_input_data[830 % IN_WIDTH];
                870 / IN_WIDTH: pong_storage_data_319 <= (fillup_transition == 1'b1) ? i_input_data[870 % IN_WIDTH] : pong_storage_data_319 ^ i_input_data[870 % IN_WIDTH];
                default: pong_storage_data_319 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_319;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_319 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_319;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_319 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_319;
            end
        end
    end
end

logic ping_storage_data_320;
logic pong_storage_data_320;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_320 <= 1'b0;
        pong_storage_data_320 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                67 / IN_WIDTH: ping_storage_data_320 <= (fillup_transition == 1'b1) ? i_input_data[67 % IN_WIDTH] : ping_storage_data_320 ^ i_input_data[67 % IN_WIDTH];
                273 / IN_WIDTH: ping_storage_data_320 <= (fillup_transition == 1'b1) ? i_input_data[273 % IN_WIDTH] : ping_storage_data_320 ^ i_input_data[273 % IN_WIDTH];
                831 / IN_WIDTH: ping_storage_data_320 <= (fillup_transition == 1'b1) ? i_input_data[831 % IN_WIDTH] : ping_storage_data_320 ^ i_input_data[831 % IN_WIDTH];
                871 / IN_WIDTH: ping_storage_data_320 <= (fillup_transition == 1'b1) ? i_input_data[871 % IN_WIDTH] : ping_storage_data_320 ^ i_input_data[871 % IN_WIDTH];
                default: ping_storage_data_320 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_320;
                endcase
            end else begin
                case (input_count)
                67 / IN_WIDTH: pong_storage_data_320 <= (fillup_transition == 1'b1) ? i_input_data[67 % IN_WIDTH] : pong_storage_data_320 ^ i_input_data[67 % IN_WIDTH];
                273 / IN_WIDTH: pong_storage_data_320 <= (fillup_transition == 1'b1) ? i_input_data[273 % IN_WIDTH] : pong_storage_data_320 ^ i_input_data[273 % IN_WIDTH];
                831 / IN_WIDTH: pong_storage_data_320 <= (fillup_transition == 1'b1) ? i_input_data[831 % IN_WIDTH] : pong_storage_data_320 ^ i_input_data[831 % IN_WIDTH];
                871 / IN_WIDTH: pong_storage_data_320 <= (fillup_transition == 1'b1) ? i_input_data[871 % IN_WIDTH] : pong_storage_data_320 ^ i_input_data[871 % IN_WIDTH];
                default: pong_storage_data_320 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_320;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_320 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_320;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_320 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_320;
            end
        end
    end
end

logic ping_storage_data_321;
logic pong_storage_data_321;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_321 <= 1'b0;
        pong_storage_data_321 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                68 / IN_WIDTH: ping_storage_data_321 <= (fillup_transition == 1'b1) ? i_input_data[68 % IN_WIDTH] : ping_storage_data_321 ^ i_input_data[68 % IN_WIDTH];
                274 / IN_WIDTH: ping_storage_data_321 <= (fillup_transition == 1'b1) ? i_input_data[274 % IN_WIDTH] : ping_storage_data_321 ^ i_input_data[274 % IN_WIDTH];
                832 / IN_WIDTH: ping_storage_data_321 <= (fillup_transition == 1'b1) ? i_input_data[832 % IN_WIDTH] : ping_storage_data_321 ^ i_input_data[832 % IN_WIDTH];
                872 / IN_WIDTH: ping_storage_data_321 <= (fillup_transition == 1'b1) ? i_input_data[872 % IN_WIDTH] : ping_storage_data_321 ^ i_input_data[872 % IN_WIDTH];
                default: ping_storage_data_321 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_321;
                endcase
            end else begin
                case (input_count)
                68 / IN_WIDTH: pong_storage_data_321 <= (fillup_transition == 1'b1) ? i_input_data[68 % IN_WIDTH] : pong_storage_data_321 ^ i_input_data[68 % IN_WIDTH];
                274 / IN_WIDTH: pong_storage_data_321 <= (fillup_transition == 1'b1) ? i_input_data[274 % IN_WIDTH] : pong_storage_data_321 ^ i_input_data[274 % IN_WIDTH];
                832 / IN_WIDTH: pong_storage_data_321 <= (fillup_transition == 1'b1) ? i_input_data[832 % IN_WIDTH] : pong_storage_data_321 ^ i_input_data[832 % IN_WIDTH];
                872 / IN_WIDTH: pong_storage_data_321 <= (fillup_transition == 1'b1) ? i_input_data[872 % IN_WIDTH] : pong_storage_data_321 ^ i_input_data[872 % IN_WIDTH];
                default: pong_storage_data_321 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_321;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_321 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_321;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_321 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_321;
            end
        end
    end
end

logic ping_storage_data_322;
logic pong_storage_data_322;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_322 <= 1'b0;
        pong_storage_data_322 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                69 / IN_WIDTH: ping_storage_data_322 <= (fillup_transition == 1'b1) ? i_input_data[69 % IN_WIDTH] : ping_storage_data_322 ^ i_input_data[69 % IN_WIDTH];
                275 / IN_WIDTH: ping_storage_data_322 <= (fillup_transition == 1'b1) ? i_input_data[275 % IN_WIDTH] : ping_storage_data_322 ^ i_input_data[275 % IN_WIDTH];
                833 / IN_WIDTH: ping_storage_data_322 <= (fillup_transition == 1'b1) ? i_input_data[833 % IN_WIDTH] : ping_storage_data_322 ^ i_input_data[833 % IN_WIDTH];
                873 / IN_WIDTH: ping_storage_data_322 <= (fillup_transition == 1'b1) ? i_input_data[873 % IN_WIDTH] : ping_storage_data_322 ^ i_input_data[873 % IN_WIDTH];
                default: ping_storage_data_322 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_322;
                endcase
            end else begin
                case (input_count)
                69 / IN_WIDTH: pong_storage_data_322 <= (fillup_transition == 1'b1) ? i_input_data[69 % IN_WIDTH] : pong_storage_data_322 ^ i_input_data[69 % IN_WIDTH];
                275 / IN_WIDTH: pong_storage_data_322 <= (fillup_transition == 1'b1) ? i_input_data[275 % IN_WIDTH] : pong_storage_data_322 ^ i_input_data[275 % IN_WIDTH];
                833 / IN_WIDTH: pong_storage_data_322 <= (fillup_transition == 1'b1) ? i_input_data[833 % IN_WIDTH] : pong_storage_data_322 ^ i_input_data[833 % IN_WIDTH];
                873 / IN_WIDTH: pong_storage_data_322 <= (fillup_transition == 1'b1) ? i_input_data[873 % IN_WIDTH] : pong_storage_data_322 ^ i_input_data[873 % IN_WIDTH];
                default: pong_storage_data_322 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_322;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_322 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_322;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_322 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_322;
            end
        end
    end
end

logic ping_storage_data_323;
logic pong_storage_data_323;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_323 <= 1'b0;
        pong_storage_data_323 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                70 / IN_WIDTH: ping_storage_data_323 <= (fillup_transition == 1'b1) ? i_input_data[70 % IN_WIDTH] : ping_storage_data_323 ^ i_input_data[70 % IN_WIDTH];
                276 / IN_WIDTH: ping_storage_data_323 <= (fillup_transition == 1'b1) ? i_input_data[276 % IN_WIDTH] : ping_storage_data_323 ^ i_input_data[276 % IN_WIDTH];
                834 / IN_WIDTH: ping_storage_data_323 <= (fillup_transition == 1'b1) ? i_input_data[834 % IN_WIDTH] : ping_storage_data_323 ^ i_input_data[834 % IN_WIDTH];
                874 / IN_WIDTH: ping_storage_data_323 <= (fillup_transition == 1'b1) ? i_input_data[874 % IN_WIDTH] : ping_storage_data_323 ^ i_input_data[874 % IN_WIDTH];
                default: ping_storage_data_323 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_323;
                endcase
            end else begin
                case (input_count)
                70 / IN_WIDTH: pong_storage_data_323 <= (fillup_transition == 1'b1) ? i_input_data[70 % IN_WIDTH] : pong_storage_data_323 ^ i_input_data[70 % IN_WIDTH];
                276 / IN_WIDTH: pong_storage_data_323 <= (fillup_transition == 1'b1) ? i_input_data[276 % IN_WIDTH] : pong_storage_data_323 ^ i_input_data[276 % IN_WIDTH];
                834 / IN_WIDTH: pong_storage_data_323 <= (fillup_transition == 1'b1) ? i_input_data[834 % IN_WIDTH] : pong_storage_data_323 ^ i_input_data[834 % IN_WIDTH];
                874 / IN_WIDTH: pong_storage_data_323 <= (fillup_transition == 1'b1) ? i_input_data[874 % IN_WIDTH] : pong_storage_data_323 ^ i_input_data[874 % IN_WIDTH];
                default: pong_storage_data_323 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_323;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_323 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_323;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_323 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_323;
            end
        end
    end
end

logic ping_storage_data_324;
logic pong_storage_data_324;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_324 <= 1'b0;
        pong_storage_data_324 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                71 / IN_WIDTH: ping_storage_data_324 <= (fillup_transition == 1'b1) ? i_input_data[71 % IN_WIDTH] : ping_storage_data_324 ^ i_input_data[71 % IN_WIDTH];
                277 / IN_WIDTH: ping_storage_data_324 <= (fillup_transition == 1'b1) ? i_input_data[277 % IN_WIDTH] : ping_storage_data_324 ^ i_input_data[277 % IN_WIDTH];
                835 / IN_WIDTH: ping_storage_data_324 <= (fillup_transition == 1'b1) ? i_input_data[835 % IN_WIDTH] : ping_storage_data_324 ^ i_input_data[835 % IN_WIDTH];
                875 / IN_WIDTH: ping_storage_data_324 <= (fillup_transition == 1'b1) ? i_input_data[875 % IN_WIDTH] : ping_storage_data_324 ^ i_input_data[875 % IN_WIDTH];
                default: ping_storage_data_324 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_324;
                endcase
            end else begin
                case (input_count)
                71 / IN_WIDTH: pong_storage_data_324 <= (fillup_transition == 1'b1) ? i_input_data[71 % IN_WIDTH] : pong_storage_data_324 ^ i_input_data[71 % IN_WIDTH];
                277 / IN_WIDTH: pong_storage_data_324 <= (fillup_transition == 1'b1) ? i_input_data[277 % IN_WIDTH] : pong_storage_data_324 ^ i_input_data[277 % IN_WIDTH];
                835 / IN_WIDTH: pong_storage_data_324 <= (fillup_transition == 1'b1) ? i_input_data[835 % IN_WIDTH] : pong_storage_data_324 ^ i_input_data[835 % IN_WIDTH];
                875 / IN_WIDTH: pong_storage_data_324 <= (fillup_transition == 1'b1) ? i_input_data[875 % IN_WIDTH] : pong_storage_data_324 ^ i_input_data[875 % IN_WIDTH];
                default: pong_storage_data_324 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_324;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_324 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_324;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_324 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_324;
            end
        end
    end
end

logic ping_storage_data_325;
logic pong_storage_data_325;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_325 <= 1'b0;
        pong_storage_data_325 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                72 / IN_WIDTH: ping_storage_data_325 <= (fillup_transition == 1'b1) ? i_input_data[72 % IN_WIDTH] : ping_storage_data_325 ^ i_input_data[72 % IN_WIDTH];
                278 / IN_WIDTH: ping_storage_data_325 <= (fillup_transition == 1'b1) ? i_input_data[278 % IN_WIDTH] : ping_storage_data_325 ^ i_input_data[278 % IN_WIDTH];
                836 / IN_WIDTH: ping_storage_data_325 <= (fillup_transition == 1'b1) ? i_input_data[836 % IN_WIDTH] : ping_storage_data_325 ^ i_input_data[836 % IN_WIDTH];
                876 / IN_WIDTH: ping_storage_data_325 <= (fillup_transition == 1'b1) ? i_input_data[876 % IN_WIDTH] : ping_storage_data_325 ^ i_input_data[876 % IN_WIDTH];
                default: ping_storage_data_325 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_325;
                endcase
            end else begin
                case (input_count)
                72 / IN_WIDTH: pong_storage_data_325 <= (fillup_transition == 1'b1) ? i_input_data[72 % IN_WIDTH] : pong_storage_data_325 ^ i_input_data[72 % IN_WIDTH];
                278 / IN_WIDTH: pong_storage_data_325 <= (fillup_transition == 1'b1) ? i_input_data[278 % IN_WIDTH] : pong_storage_data_325 ^ i_input_data[278 % IN_WIDTH];
                836 / IN_WIDTH: pong_storage_data_325 <= (fillup_transition == 1'b1) ? i_input_data[836 % IN_WIDTH] : pong_storage_data_325 ^ i_input_data[836 % IN_WIDTH];
                876 / IN_WIDTH: pong_storage_data_325 <= (fillup_transition == 1'b1) ? i_input_data[876 % IN_WIDTH] : pong_storage_data_325 ^ i_input_data[876 % IN_WIDTH];
                default: pong_storage_data_325 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_325;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_325 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_325;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_325 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_325;
            end
        end
    end
end

logic ping_storage_data_326;
logic pong_storage_data_326;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_326 <= 1'b0;
        pong_storage_data_326 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                73 / IN_WIDTH: ping_storage_data_326 <= (fillup_transition == 1'b1) ? i_input_data[73 % IN_WIDTH] : ping_storage_data_326 ^ i_input_data[73 % IN_WIDTH];
                279 / IN_WIDTH: ping_storage_data_326 <= (fillup_transition == 1'b1) ? i_input_data[279 % IN_WIDTH] : ping_storage_data_326 ^ i_input_data[279 % IN_WIDTH];
                837 / IN_WIDTH: ping_storage_data_326 <= (fillup_transition == 1'b1) ? i_input_data[837 % IN_WIDTH] : ping_storage_data_326 ^ i_input_data[837 % IN_WIDTH];
                877 / IN_WIDTH: ping_storage_data_326 <= (fillup_transition == 1'b1) ? i_input_data[877 % IN_WIDTH] : ping_storage_data_326 ^ i_input_data[877 % IN_WIDTH];
                default: ping_storage_data_326 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_326;
                endcase
            end else begin
                case (input_count)
                73 / IN_WIDTH: pong_storage_data_326 <= (fillup_transition == 1'b1) ? i_input_data[73 % IN_WIDTH] : pong_storage_data_326 ^ i_input_data[73 % IN_WIDTH];
                279 / IN_WIDTH: pong_storage_data_326 <= (fillup_transition == 1'b1) ? i_input_data[279 % IN_WIDTH] : pong_storage_data_326 ^ i_input_data[279 % IN_WIDTH];
                837 / IN_WIDTH: pong_storage_data_326 <= (fillup_transition == 1'b1) ? i_input_data[837 % IN_WIDTH] : pong_storage_data_326 ^ i_input_data[837 % IN_WIDTH];
                877 / IN_WIDTH: pong_storage_data_326 <= (fillup_transition == 1'b1) ? i_input_data[877 % IN_WIDTH] : pong_storage_data_326 ^ i_input_data[877 % IN_WIDTH];
                default: pong_storage_data_326 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_326;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_326 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_326;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_326 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_326;
            end
        end
    end
end

logic ping_storage_data_327;
logic pong_storage_data_327;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_327 <= 1'b0;
        pong_storage_data_327 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                74 / IN_WIDTH: ping_storage_data_327 <= (fillup_transition == 1'b1) ? i_input_data[74 % IN_WIDTH] : ping_storage_data_327 ^ i_input_data[74 % IN_WIDTH];
                280 / IN_WIDTH: ping_storage_data_327 <= (fillup_transition == 1'b1) ? i_input_data[280 % IN_WIDTH] : ping_storage_data_327 ^ i_input_data[280 % IN_WIDTH];
                838 / IN_WIDTH: ping_storage_data_327 <= (fillup_transition == 1'b1) ? i_input_data[838 % IN_WIDTH] : ping_storage_data_327 ^ i_input_data[838 % IN_WIDTH];
                878 / IN_WIDTH: ping_storage_data_327 <= (fillup_transition == 1'b1) ? i_input_data[878 % IN_WIDTH] : ping_storage_data_327 ^ i_input_data[878 % IN_WIDTH];
                default: ping_storage_data_327 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_327;
                endcase
            end else begin
                case (input_count)
                74 / IN_WIDTH: pong_storage_data_327 <= (fillup_transition == 1'b1) ? i_input_data[74 % IN_WIDTH] : pong_storage_data_327 ^ i_input_data[74 % IN_WIDTH];
                280 / IN_WIDTH: pong_storage_data_327 <= (fillup_transition == 1'b1) ? i_input_data[280 % IN_WIDTH] : pong_storage_data_327 ^ i_input_data[280 % IN_WIDTH];
                838 / IN_WIDTH: pong_storage_data_327 <= (fillup_transition == 1'b1) ? i_input_data[838 % IN_WIDTH] : pong_storage_data_327 ^ i_input_data[838 % IN_WIDTH];
                878 / IN_WIDTH: pong_storage_data_327 <= (fillup_transition == 1'b1) ? i_input_data[878 % IN_WIDTH] : pong_storage_data_327 ^ i_input_data[878 % IN_WIDTH];
                default: pong_storage_data_327 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_327;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_327 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_327;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_327 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_327;
            end
        end
    end
end

logic ping_storage_data_328;
logic pong_storage_data_328;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_328 <= 1'b0;
        pong_storage_data_328 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                75 / IN_WIDTH: ping_storage_data_328 <= (fillup_transition == 1'b1) ? i_input_data[75 % IN_WIDTH] : ping_storage_data_328 ^ i_input_data[75 % IN_WIDTH];
                281 / IN_WIDTH: ping_storage_data_328 <= (fillup_transition == 1'b1) ? i_input_data[281 % IN_WIDTH] : ping_storage_data_328 ^ i_input_data[281 % IN_WIDTH];
                839 / IN_WIDTH: ping_storage_data_328 <= (fillup_transition == 1'b1) ? i_input_data[839 % IN_WIDTH] : ping_storage_data_328 ^ i_input_data[839 % IN_WIDTH];
                879 / IN_WIDTH: ping_storage_data_328 <= (fillup_transition == 1'b1) ? i_input_data[879 % IN_WIDTH] : ping_storage_data_328 ^ i_input_data[879 % IN_WIDTH];
                default: ping_storage_data_328 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_328;
                endcase
            end else begin
                case (input_count)
                75 / IN_WIDTH: pong_storage_data_328 <= (fillup_transition == 1'b1) ? i_input_data[75 % IN_WIDTH] : pong_storage_data_328 ^ i_input_data[75 % IN_WIDTH];
                281 / IN_WIDTH: pong_storage_data_328 <= (fillup_transition == 1'b1) ? i_input_data[281 % IN_WIDTH] : pong_storage_data_328 ^ i_input_data[281 % IN_WIDTH];
                839 / IN_WIDTH: pong_storage_data_328 <= (fillup_transition == 1'b1) ? i_input_data[839 % IN_WIDTH] : pong_storage_data_328 ^ i_input_data[839 % IN_WIDTH];
                879 / IN_WIDTH: pong_storage_data_328 <= (fillup_transition == 1'b1) ? i_input_data[879 % IN_WIDTH] : pong_storage_data_328 ^ i_input_data[879 % IN_WIDTH];
                default: pong_storage_data_328 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_328;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_328 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_328;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_328 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_328;
            end
        end
    end
end

logic ping_storage_data_329;
logic pong_storage_data_329;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_329 <= 1'b0;
        pong_storage_data_329 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                76 / IN_WIDTH: ping_storage_data_329 <= (fillup_transition == 1'b1) ? i_input_data[76 % IN_WIDTH] : ping_storage_data_329 ^ i_input_data[76 % IN_WIDTH];
                282 / IN_WIDTH: ping_storage_data_329 <= (fillup_transition == 1'b1) ? i_input_data[282 % IN_WIDTH] : ping_storage_data_329 ^ i_input_data[282 % IN_WIDTH];
                840 / IN_WIDTH: ping_storage_data_329 <= (fillup_transition == 1'b1) ? i_input_data[840 % IN_WIDTH] : ping_storage_data_329 ^ i_input_data[840 % IN_WIDTH];
                880 / IN_WIDTH: ping_storage_data_329 <= (fillup_transition == 1'b1) ? i_input_data[880 % IN_WIDTH] : ping_storage_data_329 ^ i_input_data[880 % IN_WIDTH];
                default: ping_storage_data_329 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_329;
                endcase
            end else begin
                case (input_count)
                76 / IN_WIDTH: pong_storage_data_329 <= (fillup_transition == 1'b1) ? i_input_data[76 % IN_WIDTH] : pong_storage_data_329 ^ i_input_data[76 % IN_WIDTH];
                282 / IN_WIDTH: pong_storage_data_329 <= (fillup_transition == 1'b1) ? i_input_data[282 % IN_WIDTH] : pong_storage_data_329 ^ i_input_data[282 % IN_WIDTH];
                840 / IN_WIDTH: pong_storage_data_329 <= (fillup_transition == 1'b1) ? i_input_data[840 % IN_WIDTH] : pong_storage_data_329 ^ i_input_data[840 % IN_WIDTH];
                880 / IN_WIDTH: pong_storage_data_329 <= (fillup_transition == 1'b1) ? i_input_data[880 % IN_WIDTH] : pong_storage_data_329 ^ i_input_data[880 % IN_WIDTH];
                default: pong_storage_data_329 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_329;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_329 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_329;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_329 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_329;
            end
        end
    end
end

logic ping_storage_data_330;
logic pong_storage_data_330;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_330 <= 1'b0;
        pong_storage_data_330 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                77 / IN_WIDTH: ping_storage_data_330 <= (fillup_transition == 1'b1) ? i_input_data[77 % IN_WIDTH] : ping_storage_data_330 ^ i_input_data[77 % IN_WIDTH];
                283 / IN_WIDTH: ping_storage_data_330 <= (fillup_transition == 1'b1) ? i_input_data[283 % IN_WIDTH] : ping_storage_data_330 ^ i_input_data[283 % IN_WIDTH];
                841 / IN_WIDTH: ping_storage_data_330 <= (fillup_transition == 1'b1) ? i_input_data[841 % IN_WIDTH] : ping_storage_data_330 ^ i_input_data[841 % IN_WIDTH];
                881 / IN_WIDTH: ping_storage_data_330 <= (fillup_transition == 1'b1) ? i_input_data[881 % IN_WIDTH] : ping_storage_data_330 ^ i_input_data[881 % IN_WIDTH];
                default: ping_storage_data_330 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_330;
                endcase
            end else begin
                case (input_count)
                77 / IN_WIDTH: pong_storage_data_330 <= (fillup_transition == 1'b1) ? i_input_data[77 % IN_WIDTH] : pong_storage_data_330 ^ i_input_data[77 % IN_WIDTH];
                283 / IN_WIDTH: pong_storage_data_330 <= (fillup_transition == 1'b1) ? i_input_data[283 % IN_WIDTH] : pong_storage_data_330 ^ i_input_data[283 % IN_WIDTH];
                841 / IN_WIDTH: pong_storage_data_330 <= (fillup_transition == 1'b1) ? i_input_data[841 % IN_WIDTH] : pong_storage_data_330 ^ i_input_data[841 % IN_WIDTH];
                881 / IN_WIDTH: pong_storage_data_330 <= (fillup_transition == 1'b1) ? i_input_data[881 % IN_WIDTH] : pong_storage_data_330 ^ i_input_data[881 % IN_WIDTH];
                default: pong_storage_data_330 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_330;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_330 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_330;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_330 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_330;
            end
        end
    end
end

logic ping_storage_data_331;
logic pong_storage_data_331;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_331 <= 1'b0;
        pong_storage_data_331 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                78 / IN_WIDTH: ping_storage_data_331 <= (fillup_transition == 1'b1) ? i_input_data[78 % IN_WIDTH] : ping_storage_data_331 ^ i_input_data[78 % IN_WIDTH];
                284 / IN_WIDTH: ping_storage_data_331 <= (fillup_transition == 1'b1) ? i_input_data[284 % IN_WIDTH] : ping_storage_data_331 ^ i_input_data[284 % IN_WIDTH];
                842 / IN_WIDTH: ping_storage_data_331 <= (fillup_transition == 1'b1) ? i_input_data[842 % IN_WIDTH] : ping_storage_data_331 ^ i_input_data[842 % IN_WIDTH];
                882 / IN_WIDTH: ping_storage_data_331 <= (fillup_transition == 1'b1) ? i_input_data[882 % IN_WIDTH] : ping_storage_data_331 ^ i_input_data[882 % IN_WIDTH];
                default: ping_storage_data_331 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_331;
                endcase
            end else begin
                case (input_count)
                78 / IN_WIDTH: pong_storage_data_331 <= (fillup_transition == 1'b1) ? i_input_data[78 % IN_WIDTH] : pong_storage_data_331 ^ i_input_data[78 % IN_WIDTH];
                284 / IN_WIDTH: pong_storage_data_331 <= (fillup_transition == 1'b1) ? i_input_data[284 % IN_WIDTH] : pong_storage_data_331 ^ i_input_data[284 % IN_WIDTH];
                842 / IN_WIDTH: pong_storage_data_331 <= (fillup_transition == 1'b1) ? i_input_data[842 % IN_WIDTH] : pong_storage_data_331 ^ i_input_data[842 % IN_WIDTH];
                882 / IN_WIDTH: pong_storage_data_331 <= (fillup_transition == 1'b1) ? i_input_data[882 % IN_WIDTH] : pong_storage_data_331 ^ i_input_data[882 % IN_WIDTH];
                default: pong_storage_data_331 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_331;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_331 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_331;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_331 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_331;
            end
        end
    end
end

logic ping_storage_data_332;
logic pong_storage_data_332;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_332 <= 1'b0;
        pong_storage_data_332 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                79 / IN_WIDTH: ping_storage_data_332 <= (fillup_transition == 1'b1) ? i_input_data[79 % IN_WIDTH] : ping_storage_data_332 ^ i_input_data[79 % IN_WIDTH];
                285 / IN_WIDTH: ping_storage_data_332 <= (fillup_transition == 1'b1) ? i_input_data[285 % IN_WIDTH] : ping_storage_data_332 ^ i_input_data[285 % IN_WIDTH];
                843 / IN_WIDTH: ping_storage_data_332 <= (fillup_transition == 1'b1) ? i_input_data[843 % IN_WIDTH] : ping_storage_data_332 ^ i_input_data[843 % IN_WIDTH];
                883 / IN_WIDTH: ping_storage_data_332 <= (fillup_transition == 1'b1) ? i_input_data[883 % IN_WIDTH] : ping_storage_data_332 ^ i_input_data[883 % IN_WIDTH];
                default: ping_storage_data_332 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_332;
                endcase
            end else begin
                case (input_count)
                79 / IN_WIDTH: pong_storage_data_332 <= (fillup_transition == 1'b1) ? i_input_data[79 % IN_WIDTH] : pong_storage_data_332 ^ i_input_data[79 % IN_WIDTH];
                285 / IN_WIDTH: pong_storage_data_332 <= (fillup_transition == 1'b1) ? i_input_data[285 % IN_WIDTH] : pong_storage_data_332 ^ i_input_data[285 % IN_WIDTH];
                843 / IN_WIDTH: pong_storage_data_332 <= (fillup_transition == 1'b1) ? i_input_data[843 % IN_WIDTH] : pong_storage_data_332 ^ i_input_data[843 % IN_WIDTH];
                883 / IN_WIDTH: pong_storage_data_332 <= (fillup_transition == 1'b1) ? i_input_data[883 % IN_WIDTH] : pong_storage_data_332 ^ i_input_data[883 % IN_WIDTH];
                default: pong_storage_data_332 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_332;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_332 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_332;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_332 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_332;
            end
        end
    end
end

logic ping_storage_data_333;
logic pong_storage_data_333;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_333 <= 1'b0;
        pong_storage_data_333 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                80 / IN_WIDTH: ping_storage_data_333 <= (fillup_transition == 1'b1) ? i_input_data[80 % IN_WIDTH] : ping_storage_data_333 ^ i_input_data[80 % IN_WIDTH];
                286 / IN_WIDTH: ping_storage_data_333 <= (fillup_transition == 1'b1) ? i_input_data[286 % IN_WIDTH] : ping_storage_data_333 ^ i_input_data[286 % IN_WIDTH];
                844 / IN_WIDTH: ping_storage_data_333 <= (fillup_transition == 1'b1) ? i_input_data[844 % IN_WIDTH] : ping_storage_data_333 ^ i_input_data[844 % IN_WIDTH];
                884 / IN_WIDTH: ping_storage_data_333 <= (fillup_transition == 1'b1) ? i_input_data[884 % IN_WIDTH] : ping_storage_data_333 ^ i_input_data[884 % IN_WIDTH];
                default: ping_storage_data_333 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_333;
                endcase
            end else begin
                case (input_count)
                80 / IN_WIDTH: pong_storage_data_333 <= (fillup_transition == 1'b1) ? i_input_data[80 % IN_WIDTH] : pong_storage_data_333 ^ i_input_data[80 % IN_WIDTH];
                286 / IN_WIDTH: pong_storage_data_333 <= (fillup_transition == 1'b1) ? i_input_data[286 % IN_WIDTH] : pong_storage_data_333 ^ i_input_data[286 % IN_WIDTH];
                844 / IN_WIDTH: pong_storage_data_333 <= (fillup_transition == 1'b1) ? i_input_data[844 % IN_WIDTH] : pong_storage_data_333 ^ i_input_data[844 % IN_WIDTH];
                884 / IN_WIDTH: pong_storage_data_333 <= (fillup_transition == 1'b1) ? i_input_data[884 % IN_WIDTH] : pong_storage_data_333 ^ i_input_data[884 % IN_WIDTH];
                default: pong_storage_data_333 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_333;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_333 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_333;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_333 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_333;
            end
        end
    end
end

logic ping_storage_data_334;
logic pong_storage_data_334;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_334 <= 1'b0;
        pong_storage_data_334 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                81 / IN_WIDTH: ping_storage_data_334 <= (fillup_transition == 1'b1) ? i_input_data[81 % IN_WIDTH] : ping_storage_data_334 ^ i_input_data[81 % IN_WIDTH];
                287 / IN_WIDTH: ping_storage_data_334 <= (fillup_transition == 1'b1) ? i_input_data[287 % IN_WIDTH] : ping_storage_data_334 ^ i_input_data[287 % IN_WIDTH];
                845 / IN_WIDTH: ping_storage_data_334 <= (fillup_transition == 1'b1) ? i_input_data[845 % IN_WIDTH] : ping_storage_data_334 ^ i_input_data[845 % IN_WIDTH];
                885 / IN_WIDTH: ping_storage_data_334 <= (fillup_transition == 1'b1) ? i_input_data[885 % IN_WIDTH] : ping_storage_data_334 ^ i_input_data[885 % IN_WIDTH];
                default: ping_storage_data_334 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_334;
                endcase
            end else begin
                case (input_count)
                81 / IN_WIDTH: pong_storage_data_334 <= (fillup_transition == 1'b1) ? i_input_data[81 % IN_WIDTH] : pong_storage_data_334 ^ i_input_data[81 % IN_WIDTH];
                287 / IN_WIDTH: pong_storage_data_334 <= (fillup_transition == 1'b1) ? i_input_data[287 % IN_WIDTH] : pong_storage_data_334 ^ i_input_data[287 % IN_WIDTH];
                845 / IN_WIDTH: pong_storage_data_334 <= (fillup_transition == 1'b1) ? i_input_data[845 % IN_WIDTH] : pong_storage_data_334 ^ i_input_data[845 % IN_WIDTH];
                885 / IN_WIDTH: pong_storage_data_334 <= (fillup_transition == 1'b1) ? i_input_data[885 % IN_WIDTH] : pong_storage_data_334 ^ i_input_data[885 % IN_WIDTH];
                default: pong_storage_data_334 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_334;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_334 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_334;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_334 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_334;
            end
        end
    end
end

logic ping_storage_data_335;
logic pong_storage_data_335;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_335 <= 1'b0;
        pong_storage_data_335 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                82 / IN_WIDTH: ping_storage_data_335 <= (fillup_transition == 1'b1) ? i_input_data[82 % IN_WIDTH] : ping_storage_data_335 ^ i_input_data[82 % IN_WIDTH];
                192 / IN_WIDTH: ping_storage_data_335 <= (fillup_transition == 1'b1) ? i_input_data[192 % IN_WIDTH] : ping_storage_data_335 ^ i_input_data[192 % IN_WIDTH];
                846 / IN_WIDTH: ping_storage_data_335 <= (fillup_transition == 1'b1) ? i_input_data[846 % IN_WIDTH] : ping_storage_data_335 ^ i_input_data[846 % IN_WIDTH];
                886 / IN_WIDTH: ping_storage_data_335 <= (fillup_transition == 1'b1) ? i_input_data[886 % IN_WIDTH] : ping_storage_data_335 ^ i_input_data[886 % IN_WIDTH];
                default: ping_storage_data_335 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_335;
                endcase
            end else begin
                case (input_count)
                82 / IN_WIDTH: pong_storage_data_335 <= (fillup_transition == 1'b1) ? i_input_data[82 % IN_WIDTH] : pong_storage_data_335 ^ i_input_data[82 % IN_WIDTH];
                192 / IN_WIDTH: pong_storage_data_335 <= (fillup_transition == 1'b1) ? i_input_data[192 % IN_WIDTH] : pong_storage_data_335 ^ i_input_data[192 % IN_WIDTH];
                846 / IN_WIDTH: pong_storage_data_335 <= (fillup_transition == 1'b1) ? i_input_data[846 % IN_WIDTH] : pong_storage_data_335 ^ i_input_data[846 % IN_WIDTH];
                886 / IN_WIDTH: pong_storage_data_335 <= (fillup_transition == 1'b1) ? i_input_data[886 % IN_WIDTH] : pong_storage_data_335 ^ i_input_data[886 % IN_WIDTH];
                default: pong_storage_data_335 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_335;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_335 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_335;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_335 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_335;
            end
        end
    end
end

logic ping_storage_data_336;
logic pong_storage_data_336;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_336 <= 1'b0;
        pong_storage_data_336 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                83 / IN_WIDTH: ping_storage_data_336 <= (fillup_transition == 1'b1) ? i_input_data[83 % IN_WIDTH] : ping_storage_data_336 ^ i_input_data[83 % IN_WIDTH];
                193 / IN_WIDTH: ping_storage_data_336 <= (fillup_transition == 1'b1) ? i_input_data[193 % IN_WIDTH] : ping_storage_data_336 ^ i_input_data[193 % IN_WIDTH];
                847 / IN_WIDTH: ping_storage_data_336 <= (fillup_transition == 1'b1) ? i_input_data[847 % IN_WIDTH] : ping_storage_data_336 ^ i_input_data[847 % IN_WIDTH];
                887 / IN_WIDTH: ping_storage_data_336 <= (fillup_transition == 1'b1) ? i_input_data[887 % IN_WIDTH] : ping_storage_data_336 ^ i_input_data[887 % IN_WIDTH];
                default: ping_storage_data_336 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_336;
                endcase
            end else begin
                case (input_count)
                83 / IN_WIDTH: pong_storage_data_336 <= (fillup_transition == 1'b1) ? i_input_data[83 % IN_WIDTH] : pong_storage_data_336 ^ i_input_data[83 % IN_WIDTH];
                193 / IN_WIDTH: pong_storage_data_336 <= (fillup_transition == 1'b1) ? i_input_data[193 % IN_WIDTH] : pong_storage_data_336 ^ i_input_data[193 % IN_WIDTH];
                847 / IN_WIDTH: pong_storage_data_336 <= (fillup_transition == 1'b1) ? i_input_data[847 % IN_WIDTH] : pong_storage_data_336 ^ i_input_data[847 % IN_WIDTH];
                887 / IN_WIDTH: pong_storage_data_336 <= (fillup_transition == 1'b1) ? i_input_data[887 % IN_WIDTH] : pong_storage_data_336 ^ i_input_data[887 % IN_WIDTH];
                default: pong_storage_data_336 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_336;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_336 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_336;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_336 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_336;
            end
        end
    end
end

logic ping_storage_data_337;
logic pong_storage_data_337;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_337 <= 1'b0;
        pong_storage_data_337 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                84 / IN_WIDTH: ping_storage_data_337 <= (fillup_transition == 1'b1) ? i_input_data[84 % IN_WIDTH] : ping_storage_data_337 ^ i_input_data[84 % IN_WIDTH];
                194 / IN_WIDTH: ping_storage_data_337 <= (fillup_transition == 1'b1) ? i_input_data[194 % IN_WIDTH] : ping_storage_data_337 ^ i_input_data[194 % IN_WIDTH];
                848 / IN_WIDTH: ping_storage_data_337 <= (fillup_transition == 1'b1) ? i_input_data[848 % IN_WIDTH] : ping_storage_data_337 ^ i_input_data[848 % IN_WIDTH];
                888 / IN_WIDTH: ping_storage_data_337 <= (fillup_transition == 1'b1) ? i_input_data[888 % IN_WIDTH] : ping_storage_data_337 ^ i_input_data[888 % IN_WIDTH];
                default: ping_storage_data_337 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_337;
                endcase
            end else begin
                case (input_count)
                84 / IN_WIDTH: pong_storage_data_337 <= (fillup_transition == 1'b1) ? i_input_data[84 % IN_WIDTH] : pong_storage_data_337 ^ i_input_data[84 % IN_WIDTH];
                194 / IN_WIDTH: pong_storage_data_337 <= (fillup_transition == 1'b1) ? i_input_data[194 % IN_WIDTH] : pong_storage_data_337 ^ i_input_data[194 % IN_WIDTH];
                848 / IN_WIDTH: pong_storage_data_337 <= (fillup_transition == 1'b1) ? i_input_data[848 % IN_WIDTH] : pong_storage_data_337 ^ i_input_data[848 % IN_WIDTH];
                888 / IN_WIDTH: pong_storage_data_337 <= (fillup_transition == 1'b1) ? i_input_data[888 % IN_WIDTH] : pong_storage_data_337 ^ i_input_data[888 % IN_WIDTH];
                default: pong_storage_data_337 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_337;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_337 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_337;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_337 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_337;
            end
        end
    end
end

logic ping_storage_data_338;
logic pong_storage_data_338;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_338 <= 1'b0;
        pong_storage_data_338 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                85 / IN_WIDTH: ping_storage_data_338 <= (fillup_transition == 1'b1) ? i_input_data[85 % IN_WIDTH] : ping_storage_data_338 ^ i_input_data[85 % IN_WIDTH];
                195 / IN_WIDTH: ping_storage_data_338 <= (fillup_transition == 1'b1) ? i_input_data[195 % IN_WIDTH] : ping_storage_data_338 ^ i_input_data[195 % IN_WIDTH];
                849 / IN_WIDTH: ping_storage_data_338 <= (fillup_transition == 1'b1) ? i_input_data[849 % IN_WIDTH] : ping_storage_data_338 ^ i_input_data[849 % IN_WIDTH];
                889 / IN_WIDTH: ping_storage_data_338 <= (fillup_transition == 1'b1) ? i_input_data[889 % IN_WIDTH] : ping_storage_data_338 ^ i_input_data[889 % IN_WIDTH];
                default: ping_storage_data_338 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_338;
                endcase
            end else begin
                case (input_count)
                85 / IN_WIDTH: pong_storage_data_338 <= (fillup_transition == 1'b1) ? i_input_data[85 % IN_WIDTH] : pong_storage_data_338 ^ i_input_data[85 % IN_WIDTH];
                195 / IN_WIDTH: pong_storage_data_338 <= (fillup_transition == 1'b1) ? i_input_data[195 % IN_WIDTH] : pong_storage_data_338 ^ i_input_data[195 % IN_WIDTH];
                849 / IN_WIDTH: pong_storage_data_338 <= (fillup_transition == 1'b1) ? i_input_data[849 % IN_WIDTH] : pong_storage_data_338 ^ i_input_data[849 % IN_WIDTH];
                889 / IN_WIDTH: pong_storage_data_338 <= (fillup_transition == 1'b1) ? i_input_data[889 % IN_WIDTH] : pong_storage_data_338 ^ i_input_data[889 % IN_WIDTH];
                default: pong_storage_data_338 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_338;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_338 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_338;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_338 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_338;
            end
        end
    end
end

logic ping_storage_data_339;
logic pong_storage_data_339;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_339 <= 1'b0;
        pong_storage_data_339 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                86 / IN_WIDTH: ping_storage_data_339 <= (fillup_transition == 1'b1) ? i_input_data[86 % IN_WIDTH] : ping_storage_data_339 ^ i_input_data[86 % IN_WIDTH];
                196 / IN_WIDTH: ping_storage_data_339 <= (fillup_transition == 1'b1) ? i_input_data[196 % IN_WIDTH] : ping_storage_data_339 ^ i_input_data[196 % IN_WIDTH];
                850 / IN_WIDTH: ping_storage_data_339 <= (fillup_transition == 1'b1) ? i_input_data[850 % IN_WIDTH] : ping_storage_data_339 ^ i_input_data[850 % IN_WIDTH];
                890 / IN_WIDTH: ping_storage_data_339 <= (fillup_transition == 1'b1) ? i_input_data[890 % IN_WIDTH] : ping_storage_data_339 ^ i_input_data[890 % IN_WIDTH];
                default: ping_storage_data_339 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_339;
                endcase
            end else begin
                case (input_count)
                86 / IN_WIDTH: pong_storage_data_339 <= (fillup_transition == 1'b1) ? i_input_data[86 % IN_WIDTH] : pong_storage_data_339 ^ i_input_data[86 % IN_WIDTH];
                196 / IN_WIDTH: pong_storage_data_339 <= (fillup_transition == 1'b1) ? i_input_data[196 % IN_WIDTH] : pong_storage_data_339 ^ i_input_data[196 % IN_WIDTH];
                850 / IN_WIDTH: pong_storage_data_339 <= (fillup_transition == 1'b1) ? i_input_data[850 % IN_WIDTH] : pong_storage_data_339 ^ i_input_data[850 % IN_WIDTH];
                890 / IN_WIDTH: pong_storage_data_339 <= (fillup_transition == 1'b1) ? i_input_data[890 % IN_WIDTH] : pong_storage_data_339 ^ i_input_data[890 % IN_WIDTH];
                default: pong_storage_data_339 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_339;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_339 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_339;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_339 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_339;
            end
        end
    end
end

logic ping_storage_data_340;
logic pong_storage_data_340;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_340 <= 1'b0;
        pong_storage_data_340 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                87 / IN_WIDTH: ping_storage_data_340 <= (fillup_transition == 1'b1) ? i_input_data[87 % IN_WIDTH] : ping_storage_data_340 ^ i_input_data[87 % IN_WIDTH];
                197 / IN_WIDTH: ping_storage_data_340 <= (fillup_transition == 1'b1) ? i_input_data[197 % IN_WIDTH] : ping_storage_data_340 ^ i_input_data[197 % IN_WIDTH];
                851 / IN_WIDTH: ping_storage_data_340 <= (fillup_transition == 1'b1) ? i_input_data[851 % IN_WIDTH] : ping_storage_data_340 ^ i_input_data[851 % IN_WIDTH];
                891 / IN_WIDTH: ping_storage_data_340 <= (fillup_transition == 1'b1) ? i_input_data[891 % IN_WIDTH] : ping_storage_data_340 ^ i_input_data[891 % IN_WIDTH];
                default: ping_storage_data_340 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_340;
                endcase
            end else begin
                case (input_count)
                87 / IN_WIDTH: pong_storage_data_340 <= (fillup_transition == 1'b1) ? i_input_data[87 % IN_WIDTH] : pong_storage_data_340 ^ i_input_data[87 % IN_WIDTH];
                197 / IN_WIDTH: pong_storage_data_340 <= (fillup_transition == 1'b1) ? i_input_data[197 % IN_WIDTH] : pong_storage_data_340 ^ i_input_data[197 % IN_WIDTH];
                851 / IN_WIDTH: pong_storage_data_340 <= (fillup_transition == 1'b1) ? i_input_data[851 % IN_WIDTH] : pong_storage_data_340 ^ i_input_data[851 % IN_WIDTH];
                891 / IN_WIDTH: pong_storage_data_340 <= (fillup_transition == 1'b1) ? i_input_data[891 % IN_WIDTH] : pong_storage_data_340 ^ i_input_data[891 % IN_WIDTH];
                default: pong_storage_data_340 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_340;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_340 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_340;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_340 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_340;
            end
        end
    end
end

logic ping_storage_data_341;
logic pong_storage_data_341;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_341 <= 1'b0;
        pong_storage_data_341 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                88 / IN_WIDTH: ping_storage_data_341 <= (fillup_transition == 1'b1) ? i_input_data[88 % IN_WIDTH] : ping_storage_data_341 ^ i_input_data[88 % IN_WIDTH];
                198 / IN_WIDTH: ping_storage_data_341 <= (fillup_transition == 1'b1) ? i_input_data[198 % IN_WIDTH] : ping_storage_data_341 ^ i_input_data[198 % IN_WIDTH];
                852 / IN_WIDTH: ping_storage_data_341 <= (fillup_transition == 1'b1) ? i_input_data[852 % IN_WIDTH] : ping_storage_data_341 ^ i_input_data[852 % IN_WIDTH];
                892 / IN_WIDTH: ping_storage_data_341 <= (fillup_transition == 1'b1) ? i_input_data[892 % IN_WIDTH] : ping_storage_data_341 ^ i_input_data[892 % IN_WIDTH];
                default: ping_storage_data_341 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_341;
                endcase
            end else begin
                case (input_count)
                88 / IN_WIDTH: pong_storage_data_341 <= (fillup_transition == 1'b1) ? i_input_data[88 % IN_WIDTH] : pong_storage_data_341 ^ i_input_data[88 % IN_WIDTH];
                198 / IN_WIDTH: pong_storage_data_341 <= (fillup_transition == 1'b1) ? i_input_data[198 % IN_WIDTH] : pong_storage_data_341 ^ i_input_data[198 % IN_WIDTH];
                852 / IN_WIDTH: pong_storage_data_341 <= (fillup_transition == 1'b1) ? i_input_data[852 % IN_WIDTH] : pong_storage_data_341 ^ i_input_data[852 % IN_WIDTH];
                892 / IN_WIDTH: pong_storage_data_341 <= (fillup_transition == 1'b1) ? i_input_data[892 % IN_WIDTH] : pong_storage_data_341 ^ i_input_data[892 % IN_WIDTH];
                default: pong_storage_data_341 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_341;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_341 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_341;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_341 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_341;
            end
        end
    end
end

logic ping_storage_data_342;
logic pong_storage_data_342;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_342 <= 1'b0;
        pong_storage_data_342 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                89 / IN_WIDTH: ping_storage_data_342 <= (fillup_transition == 1'b1) ? i_input_data[89 % IN_WIDTH] : ping_storage_data_342 ^ i_input_data[89 % IN_WIDTH];
                199 / IN_WIDTH: ping_storage_data_342 <= (fillup_transition == 1'b1) ? i_input_data[199 % IN_WIDTH] : ping_storage_data_342 ^ i_input_data[199 % IN_WIDTH];
                853 / IN_WIDTH: ping_storage_data_342 <= (fillup_transition == 1'b1) ? i_input_data[853 % IN_WIDTH] : ping_storage_data_342 ^ i_input_data[853 % IN_WIDTH];
                893 / IN_WIDTH: ping_storage_data_342 <= (fillup_transition == 1'b1) ? i_input_data[893 % IN_WIDTH] : ping_storage_data_342 ^ i_input_data[893 % IN_WIDTH];
                default: ping_storage_data_342 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_342;
                endcase
            end else begin
                case (input_count)
                89 / IN_WIDTH: pong_storage_data_342 <= (fillup_transition == 1'b1) ? i_input_data[89 % IN_WIDTH] : pong_storage_data_342 ^ i_input_data[89 % IN_WIDTH];
                199 / IN_WIDTH: pong_storage_data_342 <= (fillup_transition == 1'b1) ? i_input_data[199 % IN_WIDTH] : pong_storage_data_342 ^ i_input_data[199 % IN_WIDTH];
                853 / IN_WIDTH: pong_storage_data_342 <= (fillup_transition == 1'b1) ? i_input_data[853 % IN_WIDTH] : pong_storage_data_342 ^ i_input_data[853 % IN_WIDTH];
                893 / IN_WIDTH: pong_storage_data_342 <= (fillup_transition == 1'b1) ? i_input_data[893 % IN_WIDTH] : pong_storage_data_342 ^ i_input_data[893 % IN_WIDTH];
                default: pong_storage_data_342 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_342;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_342 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_342;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_342 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_342;
            end
        end
    end
end

logic ping_storage_data_343;
logic pong_storage_data_343;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_343 <= 1'b0;
        pong_storage_data_343 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                90 / IN_WIDTH: ping_storage_data_343 <= (fillup_transition == 1'b1) ? i_input_data[90 % IN_WIDTH] : ping_storage_data_343 ^ i_input_data[90 % IN_WIDTH];
                200 / IN_WIDTH: ping_storage_data_343 <= (fillup_transition == 1'b1) ? i_input_data[200 % IN_WIDTH] : ping_storage_data_343 ^ i_input_data[200 % IN_WIDTH];
                854 / IN_WIDTH: ping_storage_data_343 <= (fillup_transition == 1'b1) ? i_input_data[854 % IN_WIDTH] : ping_storage_data_343 ^ i_input_data[854 % IN_WIDTH];
                894 / IN_WIDTH: ping_storage_data_343 <= (fillup_transition == 1'b1) ? i_input_data[894 % IN_WIDTH] : ping_storage_data_343 ^ i_input_data[894 % IN_WIDTH];
                default: ping_storage_data_343 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_343;
                endcase
            end else begin
                case (input_count)
                90 / IN_WIDTH: pong_storage_data_343 <= (fillup_transition == 1'b1) ? i_input_data[90 % IN_WIDTH] : pong_storage_data_343 ^ i_input_data[90 % IN_WIDTH];
                200 / IN_WIDTH: pong_storage_data_343 <= (fillup_transition == 1'b1) ? i_input_data[200 % IN_WIDTH] : pong_storage_data_343 ^ i_input_data[200 % IN_WIDTH];
                854 / IN_WIDTH: pong_storage_data_343 <= (fillup_transition == 1'b1) ? i_input_data[854 % IN_WIDTH] : pong_storage_data_343 ^ i_input_data[854 % IN_WIDTH];
                894 / IN_WIDTH: pong_storage_data_343 <= (fillup_transition == 1'b1) ? i_input_data[894 % IN_WIDTH] : pong_storage_data_343 ^ i_input_data[894 % IN_WIDTH];
                default: pong_storage_data_343 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_343;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_343 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_343;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_343 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_343;
            end
        end
    end
end

logic ping_storage_data_344;
logic pong_storage_data_344;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_344 <= 1'b0;
        pong_storage_data_344 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                91 / IN_WIDTH: ping_storage_data_344 <= (fillup_transition == 1'b1) ? i_input_data[91 % IN_WIDTH] : ping_storage_data_344 ^ i_input_data[91 % IN_WIDTH];
                201 / IN_WIDTH: ping_storage_data_344 <= (fillup_transition == 1'b1) ? i_input_data[201 % IN_WIDTH] : ping_storage_data_344 ^ i_input_data[201 % IN_WIDTH];
                855 / IN_WIDTH: ping_storage_data_344 <= (fillup_transition == 1'b1) ? i_input_data[855 % IN_WIDTH] : ping_storage_data_344 ^ i_input_data[855 % IN_WIDTH];
                895 / IN_WIDTH: ping_storage_data_344 <= (fillup_transition == 1'b1) ? i_input_data[895 % IN_WIDTH] : ping_storage_data_344 ^ i_input_data[895 % IN_WIDTH];
                default: ping_storage_data_344 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_344;
                endcase
            end else begin
                case (input_count)
                91 / IN_WIDTH: pong_storage_data_344 <= (fillup_transition == 1'b1) ? i_input_data[91 % IN_WIDTH] : pong_storage_data_344 ^ i_input_data[91 % IN_WIDTH];
                201 / IN_WIDTH: pong_storage_data_344 <= (fillup_transition == 1'b1) ? i_input_data[201 % IN_WIDTH] : pong_storage_data_344 ^ i_input_data[201 % IN_WIDTH];
                855 / IN_WIDTH: pong_storage_data_344 <= (fillup_transition == 1'b1) ? i_input_data[855 % IN_WIDTH] : pong_storage_data_344 ^ i_input_data[855 % IN_WIDTH];
                895 / IN_WIDTH: pong_storage_data_344 <= (fillup_transition == 1'b1) ? i_input_data[895 % IN_WIDTH] : pong_storage_data_344 ^ i_input_data[895 % IN_WIDTH];
                default: pong_storage_data_344 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_344;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_344 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_344;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_344 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_344;
            end
        end
    end
end

logic ping_storage_data_345;
logic pong_storage_data_345;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_345 <= 1'b0;
        pong_storage_data_345 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                92 / IN_WIDTH: ping_storage_data_345 <= (fillup_transition == 1'b1) ? i_input_data[92 % IN_WIDTH] : ping_storage_data_345 ^ i_input_data[92 % IN_WIDTH];
                202 / IN_WIDTH: ping_storage_data_345 <= (fillup_transition == 1'b1) ? i_input_data[202 % IN_WIDTH] : ping_storage_data_345 ^ i_input_data[202 % IN_WIDTH];
                856 / IN_WIDTH: ping_storage_data_345 <= (fillup_transition == 1'b1) ? i_input_data[856 % IN_WIDTH] : ping_storage_data_345 ^ i_input_data[856 % IN_WIDTH];
                896 / IN_WIDTH: ping_storage_data_345 <= (fillup_transition == 1'b1) ? i_input_data[896 % IN_WIDTH] : ping_storage_data_345 ^ i_input_data[896 % IN_WIDTH];
                default: ping_storage_data_345 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_345;
                endcase
            end else begin
                case (input_count)
                92 / IN_WIDTH: pong_storage_data_345 <= (fillup_transition == 1'b1) ? i_input_data[92 % IN_WIDTH] : pong_storage_data_345 ^ i_input_data[92 % IN_WIDTH];
                202 / IN_WIDTH: pong_storage_data_345 <= (fillup_transition == 1'b1) ? i_input_data[202 % IN_WIDTH] : pong_storage_data_345 ^ i_input_data[202 % IN_WIDTH];
                856 / IN_WIDTH: pong_storage_data_345 <= (fillup_transition == 1'b1) ? i_input_data[856 % IN_WIDTH] : pong_storage_data_345 ^ i_input_data[856 % IN_WIDTH];
                896 / IN_WIDTH: pong_storage_data_345 <= (fillup_transition == 1'b1) ? i_input_data[896 % IN_WIDTH] : pong_storage_data_345 ^ i_input_data[896 % IN_WIDTH];
                default: pong_storage_data_345 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_345;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_345 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_345;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_345 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_345;
            end
        end
    end
end

logic ping_storage_data_346;
logic pong_storage_data_346;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_346 <= 1'b0;
        pong_storage_data_346 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                93 / IN_WIDTH: ping_storage_data_346 <= (fillup_transition == 1'b1) ? i_input_data[93 % IN_WIDTH] : ping_storage_data_346 ^ i_input_data[93 % IN_WIDTH];
                203 / IN_WIDTH: ping_storage_data_346 <= (fillup_transition == 1'b1) ? i_input_data[203 % IN_WIDTH] : ping_storage_data_346 ^ i_input_data[203 % IN_WIDTH];
                857 / IN_WIDTH: ping_storage_data_346 <= (fillup_transition == 1'b1) ? i_input_data[857 % IN_WIDTH] : ping_storage_data_346 ^ i_input_data[857 % IN_WIDTH];
                897 / IN_WIDTH: ping_storage_data_346 <= (fillup_transition == 1'b1) ? i_input_data[897 % IN_WIDTH] : ping_storage_data_346 ^ i_input_data[897 % IN_WIDTH];
                default: ping_storage_data_346 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_346;
                endcase
            end else begin
                case (input_count)
                93 / IN_WIDTH: pong_storage_data_346 <= (fillup_transition == 1'b1) ? i_input_data[93 % IN_WIDTH] : pong_storage_data_346 ^ i_input_data[93 % IN_WIDTH];
                203 / IN_WIDTH: pong_storage_data_346 <= (fillup_transition == 1'b1) ? i_input_data[203 % IN_WIDTH] : pong_storage_data_346 ^ i_input_data[203 % IN_WIDTH];
                857 / IN_WIDTH: pong_storage_data_346 <= (fillup_transition == 1'b1) ? i_input_data[857 % IN_WIDTH] : pong_storage_data_346 ^ i_input_data[857 % IN_WIDTH];
                897 / IN_WIDTH: pong_storage_data_346 <= (fillup_transition == 1'b1) ? i_input_data[897 % IN_WIDTH] : pong_storage_data_346 ^ i_input_data[897 % IN_WIDTH];
                default: pong_storage_data_346 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_346;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_346 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_346;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_346 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_346;
            end
        end
    end
end

logic ping_storage_data_347;
logic pong_storage_data_347;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_347 <= 1'b0;
        pong_storage_data_347 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                94 / IN_WIDTH: ping_storage_data_347 <= (fillup_transition == 1'b1) ? i_input_data[94 % IN_WIDTH] : ping_storage_data_347 ^ i_input_data[94 % IN_WIDTH];
                204 / IN_WIDTH: ping_storage_data_347 <= (fillup_transition == 1'b1) ? i_input_data[204 % IN_WIDTH] : ping_storage_data_347 ^ i_input_data[204 % IN_WIDTH];
                858 / IN_WIDTH: ping_storage_data_347 <= (fillup_transition == 1'b1) ? i_input_data[858 % IN_WIDTH] : ping_storage_data_347 ^ i_input_data[858 % IN_WIDTH];
                898 / IN_WIDTH: ping_storage_data_347 <= (fillup_transition == 1'b1) ? i_input_data[898 % IN_WIDTH] : ping_storage_data_347 ^ i_input_data[898 % IN_WIDTH];
                default: ping_storage_data_347 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_347;
                endcase
            end else begin
                case (input_count)
                94 / IN_WIDTH: pong_storage_data_347 <= (fillup_transition == 1'b1) ? i_input_data[94 % IN_WIDTH] : pong_storage_data_347 ^ i_input_data[94 % IN_WIDTH];
                204 / IN_WIDTH: pong_storage_data_347 <= (fillup_transition == 1'b1) ? i_input_data[204 % IN_WIDTH] : pong_storage_data_347 ^ i_input_data[204 % IN_WIDTH];
                858 / IN_WIDTH: pong_storage_data_347 <= (fillup_transition == 1'b1) ? i_input_data[858 % IN_WIDTH] : pong_storage_data_347 ^ i_input_data[858 % IN_WIDTH];
                898 / IN_WIDTH: pong_storage_data_347 <= (fillup_transition == 1'b1) ? i_input_data[898 % IN_WIDTH] : pong_storage_data_347 ^ i_input_data[898 % IN_WIDTH];
                default: pong_storage_data_347 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_347;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_347 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_347;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_347 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_347;
            end
        end
    end
end

logic ping_storage_data_348;
logic pong_storage_data_348;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_348 <= 1'b0;
        pong_storage_data_348 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                95 / IN_WIDTH: ping_storage_data_348 <= (fillup_transition == 1'b1) ? i_input_data[95 % IN_WIDTH] : ping_storage_data_348 ^ i_input_data[95 % IN_WIDTH];
                205 / IN_WIDTH: ping_storage_data_348 <= (fillup_transition == 1'b1) ? i_input_data[205 % IN_WIDTH] : ping_storage_data_348 ^ i_input_data[205 % IN_WIDTH];
                859 / IN_WIDTH: ping_storage_data_348 <= (fillup_transition == 1'b1) ? i_input_data[859 % IN_WIDTH] : ping_storage_data_348 ^ i_input_data[859 % IN_WIDTH];
                899 / IN_WIDTH: ping_storage_data_348 <= (fillup_transition == 1'b1) ? i_input_data[899 % IN_WIDTH] : ping_storage_data_348 ^ i_input_data[899 % IN_WIDTH];
                default: ping_storage_data_348 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_348;
                endcase
            end else begin
                case (input_count)
                95 / IN_WIDTH: pong_storage_data_348 <= (fillup_transition == 1'b1) ? i_input_data[95 % IN_WIDTH] : pong_storage_data_348 ^ i_input_data[95 % IN_WIDTH];
                205 / IN_WIDTH: pong_storage_data_348 <= (fillup_transition == 1'b1) ? i_input_data[205 % IN_WIDTH] : pong_storage_data_348 ^ i_input_data[205 % IN_WIDTH];
                859 / IN_WIDTH: pong_storage_data_348 <= (fillup_transition == 1'b1) ? i_input_data[859 % IN_WIDTH] : pong_storage_data_348 ^ i_input_data[859 % IN_WIDTH];
                899 / IN_WIDTH: pong_storage_data_348 <= (fillup_transition == 1'b1) ? i_input_data[899 % IN_WIDTH] : pong_storage_data_348 ^ i_input_data[899 % IN_WIDTH];
                default: pong_storage_data_348 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_348;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_348 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_348;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_348 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_348;
            end
        end
    end
end

logic ping_storage_data_349;
logic pong_storage_data_349;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_349 <= 1'b0;
        pong_storage_data_349 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                0 / IN_WIDTH: ping_storage_data_349 <= (fillup_transition == 1'b1) ? i_input_data[0 % IN_WIDTH] : ping_storage_data_349 ^ i_input_data[0 % IN_WIDTH];
                206 / IN_WIDTH: ping_storage_data_349 <= (fillup_transition == 1'b1) ? i_input_data[206 % IN_WIDTH] : ping_storage_data_349 ^ i_input_data[206 % IN_WIDTH];
                860 / IN_WIDTH: ping_storage_data_349 <= (fillup_transition == 1'b1) ? i_input_data[860 % IN_WIDTH] : ping_storage_data_349 ^ i_input_data[860 % IN_WIDTH];
                900 / IN_WIDTH: ping_storage_data_349 <= (fillup_transition == 1'b1) ? i_input_data[900 % IN_WIDTH] : ping_storage_data_349 ^ i_input_data[900 % IN_WIDTH];
                default: ping_storage_data_349 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_349;
                endcase
            end else begin
                case (input_count)
                0 / IN_WIDTH: pong_storage_data_349 <= (fillup_transition == 1'b1) ? i_input_data[0 % IN_WIDTH] : pong_storage_data_349 ^ i_input_data[0 % IN_WIDTH];
                206 / IN_WIDTH: pong_storage_data_349 <= (fillup_transition == 1'b1) ? i_input_data[206 % IN_WIDTH] : pong_storage_data_349 ^ i_input_data[206 % IN_WIDTH];
                860 / IN_WIDTH: pong_storage_data_349 <= (fillup_transition == 1'b1) ? i_input_data[860 % IN_WIDTH] : pong_storage_data_349 ^ i_input_data[860 % IN_WIDTH];
                900 / IN_WIDTH: pong_storage_data_349 <= (fillup_transition == 1'b1) ? i_input_data[900 % IN_WIDTH] : pong_storage_data_349 ^ i_input_data[900 % IN_WIDTH];
                default: pong_storage_data_349 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_349;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_349 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_349;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_349 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_349;
            end
        end
    end
end

logic ping_storage_data_350;
logic pong_storage_data_350;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_350 <= 1'b0;
        pong_storage_data_350 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                1 / IN_WIDTH: ping_storage_data_350 <= (fillup_transition == 1'b1) ? i_input_data[1 % IN_WIDTH] : ping_storage_data_350 ^ i_input_data[1 % IN_WIDTH];
                207 / IN_WIDTH: ping_storage_data_350 <= (fillup_transition == 1'b1) ? i_input_data[207 % IN_WIDTH] : ping_storage_data_350 ^ i_input_data[207 % IN_WIDTH];
                861 / IN_WIDTH: ping_storage_data_350 <= (fillup_transition == 1'b1) ? i_input_data[861 % IN_WIDTH] : ping_storage_data_350 ^ i_input_data[861 % IN_WIDTH];
                901 / IN_WIDTH: ping_storage_data_350 <= (fillup_transition == 1'b1) ? i_input_data[901 % IN_WIDTH] : ping_storage_data_350 ^ i_input_data[901 % IN_WIDTH];
                default: ping_storage_data_350 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_350;
                endcase
            end else begin
                case (input_count)
                1 / IN_WIDTH: pong_storage_data_350 <= (fillup_transition == 1'b1) ? i_input_data[1 % IN_WIDTH] : pong_storage_data_350 ^ i_input_data[1 % IN_WIDTH];
                207 / IN_WIDTH: pong_storage_data_350 <= (fillup_transition == 1'b1) ? i_input_data[207 % IN_WIDTH] : pong_storage_data_350 ^ i_input_data[207 % IN_WIDTH];
                861 / IN_WIDTH: pong_storage_data_350 <= (fillup_transition == 1'b1) ? i_input_data[861 % IN_WIDTH] : pong_storage_data_350 ^ i_input_data[861 % IN_WIDTH];
                901 / IN_WIDTH: pong_storage_data_350 <= (fillup_transition == 1'b1) ? i_input_data[901 % IN_WIDTH] : pong_storage_data_350 ^ i_input_data[901 % IN_WIDTH];
                default: pong_storage_data_350 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_350;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_350 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_350;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_350 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_350;
            end
        end
    end
end

logic ping_storage_data_351;
logic pong_storage_data_351;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_351 <= 1'b0;
        pong_storage_data_351 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                2 / IN_WIDTH: ping_storage_data_351 <= (fillup_transition == 1'b1) ? i_input_data[2 % IN_WIDTH] : ping_storage_data_351 ^ i_input_data[2 % IN_WIDTH];
                208 / IN_WIDTH: ping_storage_data_351 <= (fillup_transition == 1'b1) ? i_input_data[208 % IN_WIDTH] : ping_storage_data_351 ^ i_input_data[208 % IN_WIDTH];
                862 / IN_WIDTH: ping_storage_data_351 <= (fillup_transition == 1'b1) ? i_input_data[862 % IN_WIDTH] : ping_storage_data_351 ^ i_input_data[862 % IN_WIDTH];
                902 / IN_WIDTH: ping_storage_data_351 <= (fillup_transition == 1'b1) ? i_input_data[902 % IN_WIDTH] : ping_storage_data_351 ^ i_input_data[902 % IN_WIDTH];
                default: ping_storage_data_351 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_351;
                endcase
            end else begin
                case (input_count)
                2 / IN_WIDTH: pong_storage_data_351 <= (fillup_transition == 1'b1) ? i_input_data[2 % IN_WIDTH] : pong_storage_data_351 ^ i_input_data[2 % IN_WIDTH];
                208 / IN_WIDTH: pong_storage_data_351 <= (fillup_transition == 1'b1) ? i_input_data[208 % IN_WIDTH] : pong_storage_data_351 ^ i_input_data[208 % IN_WIDTH];
                862 / IN_WIDTH: pong_storage_data_351 <= (fillup_transition == 1'b1) ? i_input_data[862 % IN_WIDTH] : pong_storage_data_351 ^ i_input_data[862 % IN_WIDTH];
                902 / IN_WIDTH: pong_storage_data_351 <= (fillup_transition == 1'b1) ? i_input_data[902 % IN_WIDTH] : pong_storage_data_351 ^ i_input_data[902 % IN_WIDTH];
                default: pong_storage_data_351 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_351;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_351 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_351;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_351 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_351;
            end
        end
    end
end

logic ping_storage_data_352;
logic pong_storage_data_352;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_352 <= 1'b0;
        pong_storage_data_352 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                3 / IN_WIDTH: ping_storage_data_352 <= (fillup_transition == 1'b1) ? i_input_data[3 % IN_WIDTH] : ping_storage_data_352 ^ i_input_data[3 % IN_WIDTH];
                209 / IN_WIDTH: ping_storage_data_352 <= (fillup_transition == 1'b1) ? i_input_data[209 % IN_WIDTH] : ping_storage_data_352 ^ i_input_data[209 % IN_WIDTH];
                863 / IN_WIDTH: ping_storage_data_352 <= (fillup_transition == 1'b1) ? i_input_data[863 % IN_WIDTH] : ping_storage_data_352 ^ i_input_data[863 % IN_WIDTH];
                903 / IN_WIDTH: ping_storage_data_352 <= (fillup_transition == 1'b1) ? i_input_data[903 % IN_WIDTH] : ping_storage_data_352 ^ i_input_data[903 % IN_WIDTH];
                default: ping_storage_data_352 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_352;
                endcase
            end else begin
                case (input_count)
                3 / IN_WIDTH: pong_storage_data_352 <= (fillup_transition == 1'b1) ? i_input_data[3 % IN_WIDTH] : pong_storage_data_352 ^ i_input_data[3 % IN_WIDTH];
                209 / IN_WIDTH: pong_storage_data_352 <= (fillup_transition == 1'b1) ? i_input_data[209 % IN_WIDTH] : pong_storage_data_352 ^ i_input_data[209 % IN_WIDTH];
                863 / IN_WIDTH: pong_storage_data_352 <= (fillup_transition == 1'b1) ? i_input_data[863 % IN_WIDTH] : pong_storage_data_352 ^ i_input_data[863 % IN_WIDTH];
                903 / IN_WIDTH: pong_storage_data_352 <= (fillup_transition == 1'b1) ? i_input_data[903 % IN_WIDTH] : pong_storage_data_352 ^ i_input_data[903 % IN_WIDTH];
                default: pong_storage_data_352 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_352;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_352 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_352;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_352 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_352;
            end
        end
    end
end

logic ping_storage_data_353;
logic pong_storage_data_353;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_353 <= 1'b0;
        pong_storage_data_353 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                4 / IN_WIDTH: ping_storage_data_353 <= (fillup_transition == 1'b1) ? i_input_data[4 % IN_WIDTH] : ping_storage_data_353 ^ i_input_data[4 % IN_WIDTH];
                210 / IN_WIDTH: ping_storage_data_353 <= (fillup_transition == 1'b1) ? i_input_data[210 % IN_WIDTH] : ping_storage_data_353 ^ i_input_data[210 % IN_WIDTH];
                768 / IN_WIDTH: ping_storage_data_353 <= (fillup_transition == 1'b1) ? i_input_data[768 % IN_WIDTH] : ping_storage_data_353 ^ i_input_data[768 % IN_WIDTH];
                904 / IN_WIDTH: ping_storage_data_353 <= (fillup_transition == 1'b1) ? i_input_data[904 % IN_WIDTH] : ping_storage_data_353 ^ i_input_data[904 % IN_WIDTH];
                default: ping_storage_data_353 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_353;
                endcase
            end else begin
                case (input_count)
                4 / IN_WIDTH: pong_storage_data_353 <= (fillup_transition == 1'b1) ? i_input_data[4 % IN_WIDTH] : pong_storage_data_353 ^ i_input_data[4 % IN_WIDTH];
                210 / IN_WIDTH: pong_storage_data_353 <= (fillup_transition == 1'b1) ? i_input_data[210 % IN_WIDTH] : pong_storage_data_353 ^ i_input_data[210 % IN_WIDTH];
                768 / IN_WIDTH: pong_storage_data_353 <= (fillup_transition == 1'b1) ? i_input_data[768 % IN_WIDTH] : pong_storage_data_353 ^ i_input_data[768 % IN_WIDTH];
                904 / IN_WIDTH: pong_storage_data_353 <= (fillup_transition == 1'b1) ? i_input_data[904 % IN_WIDTH] : pong_storage_data_353 ^ i_input_data[904 % IN_WIDTH];
                default: pong_storage_data_353 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_353;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_353 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_353;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_353 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_353;
            end
        end
    end
end

logic ping_storage_data_354;
logic pong_storage_data_354;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_354 <= 1'b0;
        pong_storage_data_354 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                5 / IN_WIDTH: ping_storage_data_354 <= (fillup_transition == 1'b1) ? i_input_data[5 % IN_WIDTH] : ping_storage_data_354 ^ i_input_data[5 % IN_WIDTH];
                211 / IN_WIDTH: ping_storage_data_354 <= (fillup_transition == 1'b1) ? i_input_data[211 % IN_WIDTH] : ping_storage_data_354 ^ i_input_data[211 % IN_WIDTH];
                769 / IN_WIDTH: ping_storage_data_354 <= (fillup_transition == 1'b1) ? i_input_data[769 % IN_WIDTH] : ping_storage_data_354 ^ i_input_data[769 % IN_WIDTH];
                905 / IN_WIDTH: ping_storage_data_354 <= (fillup_transition == 1'b1) ? i_input_data[905 % IN_WIDTH] : ping_storage_data_354 ^ i_input_data[905 % IN_WIDTH];
                default: ping_storage_data_354 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_354;
                endcase
            end else begin
                case (input_count)
                5 / IN_WIDTH: pong_storage_data_354 <= (fillup_transition == 1'b1) ? i_input_data[5 % IN_WIDTH] : pong_storage_data_354 ^ i_input_data[5 % IN_WIDTH];
                211 / IN_WIDTH: pong_storage_data_354 <= (fillup_transition == 1'b1) ? i_input_data[211 % IN_WIDTH] : pong_storage_data_354 ^ i_input_data[211 % IN_WIDTH];
                769 / IN_WIDTH: pong_storage_data_354 <= (fillup_transition == 1'b1) ? i_input_data[769 % IN_WIDTH] : pong_storage_data_354 ^ i_input_data[769 % IN_WIDTH];
                905 / IN_WIDTH: pong_storage_data_354 <= (fillup_transition == 1'b1) ? i_input_data[905 % IN_WIDTH] : pong_storage_data_354 ^ i_input_data[905 % IN_WIDTH];
                default: pong_storage_data_354 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_354;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_354 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_354;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_354 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_354;
            end
        end
    end
end

logic ping_storage_data_355;
logic pong_storage_data_355;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_355 <= 1'b0;
        pong_storage_data_355 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                6 / IN_WIDTH: ping_storage_data_355 <= (fillup_transition == 1'b1) ? i_input_data[6 % IN_WIDTH] : ping_storage_data_355 ^ i_input_data[6 % IN_WIDTH];
                212 / IN_WIDTH: ping_storage_data_355 <= (fillup_transition == 1'b1) ? i_input_data[212 % IN_WIDTH] : ping_storage_data_355 ^ i_input_data[212 % IN_WIDTH];
                770 / IN_WIDTH: ping_storage_data_355 <= (fillup_transition == 1'b1) ? i_input_data[770 % IN_WIDTH] : ping_storage_data_355 ^ i_input_data[770 % IN_WIDTH];
                906 / IN_WIDTH: ping_storage_data_355 <= (fillup_transition == 1'b1) ? i_input_data[906 % IN_WIDTH] : ping_storage_data_355 ^ i_input_data[906 % IN_WIDTH];
                default: ping_storage_data_355 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_355;
                endcase
            end else begin
                case (input_count)
                6 / IN_WIDTH: pong_storage_data_355 <= (fillup_transition == 1'b1) ? i_input_data[6 % IN_WIDTH] : pong_storage_data_355 ^ i_input_data[6 % IN_WIDTH];
                212 / IN_WIDTH: pong_storage_data_355 <= (fillup_transition == 1'b1) ? i_input_data[212 % IN_WIDTH] : pong_storage_data_355 ^ i_input_data[212 % IN_WIDTH];
                770 / IN_WIDTH: pong_storage_data_355 <= (fillup_transition == 1'b1) ? i_input_data[770 % IN_WIDTH] : pong_storage_data_355 ^ i_input_data[770 % IN_WIDTH];
                906 / IN_WIDTH: pong_storage_data_355 <= (fillup_transition == 1'b1) ? i_input_data[906 % IN_WIDTH] : pong_storage_data_355 ^ i_input_data[906 % IN_WIDTH];
                default: pong_storage_data_355 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_355;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_355 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_355;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_355 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_355;
            end
        end
    end
end

logic ping_storage_data_356;
logic pong_storage_data_356;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_356 <= 1'b0;
        pong_storage_data_356 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                7 / IN_WIDTH: ping_storage_data_356 <= (fillup_transition == 1'b1) ? i_input_data[7 % IN_WIDTH] : ping_storage_data_356 ^ i_input_data[7 % IN_WIDTH];
                213 / IN_WIDTH: ping_storage_data_356 <= (fillup_transition == 1'b1) ? i_input_data[213 % IN_WIDTH] : ping_storage_data_356 ^ i_input_data[213 % IN_WIDTH];
                771 / IN_WIDTH: ping_storage_data_356 <= (fillup_transition == 1'b1) ? i_input_data[771 % IN_WIDTH] : ping_storage_data_356 ^ i_input_data[771 % IN_WIDTH];
                907 / IN_WIDTH: ping_storage_data_356 <= (fillup_transition == 1'b1) ? i_input_data[907 % IN_WIDTH] : ping_storage_data_356 ^ i_input_data[907 % IN_WIDTH];
                default: ping_storage_data_356 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_356;
                endcase
            end else begin
                case (input_count)
                7 / IN_WIDTH: pong_storage_data_356 <= (fillup_transition == 1'b1) ? i_input_data[7 % IN_WIDTH] : pong_storage_data_356 ^ i_input_data[7 % IN_WIDTH];
                213 / IN_WIDTH: pong_storage_data_356 <= (fillup_transition == 1'b1) ? i_input_data[213 % IN_WIDTH] : pong_storage_data_356 ^ i_input_data[213 % IN_WIDTH];
                771 / IN_WIDTH: pong_storage_data_356 <= (fillup_transition == 1'b1) ? i_input_data[771 % IN_WIDTH] : pong_storage_data_356 ^ i_input_data[771 % IN_WIDTH];
                907 / IN_WIDTH: pong_storage_data_356 <= (fillup_transition == 1'b1) ? i_input_data[907 % IN_WIDTH] : pong_storage_data_356 ^ i_input_data[907 % IN_WIDTH];
                default: pong_storage_data_356 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_356;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_356 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_356;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_356 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_356;
            end
        end
    end
end

logic ping_storage_data_357;
logic pong_storage_data_357;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_357 <= 1'b0;
        pong_storage_data_357 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                8 / IN_WIDTH: ping_storage_data_357 <= (fillup_transition == 1'b1) ? i_input_data[8 % IN_WIDTH] : ping_storage_data_357 ^ i_input_data[8 % IN_WIDTH];
                214 / IN_WIDTH: ping_storage_data_357 <= (fillup_transition == 1'b1) ? i_input_data[214 % IN_WIDTH] : ping_storage_data_357 ^ i_input_data[214 % IN_WIDTH];
                772 / IN_WIDTH: ping_storage_data_357 <= (fillup_transition == 1'b1) ? i_input_data[772 % IN_WIDTH] : ping_storage_data_357 ^ i_input_data[772 % IN_WIDTH];
                908 / IN_WIDTH: ping_storage_data_357 <= (fillup_transition == 1'b1) ? i_input_data[908 % IN_WIDTH] : ping_storage_data_357 ^ i_input_data[908 % IN_WIDTH];
                default: ping_storage_data_357 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_357;
                endcase
            end else begin
                case (input_count)
                8 / IN_WIDTH: pong_storage_data_357 <= (fillup_transition == 1'b1) ? i_input_data[8 % IN_WIDTH] : pong_storage_data_357 ^ i_input_data[8 % IN_WIDTH];
                214 / IN_WIDTH: pong_storage_data_357 <= (fillup_transition == 1'b1) ? i_input_data[214 % IN_WIDTH] : pong_storage_data_357 ^ i_input_data[214 % IN_WIDTH];
                772 / IN_WIDTH: pong_storage_data_357 <= (fillup_transition == 1'b1) ? i_input_data[772 % IN_WIDTH] : pong_storage_data_357 ^ i_input_data[772 % IN_WIDTH];
                908 / IN_WIDTH: pong_storage_data_357 <= (fillup_transition == 1'b1) ? i_input_data[908 % IN_WIDTH] : pong_storage_data_357 ^ i_input_data[908 % IN_WIDTH];
                default: pong_storage_data_357 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_357;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_357 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_357;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_357 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_357;
            end
        end
    end
end

logic ping_storage_data_358;
logic pong_storage_data_358;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_358 <= 1'b0;
        pong_storage_data_358 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                9 / IN_WIDTH: ping_storage_data_358 <= (fillup_transition == 1'b1) ? i_input_data[9 % IN_WIDTH] : ping_storage_data_358 ^ i_input_data[9 % IN_WIDTH];
                215 / IN_WIDTH: ping_storage_data_358 <= (fillup_transition == 1'b1) ? i_input_data[215 % IN_WIDTH] : ping_storage_data_358 ^ i_input_data[215 % IN_WIDTH];
                773 / IN_WIDTH: ping_storage_data_358 <= (fillup_transition == 1'b1) ? i_input_data[773 % IN_WIDTH] : ping_storage_data_358 ^ i_input_data[773 % IN_WIDTH];
                909 / IN_WIDTH: ping_storage_data_358 <= (fillup_transition == 1'b1) ? i_input_data[909 % IN_WIDTH] : ping_storage_data_358 ^ i_input_data[909 % IN_WIDTH];
                default: ping_storage_data_358 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_358;
                endcase
            end else begin
                case (input_count)
                9 / IN_WIDTH: pong_storage_data_358 <= (fillup_transition == 1'b1) ? i_input_data[9 % IN_WIDTH] : pong_storage_data_358 ^ i_input_data[9 % IN_WIDTH];
                215 / IN_WIDTH: pong_storage_data_358 <= (fillup_transition == 1'b1) ? i_input_data[215 % IN_WIDTH] : pong_storage_data_358 ^ i_input_data[215 % IN_WIDTH];
                773 / IN_WIDTH: pong_storage_data_358 <= (fillup_transition == 1'b1) ? i_input_data[773 % IN_WIDTH] : pong_storage_data_358 ^ i_input_data[773 % IN_WIDTH];
                909 / IN_WIDTH: pong_storage_data_358 <= (fillup_transition == 1'b1) ? i_input_data[909 % IN_WIDTH] : pong_storage_data_358 ^ i_input_data[909 % IN_WIDTH];
                default: pong_storage_data_358 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_358;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_358 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_358;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_358 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_358;
            end
        end
    end
end

logic ping_storage_data_359;
logic pong_storage_data_359;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_359 <= 1'b0;
        pong_storage_data_359 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                10 / IN_WIDTH: ping_storage_data_359 <= (fillup_transition == 1'b1) ? i_input_data[10 % IN_WIDTH] : ping_storage_data_359 ^ i_input_data[10 % IN_WIDTH];
                216 / IN_WIDTH: ping_storage_data_359 <= (fillup_transition == 1'b1) ? i_input_data[216 % IN_WIDTH] : ping_storage_data_359 ^ i_input_data[216 % IN_WIDTH];
                774 / IN_WIDTH: ping_storage_data_359 <= (fillup_transition == 1'b1) ? i_input_data[774 % IN_WIDTH] : ping_storage_data_359 ^ i_input_data[774 % IN_WIDTH];
                910 / IN_WIDTH: ping_storage_data_359 <= (fillup_transition == 1'b1) ? i_input_data[910 % IN_WIDTH] : ping_storage_data_359 ^ i_input_data[910 % IN_WIDTH];
                default: ping_storage_data_359 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_359;
                endcase
            end else begin
                case (input_count)
                10 / IN_WIDTH: pong_storage_data_359 <= (fillup_transition == 1'b1) ? i_input_data[10 % IN_WIDTH] : pong_storage_data_359 ^ i_input_data[10 % IN_WIDTH];
                216 / IN_WIDTH: pong_storage_data_359 <= (fillup_transition == 1'b1) ? i_input_data[216 % IN_WIDTH] : pong_storage_data_359 ^ i_input_data[216 % IN_WIDTH];
                774 / IN_WIDTH: pong_storage_data_359 <= (fillup_transition == 1'b1) ? i_input_data[774 % IN_WIDTH] : pong_storage_data_359 ^ i_input_data[774 % IN_WIDTH];
                910 / IN_WIDTH: pong_storage_data_359 <= (fillup_transition == 1'b1) ? i_input_data[910 % IN_WIDTH] : pong_storage_data_359 ^ i_input_data[910 % IN_WIDTH];
                default: pong_storage_data_359 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_359;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_359 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_359;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_359 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_359;
            end
        end
    end
end

logic ping_storage_data_360;
logic pong_storage_data_360;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_360 <= 1'b0;
        pong_storage_data_360 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                11 / IN_WIDTH: ping_storage_data_360 <= (fillup_transition == 1'b1) ? i_input_data[11 % IN_WIDTH] : ping_storage_data_360 ^ i_input_data[11 % IN_WIDTH];
                217 / IN_WIDTH: ping_storage_data_360 <= (fillup_transition == 1'b1) ? i_input_data[217 % IN_WIDTH] : ping_storage_data_360 ^ i_input_data[217 % IN_WIDTH];
                775 / IN_WIDTH: ping_storage_data_360 <= (fillup_transition == 1'b1) ? i_input_data[775 % IN_WIDTH] : ping_storage_data_360 ^ i_input_data[775 % IN_WIDTH];
                911 / IN_WIDTH: ping_storage_data_360 <= (fillup_transition == 1'b1) ? i_input_data[911 % IN_WIDTH] : ping_storage_data_360 ^ i_input_data[911 % IN_WIDTH];
                default: ping_storage_data_360 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_360;
                endcase
            end else begin
                case (input_count)
                11 / IN_WIDTH: pong_storage_data_360 <= (fillup_transition == 1'b1) ? i_input_data[11 % IN_WIDTH] : pong_storage_data_360 ^ i_input_data[11 % IN_WIDTH];
                217 / IN_WIDTH: pong_storage_data_360 <= (fillup_transition == 1'b1) ? i_input_data[217 % IN_WIDTH] : pong_storage_data_360 ^ i_input_data[217 % IN_WIDTH];
                775 / IN_WIDTH: pong_storage_data_360 <= (fillup_transition == 1'b1) ? i_input_data[775 % IN_WIDTH] : pong_storage_data_360 ^ i_input_data[775 % IN_WIDTH];
                911 / IN_WIDTH: pong_storage_data_360 <= (fillup_transition == 1'b1) ? i_input_data[911 % IN_WIDTH] : pong_storage_data_360 ^ i_input_data[911 % IN_WIDTH];
                default: pong_storage_data_360 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_360;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_360 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_360;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_360 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_360;
            end
        end
    end
end

logic ping_storage_data_361;
logic pong_storage_data_361;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_361 <= 1'b0;
        pong_storage_data_361 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                12 / IN_WIDTH: ping_storage_data_361 <= (fillup_transition == 1'b1) ? i_input_data[12 % IN_WIDTH] : ping_storage_data_361 ^ i_input_data[12 % IN_WIDTH];
                218 / IN_WIDTH: ping_storage_data_361 <= (fillup_transition == 1'b1) ? i_input_data[218 % IN_WIDTH] : ping_storage_data_361 ^ i_input_data[218 % IN_WIDTH];
                776 / IN_WIDTH: ping_storage_data_361 <= (fillup_transition == 1'b1) ? i_input_data[776 % IN_WIDTH] : ping_storage_data_361 ^ i_input_data[776 % IN_WIDTH];
                912 / IN_WIDTH: ping_storage_data_361 <= (fillup_transition == 1'b1) ? i_input_data[912 % IN_WIDTH] : ping_storage_data_361 ^ i_input_data[912 % IN_WIDTH];
                default: ping_storage_data_361 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_361;
                endcase
            end else begin
                case (input_count)
                12 / IN_WIDTH: pong_storage_data_361 <= (fillup_transition == 1'b1) ? i_input_data[12 % IN_WIDTH] : pong_storage_data_361 ^ i_input_data[12 % IN_WIDTH];
                218 / IN_WIDTH: pong_storage_data_361 <= (fillup_transition == 1'b1) ? i_input_data[218 % IN_WIDTH] : pong_storage_data_361 ^ i_input_data[218 % IN_WIDTH];
                776 / IN_WIDTH: pong_storage_data_361 <= (fillup_transition == 1'b1) ? i_input_data[776 % IN_WIDTH] : pong_storage_data_361 ^ i_input_data[776 % IN_WIDTH];
                912 / IN_WIDTH: pong_storage_data_361 <= (fillup_transition == 1'b1) ? i_input_data[912 % IN_WIDTH] : pong_storage_data_361 ^ i_input_data[912 % IN_WIDTH];
                default: pong_storage_data_361 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_361;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_361 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_361;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_361 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_361;
            end
        end
    end
end

logic ping_storage_data_362;
logic pong_storage_data_362;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_362 <= 1'b0;
        pong_storage_data_362 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                13 / IN_WIDTH: ping_storage_data_362 <= (fillup_transition == 1'b1) ? i_input_data[13 % IN_WIDTH] : ping_storage_data_362 ^ i_input_data[13 % IN_WIDTH];
                219 / IN_WIDTH: ping_storage_data_362 <= (fillup_transition == 1'b1) ? i_input_data[219 % IN_WIDTH] : ping_storage_data_362 ^ i_input_data[219 % IN_WIDTH];
                777 / IN_WIDTH: ping_storage_data_362 <= (fillup_transition == 1'b1) ? i_input_data[777 % IN_WIDTH] : ping_storage_data_362 ^ i_input_data[777 % IN_WIDTH];
                913 / IN_WIDTH: ping_storage_data_362 <= (fillup_transition == 1'b1) ? i_input_data[913 % IN_WIDTH] : ping_storage_data_362 ^ i_input_data[913 % IN_WIDTH];
                default: ping_storage_data_362 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_362;
                endcase
            end else begin
                case (input_count)
                13 / IN_WIDTH: pong_storage_data_362 <= (fillup_transition == 1'b1) ? i_input_data[13 % IN_WIDTH] : pong_storage_data_362 ^ i_input_data[13 % IN_WIDTH];
                219 / IN_WIDTH: pong_storage_data_362 <= (fillup_transition == 1'b1) ? i_input_data[219 % IN_WIDTH] : pong_storage_data_362 ^ i_input_data[219 % IN_WIDTH];
                777 / IN_WIDTH: pong_storage_data_362 <= (fillup_transition == 1'b1) ? i_input_data[777 % IN_WIDTH] : pong_storage_data_362 ^ i_input_data[777 % IN_WIDTH];
                913 / IN_WIDTH: pong_storage_data_362 <= (fillup_transition == 1'b1) ? i_input_data[913 % IN_WIDTH] : pong_storage_data_362 ^ i_input_data[913 % IN_WIDTH];
                default: pong_storage_data_362 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_362;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_362 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_362;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_362 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_362;
            end
        end
    end
end

logic ping_storage_data_363;
logic pong_storage_data_363;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_363 <= 1'b0;
        pong_storage_data_363 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                14 / IN_WIDTH: ping_storage_data_363 <= (fillup_transition == 1'b1) ? i_input_data[14 % IN_WIDTH] : ping_storage_data_363 ^ i_input_data[14 % IN_WIDTH];
                220 / IN_WIDTH: ping_storage_data_363 <= (fillup_transition == 1'b1) ? i_input_data[220 % IN_WIDTH] : ping_storage_data_363 ^ i_input_data[220 % IN_WIDTH];
                778 / IN_WIDTH: ping_storage_data_363 <= (fillup_transition == 1'b1) ? i_input_data[778 % IN_WIDTH] : ping_storage_data_363 ^ i_input_data[778 % IN_WIDTH];
                914 / IN_WIDTH: ping_storage_data_363 <= (fillup_transition == 1'b1) ? i_input_data[914 % IN_WIDTH] : ping_storage_data_363 ^ i_input_data[914 % IN_WIDTH];
                default: ping_storage_data_363 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_363;
                endcase
            end else begin
                case (input_count)
                14 / IN_WIDTH: pong_storage_data_363 <= (fillup_transition == 1'b1) ? i_input_data[14 % IN_WIDTH] : pong_storage_data_363 ^ i_input_data[14 % IN_WIDTH];
                220 / IN_WIDTH: pong_storage_data_363 <= (fillup_transition == 1'b1) ? i_input_data[220 % IN_WIDTH] : pong_storage_data_363 ^ i_input_data[220 % IN_WIDTH];
                778 / IN_WIDTH: pong_storage_data_363 <= (fillup_transition == 1'b1) ? i_input_data[778 % IN_WIDTH] : pong_storage_data_363 ^ i_input_data[778 % IN_WIDTH];
                914 / IN_WIDTH: pong_storage_data_363 <= (fillup_transition == 1'b1) ? i_input_data[914 % IN_WIDTH] : pong_storage_data_363 ^ i_input_data[914 % IN_WIDTH];
                default: pong_storage_data_363 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_363;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_363 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_363;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_363 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_363;
            end
        end
    end
end

logic ping_storage_data_364;
logic pong_storage_data_364;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_364 <= 1'b0;
        pong_storage_data_364 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                15 / IN_WIDTH: ping_storage_data_364 <= (fillup_transition == 1'b1) ? i_input_data[15 % IN_WIDTH] : ping_storage_data_364 ^ i_input_data[15 % IN_WIDTH];
                221 / IN_WIDTH: ping_storage_data_364 <= (fillup_transition == 1'b1) ? i_input_data[221 % IN_WIDTH] : ping_storage_data_364 ^ i_input_data[221 % IN_WIDTH];
                779 / IN_WIDTH: ping_storage_data_364 <= (fillup_transition == 1'b1) ? i_input_data[779 % IN_WIDTH] : ping_storage_data_364 ^ i_input_data[779 % IN_WIDTH];
                915 / IN_WIDTH: ping_storage_data_364 <= (fillup_transition == 1'b1) ? i_input_data[915 % IN_WIDTH] : ping_storage_data_364 ^ i_input_data[915 % IN_WIDTH];
                default: ping_storage_data_364 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_364;
                endcase
            end else begin
                case (input_count)
                15 / IN_WIDTH: pong_storage_data_364 <= (fillup_transition == 1'b1) ? i_input_data[15 % IN_WIDTH] : pong_storage_data_364 ^ i_input_data[15 % IN_WIDTH];
                221 / IN_WIDTH: pong_storage_data_364 <= (fillup_transition == 1'b1) ? i_input_data[221 % IN_WIDTH] : pong_storage_data_364 ^ i_input_data[221 % IN_WIDTH];
                779 / IN_WIDTH: pong_storage_data_364 <= (fillup_transition == 1'b1) ? i_input_data[779 % IN_WIDTH] : pong_storage_data_364 ^ i_input_data[779 % IN_WIDTH];
                915 / IN_WIDTH: pong_storage_data_364 <= (fillup_transition == 1'b1) ? i_input_data[915 % IN_WIDTH] : pong_storage_data_364 ^ i_input_data[915 % IN_WIDTH];
                default: pong_storage_data_364 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_364;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_364 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_364;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_364 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_364;
            end
        end
    end
end

logic ping_storage_data_365;
logic pong_storage_data_365;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_365 <= 1'b0;
        pong_storage_data_365 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                16 / IN_WIDTH: ping_storage_data_365 <= (fillup_transition == 1'b1) ? i_input_data[16 % IN_WIDTH] : ping_storage_data_365 ^ i_input_data[16 % IN_WIDTH];
                222 / IN_WIDTH: ping_storage_data_365 <= (fillup_transition == 1'b1) ? i_input_data[222 % IN_WIDTH] : ping_storage_data_365 ^ i_input_data[222 % IN_WIDTH];
                780 / IN_WIDTH: ping_storage_data_365 <= (fillup_transition == 1'b1) ? i_input_data[780 % IN_WIDTH] : ping_storage_data_365 ^ i_input_data[780 % IN_WIDTH];
                916 / IN_WIDTH: ping_storage_data_365 <= (fillup_transition == 1'b1) ? i_input_data[916 % IN_WIDTH] : ping_storage_data_365 ^ i_input_data[916 % IN_WIDTH];
                default: ping_storage_data_365 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_365;
                endcase
            end else begin
                case (input_count)
                16 / IN_WIDTH: pong_storage_data_365 <= (fillup_transition == 1'b1) ? i_input_data[16 % IN_WIDTH] : pong_storage_data_365 ^ i_input_data[16 % IN_WIDTH];
                222 / IN_WIDTH: pong_storage_data_365 <= (fillup_transition == 1'b1) ? i_input_data[222 % IN_WIDTH] : pong_storage_data_365 ^ i_input_data[222 % IN_WIDTH];
                780 / IN_WIDTH: pong_storage_data_365 <= (fillup_transition == 1'b1) ? i_input_data[780 % IN_WIDTH] : pong_storage_data_365 ^ i_input_data[780 % IN_WIDTH];
                916 / IN_WIDTH: pong_storage_data_365 <= (fillup_transition == 1'b1) ? i_input_data[916 % IN_WIDTH] : pong_storage_data_365 ^ i_input_data[916 % IN_WIDTH];
                default: pong_storage_data_365 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_365;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_365 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_365;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_365 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_365;
            end
        end
    end
end

logic ping_storage_data_366;
logic pong_storage_data_366;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_366 <= 1'b0;
        pong_storage_data_366 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                17 / IN_WIDTH: ping_storage_data_366 <= (fillup_transition == 1'b1) ? i_input_data[17 % IN_WIDTH] : ping_storage_data_366 ^ i_input_data[17 % IN_WIDTH];
                223 / IN_WIDTH: ping_storage_data_366 <= (fillup_transition == 1'b1) ? i_input_data[223 % IN_WIDTH] : ping_storage_data_366 ^ i_input_data[223 % IN_WIDTH];
                781 / IN_WIDTH: ping_storage_data_366 <= (fillup_transition == 1'b1) ? i_input_data[781 % IN_WIDTH] : ping_storage_data_366 ^ i_input_data[781 % IN_WIDTH];
                917 / IN_WIDTH: ping_storage_data_366 <= (fillup_transition == 1'b1) ? i_input_data[917 % IN_WIDTH] : ping_storage_data_366 ^ i_input_data[917 % IN_WIDTH];
                default: ping_storage_data_366 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_366;
                endcase
            end else begin
                case (input_count)
                17 / IN_WIDTH: pong_storage_data_366 <= (fillup_transition == 1'b1) ? i_input_data[17 % IN_WIDTH] : pong_storage_data_366 ^ i_input_data[17 % IN_WIDTH];
                223 / IN_WIDTH: pong_storage_data_366 <= (fillup_transition == 1'b1) ? i_input_data[223 % IN_WIDTH] : pong_storage_data_366 ^ i_input_data[223 % IN_WIDTH];
                781 / IN_WIDTH: pong_storage_data_366 <= (fillup_transition == 1'b1) ? i_input_data[781 % IN_WIDTH] : pong_storage_data_366 ^ i_input_data[781 % IN_WIDTH];
                917 / IN_WIDTH: pong_storage_data_366 <= (fillup_transition == 1'b1) ? i_input_data[917 % IN_WIDTH] : pong_storage_data_366 ^ i_input_data[917 % IN_WIDTH];
                default: pong_storage_data_366 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_366;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_366 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_366;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_366 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_366;
            end
        end
    end
end

logic ping_storage_data_367;
logic pong_storage_data_367;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_367 <= 1'b0;
        pong_storage_data_367 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                18 / IN_WIDTH: ping_storage_data_367 <= (fillup_transition == 1'b1) ? i_input_data[18 % IN_WIDTH] : ping_storage_data_367 ^ i_input_data[18 % IN_WIDTH];
                224 / IN_WIDTH: ping_storage_data_367 <= (fillup_transition == 1'b1) ? i_input_data[224 % IN_WIDTH] : ping_storage_data_367 ^ i_input_data[224 % IN_WIDTH];
                782 / IN_WIDTH: ping_storage_data_367 <= (fillup_transition == 1'b1) ? i_input_data[782 % IN_WIDTH] : ping_storage_data_367 ^ i_input_data[782 % IN_WIDTH];
                918 / IN_WIDTH: ping_storage_data_367 <= (fillup_transition == 1'b1) ? i_input_data[918 % IN_WIDTH] : ping_storage_data_367 ^ i_input_data[918 % IN_WIDTH];
                default: ping_storage_data_367 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_367;
                endcase
            end else begin
                case (input_count)
                18 / IN_WIDTH: pong_storage_data_367 <= (fillup_transition == 1'b1) ? i_input_data[18 % IN_WIDTH] : pong_storage_data_367 ^ i_input_data[18 % IN_WIDTH];
                224 / IN_WIDTH: pong_storage_data_367 <= (fillup_transition == 1'b1) ? i_input_data[224 % IN_WIDTH] : pong_storage_data_367 ^ i_input_data[224 % IN_WIDTH];
                782 / IN_WIDTH: pong_storage_data_367 <= (fillup_transition == 1'b1) ? i_input_data[782 % IN_WIDTH] : pong_storage_data_367 ^ i_input_data[782 % IN_WIDTH];
                918 / IN_WIDTH: pong_storage_data_367 <= (fillup_transition == 1'b1) ? i_input_data[918 % IN_WIDTH] : pong_storage_data_367 ^ i_input_data[918 % IN_WIDTH];
                default: pong_storage_data_367 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_367;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_367 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_367;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_367 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_367;
            end
        end
    end
end

logic ping_storage_data_368;
logic pong_storage_data_368;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_368 <= 1'b0;
        pong_storage_data_368 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                19 / IN_WIDTH: ping_storage_data_368 <= (fillup_transition == 1'b1) ? i_input_data[19 % IN_WIDTH] : ping_storage_data_368 ^ i_input_data[19 % IN_WIDTH];
                225 / IN_WIDTH: ping_storage_data_368 <= (fillup_transition == 1'b1) ? i_input_data[225 % IN_WIDTH] : ping_storage_data_368 ^ i_input_data[225 % IN_WIDTH];
                783 / IN_WIDTH: ping_storage_data_368 <= (fillup_transition == 1'b1) ? i_input_data[783 % IN_WIDTH] : ping_storage_data_368 ^ i_input_data[783 % IN_WIDTH];
                919 / IN_WIDTH: ping_storage_data_368 <= (fillup_transition == 1'b1) ? i_input_data[919 % IN_WIDTH] : ping_storage_data_368 ^ i_input_data[919 % IN_WIDTH];
                default: ping_storage_data_368 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_368;
                endcase
            end else begin
                case (input_count)
                19 / IN_WIDTH: pong_storage_data_368 <= (fillup_transition == 1'b1) ? i_input_data[19 % IN_WIDTH] : pong_storage_data_368 ^ i_input_data[19 % IN_WIDTH];
                225 / IN_WIDTH: pong_storage_data_368 <= (fillup_transition == 1'b1) ? i_input_data[225 % IN_WIDTH] : pong_storage_data_368 ^ i_input_data[225 % IN_WIDTH];
                783 / IN_WIDTH: pong_storage_data_368 <= (fillup_transition == 1'b1) ? i_input_data[783 % IN_WIDTH] : pong_storage_data_368 ^ i_input_data[783 % IN_WIDTH];
                919 / IN_WIDTH: pong_storage_data_368 <= (fillup_transition == 1'b1) ? i_input_data[919 % IN_WIDTH] : pong_storage_data_368 ^ i_input_data[919 % IN_WIDTH];
                default: pong_storage_data_368 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_368;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_368 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_368;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_368 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_368;
            end
        end
    end
end

logic ping_storage_data_369;
logic pong_storage_data_369;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_369 <= 1'b0;
        pong_storage_data_369 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                20 / IN_WIDTH: ping_storage_data_369 <= (fillup_transition == 1'b1) ? i_input_data[20 % IN_WIDTH] : ping_storage_data_369 ^ i_input_data[20 % IN_WIDTH];
                226 / IN_WIDTH: ping_storage_data_369 <= (fillup_transition == 1'b1) ? i_input_data[226 % IN_WIDTH] : ping_storage_data_369 ^ i_input_data[226 % IN_WIDTH];
                784 / IN_WIDTH: ping_storage_data_369 <= (fillup_transition == 1'b1) ? i_input_data[784 % IN_WIDTH] : ping_storage_data_369 ^ i_input_data[784 % IN_WIDTH];
                920 / IN_WIDTH: ping_storage_data_369 <= (fillup_transition == 1'b1) ? i_input_data[920 % IN_WIDTH] : ping_storage_data_369 ^ i_input_data[920 % IN_WIDTH];
                default: ping_storage_data_369 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_369;
                endcase
            end else begin
                case (input_count)
                20 / IN_WIDTH: pong_storage_data_369 <= (fillup_transition == 1'b1) ? i_input_data[20 % IN_WIDTH] : pong_storage_data_369 ^ i_input_data[20 % IN_WIDTH];
                226 / IN_WIDTH: pong_storage_data_369 <= (fillup_transition == 1'b1) ? i_input_data[226 % IN_WIDTH] : pong_storage_data_369 ^ i_input_data[226 % IN_WIDTH];
                784 / IN_WIDTH: pong_storage_data_369 <= (fillup_transition == 1'b1) ? i_input_data[784 % IN_WIDTH] : pong_storage_data_369 ^ i_input_data[784 % IN_WIDTH];
                920 / IN_WIDTH: pong_storage_data_369 <= (fillup_transition == 1'b1) ? i_input_data[920 % IN_WIDTH] : pong_storage_data_369 ^ i_input_data[920 % IN_WIDTH];
                default: pong_storage_data_369 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_369;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_369 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_369;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_369 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_369;
            end
        end
    end
end

logic ping_storage_data_370;
logic pong_storage_data_370;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_370 <= 1'b0;
        pong_storage_data_370 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                21 / IN_WIDTH: ping_storage_data_370 <= (fillup_transition == 1'b1) ? i_input_data[21 % IN_WIDTH] : ping_storage_data_370 ^ i_input_data[21 % IN_WIDTH];
                227 / IN_WIDTH: ping_storage_data_370 <= (fillup_transition == 1'b1) ? i_input_data[227 % IN_WIDTH] : ping_storage_data_370 ^ i_input_data[227 % IN_WIDTH];
                785 / IN_WIDTH: ping_storage_data_370 <= (fillup_transition == 1'b1) ? i_input_data[785 % IN_WIDTH] : ping_storage_data_370 ^ i_input_data[785 % IN_WIDTH];
                921 / IN_WIDTH: ping_storage_data_370 <= (fillup_transition == 1'b1) ? i_input_data[921 % IN_WIDTH] : ping_storage_data_370 ^ i_input_data[921 % IN_WIDTH];
                default: ping_storage_data_370 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_370;
                endcase
            end else begin
                case (input_count)
                21 / IN_WIDTH: pong_storage_data_370 <= (fillup_transition == 1'b1) ? i_input_data[21 % IN_WIDTH] : pong_storage_data_370 ^ i_input_data[21 % IN_WIDTH];
                227 / IN_WIDTH: pong_storage_data_370 <= (fillup_transition == 1'b1) ? i_input_data[227 % IN_WIDTH] : pong_storage_data_370 ^ i_input_data[227 % IN_WIDTH];
                785 / IN_WIDTH: pong_storage_data_370 <= (fillup_transition == 1'b1) ? i_input_data[785 % IN_WIDTH] : pong_storage_data_370 ^ i_input_data[785 % IN_WIDTH];
                921 / IN_WIDTH: pong_storage_data_370 <= (fillup_transition == 1'b1) ? i_input_data[921 % IN_WIDTH] : pong_storage_data_370 ^ i_input_data[921 % IN_WIDTH];
                default: pong_storage_data_370 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_370;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_370 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_370;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_370 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_370;
            end
        end
    end
end

logic ping_storage_data_371;
logic pong_storage_data_371;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_371 <= 1'b0;
        pong_storage_data_371 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                22 / IN_WIDTH: ping_storage_data_371 <= (fillup_transition == 1'b1) ? i_input_data[22 % IN_WIDTH] : ping_storage_data_371 ^ i_input_data[22 % IN_WIDTH];
                228 / IN_WIDTH: ping_storage_data_371 <= (fillup_transition == 1'b1) ? i_input_data[228 % IN_WIDTH] : ping_storage_data_371 ^ i_input_data[228 % IN_WIDTH];
                786 / IN_WIDTH: ping_storage_data_371 <= (fillup_transition == 1'b1) ? i_input_data[786 % IN_WIDTH] : ping_storage_data_371 ^ i_input_data[786 % IN_WIDTH];
                922 / IN_WIDTH: ping_storage_data_371 <= (fillup_transition == 1'b1) ? i_input_data[922 % IN_WIDTH] : ping_storage_data_371 ^ i_input_data[922 % IN_WIDTH];
                default: ping_storage_data_371 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_371;
                endcase
            end else begin
                case (input_count)
                22 / IN_WIDTH: pong_storage_data_371 <= (fillup_transition == 1'b1) ? i_input_data[22 % IN_WIDTH] : pong_storage_data_371 ^ i_input_data[22 % IN_WIDTH];
                228 / IN_WIDTH: pong_storage_data_371 <= (fillup_transition == 1'b1) ? i_input_data[228 % IN_WIDTH] : pong_storage_data_371 ^ i_input_data[228 % IN_WIDTH];
                786 / IN_WIDTH: pong_storage_data_371 <= (fillup_transition == 1'b1) ? i_input_data[786 % IN_WIDTH] : pong_storage_data_371 ^ i_input_data[786 % IN_WIDTH];
                922 / IN_WIDTH: pong_storage_data_371 <= (fillup_transition == 1'b1) ? i_input_data[922 % IN_WIDTH] : pong_storage_data_371 ^ i_input_data[922 % IN_WIDTH];
                default: pong_storage_data_371 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_371;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_371 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_371;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_371 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_371;
            end
        end
    end
end

logic ping_storage_data_372;
logic pong_storage_data_372;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_372 <= 1'b0;
        pong_storage_data_372 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                23 / IN_WIDTH: ping_storage_data_372 <= (fillup_transition == 1'b1) ? i_input_data[23 % IN_WIDTH] : ping_storage_data_372 ^ i_input_data[23 % IN_WIDTH];
                229 / IN_WIDTH: ping_storage_data_372 <= (fillup_transition == 1'b1) ? i_input_data[229 % IN_WIDTH] : ping_storage_data_372 ^ i_input_data[229 % IN_WIDTH];
                787 / IN_WIDTH: ping_storage_data_372 <= (fillup_transition == 1'b1) ? i_input_data[787 % IN_WIDTH] : ping_storage_data_372 ^ i_input_data[787 % IN_WIDTH];
                923 / IN_WIDTH: ping_storage_data_372 <= (fillup_transition == 1'b1) ? i_input_data[923 % IN_WIDTH] : ping_storage_data_372 ^ i_input_data[923 % IN_WIDTH];
                default: ping_storage_data_372 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_372;
                endcase
            end else begin
                case (input_count)
                23 / IN_WIDTH: pong_storage_data_372 <= (fillup_transition == 1'b1) ? i_input_data[23 % IN_WIDTH] : pong_storage_data_372 ^ i_input_data[23 % IN_WIDTH];
                229 / IN_WIDTH: pong_storage_data_372 <= (fillup_transition == 1'b1) ? i_input_data[229 % IN_WIDTH] : pong_storage_data_372 ^ i_input_data[229 % IN_WIDTH];
                787 / IN_WIDTH: pong_storage_data_372 <= (fillup_transition == 1'b1) ? i_input_data[787 % IN_WIDTH] : pong_storage_data_372 ^ i_input_data[787 % IN_WIDTH];
                923 / IN_WIDTH: pong_storage_data_372 <= (fillup_transition == 1'b1) ? i_input_data[923 % IN_WIDTH] : pong_storage_data_372 ^ i_input_data[923 % IN_WIDTH];
                default: pong_storage_data_372 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_372;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_372 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_372;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_372 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_372;
            end
        end
    end
end

logic ping_storage_data_373;
logic pong_storage_data_373;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_373 <= 1'b0;
        pong_storage_data_373 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                24 / IN_WIDTH: ping_storage_data_373 <= (fillup_transition == 1'b1) ? i_input_data[24 % IN_WIDTH] : ping_storage_data_373 ^ i_input_data[24 % IN_WIDTH];
                230 / IN_WIDTH: ping_storage_data_373 <= (fillup_transition == 1'b1) ? i_input_data[230 % IN_WIDTH] : ping_storage_data_373 ^ i_input_data[230 % IN_WIDTH];
                788 / IN_WIDTH: ping_storage_data_373 <= (fillup_transition == 1'b1) ? i_input_data[788 % IN_WIDTH] : ping_storage_data_373 ^ i_input_data[788 % IN_WIDTH];
                924 / IN_WIDTH: ping_storage_data_373 <= (fillup_transition == 1'b1) ? i_input_data[924 % IN_WIDTH] : ping_storage_data_373 ^ i_input_data[924 % IN_WIDTH];
                default: ping_storage_data_373 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_373;
                endcase
            end else begin
                case (input_count)
                24 / IN_WIDTH: pong_storage_data_373 <= (fillup_transition == 1'b1) ? i_input_data[24 % IN_WIDTH] : pong_storage_data_373 ^ i_input_data[24 % IN_WIDTH];
                230 / IN_WIDTH: pong_storage_data_373 <= (fillup_transition == 1'b1) ? i_input_data[230 % IN_WIDTH] : pong_storage_data_373 ^ i_input_data[230 % IN_WIDTH];
                788 / IN_WIDTH: pong_storage_data_373 <= (fillup_transition == 1'b1) ? i_input_data[788 % IN_WIDTH] : pong_storage_data_373 ^ i_input_data[788 % IN_WIDTH];
                924 / IN_WIDTH: pong_storage_data_373 <= (fillup_transition == 1'b1) ? i_input_data[924 % IN_WIDTH] : pong_storage_data_373 ^ i_input_data[924 % IN_WIDTH];
                default: pong_storage_data_373 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_373;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_373 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_373;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_373 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_373;
            end
        end
    end
end

logic ping_storage_data_374;
logic pong_storage_data_374;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_374 <= 1'b0;
        pong_storage_data_374 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                25 / IN_WIDTH: ping_storage_data_374 <= (fillup_transition == 1'b1) ? i_input_data[25 % IN_WIDTH] : ping_storage_data_374 ^ i_input_data[25 % IN_WIDTH];
                231 / IN_WIDTH: ping_storage_data_374 <= (fillup_transition == 1'b1) ? i_input_data[231 % IN_WIDTH] : ping_storage_data_374 ^ i_input_data[231 % IN_WIDTH];
                789 / IN_WIDTH: ping_storage_data_374 <= (fillup_transition == 1'b1) ? i_input_data[789 % IN_WIDTH] : ping_storage_data_374 ^ i_input_data[789 % IN_WIDTH];
                925 / IN_WIDTH: ping_storage_data_374 <= (fillup_transition == 1'b1) ? i_input_data[925 % IN_WIDTH] : ping_storage_data_374 ^ i_input_data[925 % IN_WIDTH];
                default: ping_storage_data_374 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_374;
                endcase
            end else begin
                case (input_count)
                25 / IN_WIDTH: pong_storage_data_374 <= (fillup_transition == 1'b1) ? i_input_data[25 % IN_WIDTH] : pong_storage_data_374 ^ i_input_data[25 % IN_WIDTH];
                231 / IN_WIDTH: pong_storage_data_374 <= (fillup_transition == 1'b1) ? i_input_data[231 % IN_WIDTH] : pong_storage_data_374 ^ i_input_data[231 % IN_WIDTH];
                789 / IN_WIDTH: pong_storage_data_374 <= (fillup_transition == 1'b1) ? i_input_data[789 % IN_WIDTH] : pong_storage_data_374 ^ i_input_data[789 % IN_WIDTH];
                925 / IN_WIDTH: pong_storage_data_374 <= (fillup_transition == 1'b1) ? i_input_data[925 % IN_WIDTH] : pong_storage_data_374 ^ i_input_data[925 % IN_WIDTH];
                default: pong_storage_data_374 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_374;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_374 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_374;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_374 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_374;
            end
        end
    end
end

logic ping_storage_data_375;
logic pong_storage_data_375;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_375 <= 1'b0;
        pong_storage_data_375 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                26 / IN_WIDTH: ping_storage_data_375 <= (fillup_transition == 1'b1) ? i_input_data[26 % IN_WIDTH] : ping_storage_data_375 ^ i_input_data[26 % IN_WIDTH];
                232 / IN_WIDTH: ping_storage_data_375 <= (fillup_transition == 1'b1) ? i_input_data[232 % IN_WIDTH] : ping_storage_data_375 ^ i_input_data[232 % IN_WIDTH];
                790 / IN_WIDTH: ping_storage_data_375 <= (fillup_transition == 1'b1) ? i_input_data[790 % IN_WIDTH] : ping_storage_data_375 ^ i_input_data[790 % IN_WIDTH];
                926 / IN_WIDTH: ping_storage_data_375 <= (fillup_transition == 1'b1) ? i_input_data[926 % IN_WIDTH] : ping_storage_data_375 ^ i_input_data[926 % IN_WIDTH];
                default: ping_storage_data_375 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_375;
                endcase
            end else begin
                case (input_count)
                26 / IN_WIDTH: pong_storage_data_375 <= (fillup_transition == 1'b1) ? i_input_data[26 % IN_WIDTH] : pong_storage_data_375 ^ i_input_data[26 % IN_WIDTH];
                232 / IN_WIDTH: pong_storage_data_375 <= (fillup_transition == 1'b1) ? i_input_data[232 % IN_WIDTH] : pong_storage_data_375 ^ i_input_data[232 % IN_WIDTH];
                790 / IN_WIDTH: pong_storage_data_375 <= (fillup_transition == 1'b1) ? i_input_data[790 % IN_WIDTH] : pong_storage_data_375 ^ i_input_data[790 % IN_WIDTH];
                926 / IN_WIDTH: pong_storage_data_375 <= (fillup_transition == 1'b1) ? i_input_data[926 % IN_WIDTH] : pong_storage_data_375 ^ i_input_data[926 % IN_WIDTH];
                default: pong_storage_data_375 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_375;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_375 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_375;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_375 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_375;
            end
        end
    end
end

logic ping_storage_data_376;
logic pong_storage_data_376;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_376 <= 1'b0;
        pong_storage_data_376 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                27 / IN_WIDTH: ping_storage_data_376 <= (fillup_transition == 1'b1) ? i_input_data[27 % IN_WIDTH] : ping_storage_data_376 ^ i_input_data[27 % IN_WIDTH];
                233 / IN_WIDTH: ping_storage_data_376 <= (fillup_transition == 1'b1) ? i_input_data[233 % IN_WIDTH] : ping_storage_data_376 ^ i_input_data[233 % IN_WIDTH];
                791 / IN_WIDTH: ping_storage_data_376 <= (fillup_transition == 1'b1) ? i_input_data[791 % IN_WIDTH] : ping_storage_data_376 ^ i_input_data[791 % IN_WIDTH];
                927 / IN_WIDTH: ping_storage_data_376 <= (fillup_transition == 1'b1) ? i_input_data[927 % IN_WIDTH] : ping_storage_data_376 ^ i_input_data[927 % IN_WIDTH];
                default: ping_storage_data_376 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_376;
                endcase
            end else begin
                case (input_count)
                27 / IN_WIDTH: pong_storage_data_376 <= (fillup_transition == 1'b1) ? i_input_data[27 % IN_WIDTH] : pong_storage_data_376 ^ i_input_data[27 % IN_WIDTH];
                233 / IN_WIDTH: pong_storage_data_376 <= (fillup_transition == 1'b1) ? i_input_data[233 % IN_WIDTH] : pong_storage_data_376 ^ i_input_data[233 % IN_WIDTH];
                791 / IN_WIDTH: pong_storage_data_376 <= (fillup_transition == 1'b1) ? i_input_data[791 % IN_WIDTH] : pong_storage_data_376 ^ i_input_data[791 % IN_WIDTH];
                927 / IN_WIDTH: pong_storage_data_376 <= (fillup_transition == 1'b1) ? i_input_data[927 % IN_WIDTH] : pong_storage_data_376 ^ i_input_data[927 % IN_WIDTH];
                default: pong_storage_data_376 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_376;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_376 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_376;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_376 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_376;
            end
        end
    end
end

logic ping_storage_data_377;
logic pong_storage_data_377;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_377 <= 1'b0;
        pong_storage_data_377 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                28 / IN_WIDTH: ping_storage_data_377 <= (fillup_transition == 1'b1) ? i_input_data[28 % IN_WIDTH] : ping_storage_data_377 ^ i_input_data[28 % IN_WIDTH];
                234 / IN_WIDTH: ping_storage_data_377 <= (fillup_transition == 1'b1) ? i_input_data[234 % IN_WIDTH] : ping_storage_data_377 ^ i_input_data[234 % IN_WIDTH];
                792 / IN_WIDTH: ping_storage_data_377 <= (fillup_transition == 1'b1) ? i_input_data[792 % IN_WIDTH] : ping_storage_data_377 ^ i_input_data[792 % IN_WIDTH];
                928 / IN_WIDTH: ping_storage_data_377 <= (fillup_transition == 1'b1) ? i_input_data[928 % IN_WIDTH] : ping_storage_data_377 ^ i_input_data[928 % IN_WIDTH];
                default: ping_storage_data_377 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_377;
                endcase
            end else begin
                case (input_count)
                28 / IN_WIDTH: pong_storage_data_377 <= (fillup_transition == 1'b1) ? i_input_data[28 % IN_WIDTH] : pong_storage_data_377 ^ i_input_data[28 % IN_WIDTH];
                234 / IN_WIDTH: pong_storage_data_377 <= (fillup_transition == 1'b1) ? i_input_data[234 % IN_WIDTH] : pong_storage_data_377 ^ i_input_data[234 % IN_WIDTH];
                792 / IN_WIDTH: pong_storage_data_377 <= (fillup_transition == 1'b1) ? i_input_data[792 % IN_WIDTH] : pong_storage_data_377 ^ i_input_data[792 % IN_WIDTH];
                928 / IN_WIDTH: pong_storage_data_377 <= (fillup_transition == 1'b1) ? i_input_data[928 % IN_WIDTH] : pong_storage_data_377 ^ i_input_data[928 % IN_WIDTH];
                default: pong_storage_data_377 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_377;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_377 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_377;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_377 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_377;
            end
        end
    end
end

logic ping_storage_data_378;
logic pong_storage_data_378;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_378 <= 1'b0;
        pong_storage_data_378 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                29 / IN_WIDTH: ping_storage_data_378 <= (fillup_transition == 1'b1) ? i_input_data[29 % IN_WIDTH] : ping_storage_data_378 ^ i_input_data[29 % IN_WIDTH];
                235 / IN_WIDTH: ping_storage_data_378 <= (fillup_transition == 1'b1) ? i_input_data[235 % IN_WIDTH] : ping_storage_data_378 ^ i_input_data[235 % IN_WIDTH];
                793 / IN_WIDTH: ping_storage_data_378 <= (fillup_transition == 1'b1) ? i_input_data[793 % IN_WIDTH] : ping_storage_data_378 ^ i_input_data[793 % IN_WIDTH];
                929 / IN_WIDTH: ping_storage_data_378 <= (fillup_transition == 1'b1) ? i_input_data[929 % IN_WIDTH] : ping_storage_data_378 ^ i_input_data[929 % IN_WIDTH];
                default: ping_storage_data_378 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_378;
                endcase
            end else begin
                case (input_count)
                29 / IN_WIDTH: pong_storage_data_378 <= (fillup_transition == 1'b1) ? i_input_data[29 % IN_WIDTH] : pong_storage_data_378 ^ i_input_data[29 % IN_WIDTH];
                235 / IN_WIDTH: pong_storage_data_378 <= (fillup_transition == 1'b1) ? i_input_data[235 % IN_WIDTH] : pong_storage_data_378 ^ i_input_data[235 % IN_WIDTH];
                793 / IN_WIDTH: pong_storage_data_378 <= (fillup_transition == 1'b1) ? i_input_data[793 % IN_WIDTH] : pong_storage_data_378 ^ i_input_data[793 % IN_WIDTH];
                929 / IN_WIDTH: pong_storage_data_378 <= (fillup_transition == 1'b1) ? i_input_data[929 % IN_WIDTH] : pong_storage_data_378 ^ i_input_data[929 % IN_WIDTH];
                default: pong_storage_data_378 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_378;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_378 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_378;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_378 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_378;
            end
        end
    end
end

logic ping_storage_data_379;
logic pong_storage_data_379;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_379 <= 1'b0;
        pong_storage_data_379 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                30 / IN_WIDTH: ping_storage_data_379 <= (fillup_transition == 1'b1) ? i_input_data[30 % IN_WIDTH] : ping_storage_data_379 ^ i_input_data[30 % IN_WIDTH];
                236 / IN_WIDTH: ping_storage_data_379 <= (fillup_transition == 1'b1) ? i_input_data[236 % IN_WIDTH] : ping_storage_data_379 ^ i_input_data[236 % IN_WIDTH];
                794 / IN_WIDTH: ping_storage_data_379 <= (fillup_transition == 1'b1) ? i_input_data[794 % IN_WIDTH] : ping_storage_data_379 ^ i_input_data[794 % IN_WIDTH];
                930 / IN_WIDTH: ping_storage_data_379 <= (fillup_transition == 1'b1) ? i_input_data[930 % IN_WIDTH] : ping_storage_data_379 ^ i_input_data[930 % IN_WIDTH];
                default: ping_storage_data_379 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_379;
                endcase
            end else begin
                case (input_count)
                30 / IN_WIDTH: pong_storage_data_379 <= (fillup_transition == 1'b1) ? i_input_data[30 % IN_WIDTH] : pong_storage_data_379 ^ i_input_data[30 % IN_WIDTH];
                236 / IN_WIDTH: pong_storage_data_379 <= (fillup_transition == 1'b1) ? i_input_data[236 % IN_WIDTH] : pong_storage_data_379 ^ i_input_data[236 % IN_WIDTH];
                794 / IN_WIDTH: pong_storage_data_379 <= (fillup_transition == 1'b1) ? i_input_data[794 % IN_WIDTH] : pong_storage_data_379 ^ i_input_data[794 % IN_WIDTH];
                930 / IN_WIDTH: pong_storage_data_379 <= (fillup_transition == 1'b1) ? i_input_data[930 % IN_WIDTH] : pong_storage_data_379 ^ i_input_data[930 % IN_WIDTH];
                default: pong_storage_data_379 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_379;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_379 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_379;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_379 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_379;
            end
        end
    end
end

logic ping_storage_data_380;
logic pong_storage_data_380;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_380 <= 1'b0;
        pong_storage_data_380 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                31 / IN_WIDTH: ping_storage_data_380 <= (fillup_transition == 1'b1) ? i_input_data[31 % IN_WIDTH] : ping_storage_data_380 ^ i_input_data[31 % IN_WIDTH];
                237 / IN_WIDTH: ping_storage_data_380 <= (fillup_transition == 1'b1) ? i_input_data[237 % IN_WIDTH] : ping_storage_data_380 ^ i_input_data[237 % IN_WIDTH];
                795 / IN_WIDTH: ping_storage_data_380 <= (fillup_transition == 1'b1) ? i_input_data[795 % IN_WIDTH] : ping_storage_data_380 ^ i_input_data[795 % IN_WIDTH];
                931 / IN_WIDTH: ping_storage_data_380 <= (fillup_transition == 1'b1) ? i_input_data[931 % IN_WIDTH] : ping_storage_data_380 ^ i_input_data[931 % IN_WIDTH];
                default: ping_storage_data_380 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_380;
                endcase
            end else begin
                case (input_count)
                31 / IN_WIDTH: pong_storage_data_380 <= (fillup_transition == 1'b1) ? i_input_data[31 % IN_WIDTH] : pong_storage_data_380 ^ i_input_data[31 % IN_WIDTH];
                237 / IN_WIDTH: pong_storage_data_380 <= (fillup_transition == 1'b1) ? i_input_data[237 % IN_WIDTH] : pong_storage_data_380 ^ i_input_data[237 % IN_WIDTH];
                795 / IN_WIDTH: pong_storage_data_380 <= (fillup_transition == 1'b1) ? i_input_data[795 % IN_WIDTH] : pong_storage_data_380 ^ i_input_data[795 % IN_WIDTH];
                931 / IN_WIDTH: pong_storage_data_380 <= (fillup_transition == 1'b1) ? i_input_data[931 % IN_WIDTH] : pong_storage_data_380 ^ i_input_data[931 % IN_WIDTH];
                default: pong_storage_data_380 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_380;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_380 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_380;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_380 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_380;
            end
        end
    end
end

logic ping_storage_data_381;
logic pong_storage_data_381;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_381 <= 1'b0;
        pong_storage_data_381 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                32 / IN_WIDTH: ping_storage_data_381 <= (fillup_transition == 1'b1) ? i_input_data[32 % IN_WIDTH] : ping_storage_data_381 ^ i_input_data[32 % IN_WIDTH];
                238 / IN_WIDTH: ping_storage_data_381 <= (fillup_transition == 1'b1) ? i_input_data[238 % IN_WIDTH] : ping_storage_data_381 ^ i_input_data[238 % IN_WIDTH];
                796 / IN_WIDTH: ping_storage_data_381 <= (fillup_transition == 1'b1) ? i_input_data[796 % IN_WIDTH] : ping_storage_data_381 ^ i_input_data[796 % IN_WIDTH];
                932 / IN_WIDTH: ping_storage_data_381 <= (fillup_transition == 1'b1) ? i_input_data[932 % IN_WIDTH] : ping_storage_data_381 ^ i_input_data[932 % IN_WIDTH];
                default: ping_storage_data_381 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_381;
                endcase
            end else begin
                case (input_count)
                32 / IN_WIDTH: pong_storage_data_381 <= (fillup_transition == 1'b1) ? i_input_data[32 % IN_WIDTH] : pong_storage_data_381 ^ i_input_data[32 % IN_WIDTH];
                238 / IN_WIDTH: pong_storage_data_381 <= (fillup_transition == 1'b1) ? i_input_data[238 % IN_WIDTH] : pong_storage_data_381 ^ i_input_data[238 % IN_WIDTH];
                796 / IN_WIDTH: pong_storage_data_381 <= (fillup_transition == 1'b1) ? i_input_data[796 % IN_WIDTH] : pong_storage_data_381 ^ i_input_data[796 % IN_WIDTH];
                932 / IN_WIDTH: pong_storage_data_381 <= (fillup_transition == 1'b1) ? i_input_data[932 % IN_WIDTH] : pong_storage_data_381 ^ i_input_data[932 % IN_WIDTH];
                default: pong_storage_data_381 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_381;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_381 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_381;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_381 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_381;
            end
        end
    end
end

logic ping_storage_data_382;
logic pong_storage_data_382;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_382 <= 1'b0;
        pong_storage_data_382 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                33 / IN_WIDTH: ping_storage_data_382 <= (fillup_transition == 1'b1) ? i_input_data[33 % IN_WIDTH] : ping_storage_data_382 ^ i_input_data[33 % IN_WIDTH];
                239 / IN_WIDTH: ping_storage_data_382 <= (fillup_transition == 1'b1) ? i_input_data[239 % IN_WIDTH] : ping_storage_data_382 ^ i_input_data[239 % IN_WIDTH];
                797 / IN_WIDTH: ping_storage_data_382 <= (fillup_transition == 1'b1) ? i_input_data[797 % IN_WIDTH] : ping_storage_data_382 ^ i_input_data[797 % IN_WIDTH];
                933 / IN_WIDTH: ping_storage_data_382 <= (fillup_transition == 1'b1) ? i_input_data[933 % IN_WIDTH] : ping_storage_data_382 ^ i_input_data[933 % IN_WIDTH];
                default: ping_storage_data_382 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_382;
                endcase
            end else begin
                case (input_count)
                33 / IN_WIDTH: pong_storage_data_382 <= (fillup_transition == 1'b1) ? i_input_data[33 % IN_WIDTH] : pong_storage_data_382 ^ i_input_data[33 % IN_WIDTH];
                239 / IN_WIDTH: pong_storage_data_382 <= (fillup_transition == 1'b1) ? i_input_data[239 % IN_WIDTH] : pong_storage_data_382 ^ i_input_data[239 % IN_WIDTH];
                797 / IN_WIDTH: pong_storage_data_382 <= (fillup_transition == 1'b1) ? i_input_data[797 % IN_WIDTH] : pong_storage_data_382 ^ i_input_data[797 % IN_WIDTH];
                933 / IN_WIDTH: pong_storage_data_382 <= (fillup_transition == 1'b1) ? i_input_data[933 % IN_WIDTH] : pong_storage_data_382 ^ i_input_data[933 % IN_WIDTH];
                default: pong_storage_data_382 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_382;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_382 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_382;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_382 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_382;
            end
        end
    end
end

logic ping_storage_data_383;
logic pong_storage_data_383;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_383 <= 1'b0;
        pong_storage_data_383 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                34 / IN_WIDTH: ping_storage_data_383 <= (fillup_transition == 1'b1) ? i_input_data[34 % IN_WIDTH] : ping_storage_data_383 ^ i_input_data[34 % IN_WIDTH];
                240 / IN_WIDTH: ping_storage_data_383 <= (fillup_transition == 1'b1) ? i_input_data[240 % IN_WIDTH] : ping_storage_data_383 ^ i_input_data[240 % IN_WIDTH];
                798 / IN_WIDTH: ping_storage_data_383 <= (fillup_transition == 1'b1) ? i_input_data[798 % IN_WIDTH] : ping_storage_data_383 ^ i_input_data[798 % IN_WIDTH];
                934 / IN_WIDTH: ping_storage_data_383 <= (fillup_transition == 1'b1) ? i_input_data[934 % IN_WIDTH] : ping_storage_data_383 ^ i_input_data[934 % IN_WIDTH];
                default: ping_storage_data_383 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_383;
                endcase
            end else begin
                case (input_count)
                34 / IN_WIDTH: pong_storage_data_383 <= (fillup_transition == 1'b1) ? i_input_data[34 % IN_WIDTH] : pong_storage_data_383 ^ i_input_data[34 % IN_WIDTH];
                240 / IN_WIDTH: pong_storage_data_383 <= (fillup_transition == 1'b1) ? i_input_data[240 % IN_WIDTH] : pong_storage_data_383 ^ i_input_data[240 % IN_WIDTH];
                798 / IN_WIDTH: pong_storage_data_383 <= (fillup_transition == 1'b1) ? i_input_data[798 % IN_WIDTH] : pong_storage_data_383 ^ i_input_data[798 % IN_WIDTH];
                934 / IN_WIDTH: pong_storage_data_383 <= (fillup_transition == 1'b1) ? i_input_data[934 % IN_WIDTH] : pong_storage_data_383 ^ i_input_data[934 % IN_WIDTH];
                default: pong_storage_data_383 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_383;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_383 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_383;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_383 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_383;
            end
        end
    end
end

logic ping_storage_data_384;
logic pong_storage_data_384;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_384 <= 1'b0;
        pong_storage_data_384 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                249 / IN_WIDTH: ping_storage_data_384 <= (fillup_transition == 1'b1) ? i_input_data[249 % IN_WIDTH] : ping_storage_data_384 ^ i_input_data[249 % IN_WIDTH];
                588 / IN_WIDTH: ping_storage_data_384 <= (fillup_transition == 1'b1) ? i_input_data[588 % IN_WIDTH] : ping_storage_data_384 ^ i_input_data[588 % IN_WIDTH];
                919 / IN_WIDTH: ping_storage_data_384 <= (fillup_transition == 1'b1) ? i_input_data[919 % IN_WIDTH] : ping_storage_data_384 ^ i_input_data[919 % IN_WIDTH];
                984 / IN_WIDTH: ping_storage_data_384 <= (fillup_transition == 1'b1) ? i_input_data[984 % IN_WIDTH] : ping_storage_data_384 ^ i_input_data[984 % IN_WIDTH];
                default: ping_storage_data_384 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_384;
                endcase
            end else begin
                case (input_count)
                249 / IN_WIDTH: pong_storage_data_384 <= (fillup_transition == 1'b1) ? i_input_data[249 % IN_WIDTH] : pong_storage_data_384 ^ i_input_data[249 % IN_WIDTH];
                588 / IN_WIDTH: pong_storage_data_384 <= (fillup_transition == 1'b1) ? i_input_data[588 % IN_WIDTH] : pong_storage_data_384 ^ i_input_data[588 % IN_WIDTH];
                919 / IN_WIDTH: pong_storage_data_384 <= (fillup_transition == 1'b1) ? i_input_data[919 % IN_WIDTH] : pong_storage_data_384 ^ i_input_data[919 % IN_WIDTH];
                984 / IN_WIDTH: pong_storage_data_384 <= (fillup_transition == 1'b1) ? i_input_data[984 % IN_WIDTH] : pong_storage_data_384 ^ i_input_data[984 % IN_WIDTH];
                default: pong_storage_data_384 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_384;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_384 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_384;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_384 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_384;
            end
        end
    end
end

logic ping_storage_data_385;
logic pong_storage_data_385;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_385 <= 1'b0;
        pong_storage_data_385 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                250 / IN_WIDTH: ping_storage_data_385 <= (fillup_transition == 1'b1) ? i_input_data[250 % IN_WIDTH] : ping_storage_data_385 ^ i_input_data[250 % IN_WIDTH];
                589 / IN_WIDTH: ping_storage_data_385 <= (fillup_transition == 1'b1) ? i_input_data[589 % IN_WIDTH] : ping_storage_data_385 ^ i_input_data[589 % IN_WIDTH];
                920 / IN_WIDTH: ping_storage_data_385 <= (fillup_transition == 1'b1) ? i_input_data[920 % IN_WIDTH] : ping_storage_data_385 ^ i_input_data[920 % IN_WIDTH];
                985 / IN_WIDTH: ping_storage_data_385 <= (fillup_transition == 1'b1) ? i_input_data[985 % IN_WIDTH] : ping_storage_data_385 ^ i_input_data[985 % IN_WIDTH];
                default: ping_storage_data_385 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_385;
                endcase
            end else begin
                case (input_count)
                250 / IN_WIDTH: pong_storage_data_385 <= (fillup_transition == 1'b1) ? i_input_data[250 % IN_WIDTH] : pong_storage_data_385 ^ i_input_data[250 % IN_WIDTH];
                589 / IN_WIDTH: pong_storage_data_385 <= (fillup_transition == 1'b1) ? i_input_data[589 % IN_WIDTH] : pong_storage_data_385 ^ i_input_data[589 % IN_WIDTH];
                920 / IN_WIDTH: pong_storage_data_385 <= (fillup_transition == 1'b1) ? i_input_data[920 % IN_WIDTH] : pong_storage_data_385 ^ i_input_data[920 % IN_WIDTH];
                985 / IN_WIDTH: pong_storage_data_385 <= (fillup_transition == 1'b1) ? i_input_data[985 % IN_WIDTH] : pong_storage_data_385 ^ i_input_data[985 % IN_WIDTH];
                default: pong_storage_data_385 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_385;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_385 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_385;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_385 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_385;
            end
        end
    end
end

logic ping_storage_data_386;
logic pong_storage_data_386;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_386 <= 1'b0;
        pong_storage_data_386 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                251 / IN_WIDTH: ping_storage_data_386 <= (fillup_transition == 1'b1) ? i_input_data[251 % IN_WIDTH] : ping_storage_data_386 ^ i_input_data[251 % IN_WIDTH];
                590 / IN_WIDTH: ping_storage_data_386 <= (fillup_transition == 1'b1) ? i_input_data[590 % IN_WIDTH] : ping_storage_data_386 ^ i_input_data[590 % IN_WIDTH];
                921 / IN_WIDTH: ping_storage_data_386 <= (fillup_transition == 1'b1) ? i_input_data[921 % IN_WIDTH] : ping_storage_data_386 ^ i_input_data[921 % IN_WIDTH];
                986 / IN_WIDTH: ping_storage_data_386 <= (fillup_transition == 1'b1) ? i_input_data[986 % IN_WIDTH] : ping_storage_data_386 ^ i_input_data[986 % IN_WIDTH];
                default: ping_storage_data_386 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_386;
                endcase
            end else begin
                case (input_count)
                251 / IN_WIDTH: pong_storage_data_386 <= (fillup_transition == 1'b1) ? i_input_data[251 % IN_WIDTH] : pong_storage_data_386 ^ i_input_data[251 % IN_WIDTH];
                590 / IN_WIDTH: pong_storage_data_386 <= (fillup_transition == 1'b1) ? i_input_data[590 % IN_WIDTH] : pong_storage_data_386 ^ i_input_data[590 % IN_WIDTH];
                921 / IN_WIDTH: pong_storage_data_386 <= (fillup_transition == 1'b1) ? i_input_data[921 % IN_WIDTH] : pong_storage_data_386 ^ i_input_data[921 % IN_WIDTH];
                986 / IN_WIDTH: pong_storage_data_386 <= (fillup_transition == 1'b1) ? i_input_data[986 % IN_WIDTH] : pong_storage_data_386 ^ i_input_data[986 % IN_WIDTH];
                default: pong_storage_data_386 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_386;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_386 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_386;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_386 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_386;
            end
        end
    end
end

logic ping_storage_data_387;
logic pong_storage_data_387;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_387 <= 1'b0;
        pong_storage_data_387 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                252 / IN_WIDTH: ping_storage_data_387 <= (fillup_transition == 1'b1) ? i_input_data[252 % IN_WIDTH] : ping_storage_data_387 ^ i_input_data[252 % IN_WIDTH];
                591 / IN_WIDTH: ping_storage_data_387 <= (fillup_transition == 1'b1) ? i_input_data[591 % IN_WIDTH] : ping_storage_data_387 ^ i_input_data[591 % IN_WIDTH];
                922 / IN_WIDTH: ping_storage_data_387 <= (fillup_transition == 1'b1) ? i_input_data[922 % IN_WIDTH] : ping_storage_data_387 ^ i_input_data[922 % IN_WIDTH];
                987 / IN_WIDTH: ping_storage_data_387 <= (fillup_transition == 1'b1) ? i_input_data[987 % IN_WIDTH] : ping_storage_data_387 ^ i_input_data[987 % IN_WIDTH];
                default: ping_storage_data_387 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_387;
                endcase
            end else begin
                case (input_count)
                252 / IN_WIDTH: pong_storage_data_387 <= (fillup_transition == 1'b1) ? i_input_data[252 % IN_WIDTH] : pong_storage_data_387 ^ i_input_data[252 % IN_WIDTH];
                591 / IN_WIDTH: pong_storage_data_387 <= (fillup_transition == 1'b1) ? i_input_data[591 % IN_WIDTH] : pong_storage_data_387 ^ i_input_data[591 % IN_WIDTH];
                922 / IN_WIDTH: pong_storage_data_387 <= (fillup_transition == 1'b1) ? i_input_data[922 % IN_WIDTH] : pong_storage_data_387 ^ i_input_data[922 % IN_WIDTH];
                987 / IN_WIDTH: pong_storage_data_387 <= (fillup_transition == 1'b1) ? i_input_data[987 % IN_WIDTH] : pong_storage_data_387 ^ i_input_data[987 % IN_WIDTH];
                default: pong_storage_data_387 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_387;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_387 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_387;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_387 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_387;
            end
        end
    end
end

logic ping_storage_data_388;
logic pong_storage_data_388;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_388 <= 1'b0;
        pong_storage_data_388 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                253 / IN_WIDTH: ping_storage_data_388 <= (fillup_transition == 1'b1) ? i_input_data[253 % IN_WIDTH] : ping_storage_data_388 ^ i_input_data[253 % IN_WIDTH];
                592 / IN_WIDTH: ping_storage_data_388 <= (fillup_transition == 1'b1) ? i_input_data[592 % IN_WIDTH] : ping_storage_data_388 ^ i_input_data[592 % IN_WIDTH];
                923 / IN_WIDTH: ping_storage_data_388 <= (fillup_transition == 1'b1) ? i_input_data[923 % IN_WIDTH] : ping_storage_data_388 ^ i_input_data[923 % IN_WIDTH];
                988 / IN_WIDTH: ping_storage_data_388 <= (fillup_transition == 1'b1) ? i_input_data[988 % IN_WIDTH] : ping_storage_data_388 ^ i_input_data[988 % IN_WIDTH];
                default: ping_storage_data_388 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_388;
                endcase
            end else begin
                case (input_count)
                253 / IN_WIDTH: pong_storage_data_388 <= (fillup_transition == 1'b1) ? i_input_data[253 % IN_WIDTH] : pong_storage_data_388 ^ i_input_data[253 % IN_WIDTH];
                592 / IN_WIDTH: pong_storage_data_388 <= (fillup_transition == 1'b1) ? i_input_data[592 % IN_WIDTH] : pong_storage_data_388 ^ i_input_data[592 % IN_WIDTH];
                923 / IN_WIDTH: pong_storage_data_388 <= (fillup_transition == 1'b1) ? i_input_data[923 % IN_WIDTH] : pong_storage_data_388 ^ i_input_data[923 % IN_WIDTH];
                988 / IN_WIDTH: pong_storage_data_388 <= (fillup_transition == 1'b1) ? i_input_data[988 % IN_WIDTH] : pong_storage_data_388 ^ i_input_data[988 % IN_WIDTH];
                default: pong_storage_data_388 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_388;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_388 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_388;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_388 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_388;
            end
        end
    end
end

logic ping_storage_data_389;
logic pong_storage_data_389;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_389 <= 1'b0;
        pong_storage_data_389 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                254 / IN_WIDTH: ping_storage_data_389 <= (fillup_transition == 1'b1) ? i_input_data[254 % IN_WIDTH] : ping_storage_data_389 ^ i_input_data[254 % IN_WIDTH];
                593 / IN_WIDTH: ping_storage_data_389 <= (fillup_transition == 1'b1) ? i_input_data[593 % IN_WIDTH] : ping_storage_data_389 ^ i_input_data[593 % IN_WIDTH];
                924 / IN_WIDTH: ping_storage_data_389 <= (fillup_transition == 1'b1) ? i_input_data[924 % IN_WIDTH] : ping_storage_data_389 ^ i_input_data[924 % IN_WIDTH];
                989 / IN_WIDTH: ping_storage_data_389 <= (fillup_transition == 1'b1) ? i_input_data[989 % IN_WIDTH] : ping_storage_data_389 ^ i_input_data[989 % IN_WIDTH];
                default: ping_storage_data_389 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_389;
                endcase
            end else begin
                case (input_count)
                254 / IN_WIDTH: pong_storage_data_389 <= (fillup_transition == 1'b1) ? i_input_data[254 % IN_WIDTH] : pong_storage_data_389 ^ i_input_data[254 % IN_WIDTH];
                593 / IN_WIDTH: pong_storage_data_389 <= (fillup_transition == 1'b1) ? i_input_data[593 % IN_WIDTH] : pong_storage_data_389 ^ i_input_data[593 % IN_WIDTH];
                924 / IN_WIDTH: pong_storage_data_389 <= (fillup_transition == 1'b1) ? i_input_data[924 % IN_WIDTH] : pong_storage_data_389 ^ i_input_data[924 % IN_WIDTH];
                989 / IN_WIDTH: pong_storage_data_389 <= (fillup_transition == 1'b1) ? i_input_data[989 % IN_WIDTH] : pong_storage_data_389 ^ i_input_data[989 % IN_WIDTH];
                default: pong_storage_data_389 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_389;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_389 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_389;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_389 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_389;
            end
        end
    end
end

logic ping_storage_data_390;
logic pong_storage_data_390;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_390 <= 1'b0;
        pong_storage_data_390 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                255 / IN_WIDTH: ping_storage_data_390 <= (fillup_transition == 1'b1) ? i_input_data[255 % IN_WIDTH] : ping_storage_data_390 ^ i_input_data[255 % IN_WIDTH];
                594 / IN_WIDTH: ping_storage_data_390 <= (fillup_transition == 1'b1) ? i_input_data[594 % IN_WIDTH] : ping_storage_data_390 ^ i_input_data[594 % IN_WIDTH];
                925 / IN_WIDTH: ping_storage_data_390 <= (fillup_transition == 1'b1) ? i_input_data[925 % IN_WIDTH] : ping_storage_data_390 ^ i_input_data[925 % IN_WIDTH];
                990 / IN_WIDTH: ping_storage_data_390 <= (fillup_transition == 1'b1) ? i_input_data[990 % IN_WIDTH] : ping_storage_data_390 ^ i_input_data[990 % IN_WIDTH];
                default: ping_storage_data_390 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_390;
                endcase
            end else begin
                case (input_count)
                255 / IN_WIDTH: pong_storage_data_390 <= (fillup_transition == 1'b1) ? i_input_data[255 % IN_WIDTH] : pong_storage_data_390 ^ i_input_data[255 % IN_WIDTH];
                594 / IN_WIDTH: pong_storage_data_390 <= (fillup_transition == 1'b1) ? i_input_data[594 % IN_WIDTH] : pong_storage_data_390 ^ i_input_data[594 % IN_WIDTH];
                925 / IN_WIDTH: pong_storage_data_390 <= (fillup_transition == 1'b1) ? i_input_data[925 % IN_WIDTH] : pong_storage_data_390 ^ i_input_data[925 % IN_WIDTH];
                990 / IN_WIDTH: pong_storage_data_390 <= (fillup_transition == 1'b1) ? i_input_data[990 % IN_WIDTH] : pong_storage_data_390 ^ i_input_data[990 % IN_WIDTH];
                default: pong_storage_data_390 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_390;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_390 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_390;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_390 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_390;
            end
        end
    end
end

logic ping_storage_data_391;
logic pong_storage_data_391;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_391 <= 1'b0;
        pong_storage_data_391 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                256 / IN_WIDTH: ping_storage_data_391 <= (fillup_transition == 1'b1) ? i_input_data[256 % IN_WIDTH] : ping_storage_data_391 ^ i_input_data[256 % IN_WIDTH];
                595 / IN_WIDTH: ping_storage_data_391 <= (fillup_transition == 1'b1) ? i_input_data[595 % IN_WIDTH] : ping_storage_data_391 ^ i_input_data[595 % IN_WIDTH];
                926 / IN_WIDTH: ping_storage_data_391 <= (fillup_transition == 1'b1) ? i_input_data[926 % IN_WIDTH] : ping_storage_data_391 ^ i_input_data[926 % IN_WIDTH];
                991 / IN_WIDTH: ping_storage_data_391 <= (fillup_transition == 1'b1) ? i_input_data[991 % IN_WIDTH] : ping_storage_data_391 ^ i_input_data[991 % IN_WIDTH];
                default: ping_storage_data_391 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_391;
                endcase
            end else begin
                case (input_count)
                256 / IN_WIDTH: pong_storage_data_391 <= (fillup_transition == 1'b1) ? i_input_data[256 % IN_WIDTH] : pong_storage_data_391 ^ i_input_data[256 % IN_WIDTH];
                595 / IN_WIDTH: pong_storage_data_391 <= (fillup_transition == 1'b1) ? i_input_data[595 % IN_WIDTH] : pong_storage_data_391 ^ i_input_data[595 % IN_WIDTH];
                926 / IN_WIDTH: pong_storage_data_391 <= (fillup_transition == 1'b1) ? i_input_data[926 % IN_WIDTH] : pong_storage_data_391 ^ i_input_data[926 % IN_WIDTH];
                991 / IN_WIDTH: pong_storage_data_391 <= (fillup_transition == 1'b1) ? i_input_data[991 % IN_WIDTH] : pong_storage_data_391 ^ i_input_data[991 % IN_WIDTH];
                default: pong_storage_data_391 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_391;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_391 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_391;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_391 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_391;
            end
        end
    end
end

logic ping_storage_data_392;
logic pong_storage_data_392;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_392 <= 1'b0;
        pong_storage_data_392 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                257 / IN_WIDTH: ping_storage_data_392 <= (fillup_transition == 1'b1) ? i_input_data[257 % IN_WIDTH] : ping_storage_data_392 ^ i_input_data[257 % IN_WIDTH];
                596 / IN_WIDTH: ping_storage_data_392 <= (fillup_transition == 1'b1) ? i_input_data[596 % IN_WIDTH] : ping_storage_data_392 ^ i_input_data[596 % IN_WIDTH];
                927 / IN_WIDTH: ping_storage_data_392 <= (fillup_transition == 1'b1) ? i_input_data[927 % IN_WIDTH] : ping_storage_data_392 ^ i_input_data[927 % IN_WIDTH];
                992 / IN_WIDTH: ping_storage_data_392 <= (fillup_transition == 1'b1) ? i_input_data[992 % IN_WIDTH] : ping_storage_data_392 ^ i_input_data[992 % IN_WIDTH];
                default: ping_storage_data_392 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_392;
                endcase
            end else begin
                case (input_count)
                257 / IN_WIDTH: pong_storage_data_392 <= (fillup_transition == 1'b1) ? i_input_data[257 % IN_WIDTH] : pong_storage_data_392 ^ i_input_data[257 % IN_WIDTH];
                596 / IN_WIDTH: pong_storage_data_392 <= (fillup_transition == 1'b1) ? i_input_data[596 % IN_WIDTH] : pong_storage_data_392 ^ i_input_data[596 % IN_WIDTH];
                927 / IN_WIDTH: pong_storage_data_392 <= (fillup_transition == 1'b1) ? i_input_data[927 % IN_WIDTH] : pong_storage_data_392 ^ i_input_data[927 % IN_WIDTH];
                992 / IN_WIDTH: pong_storage_data_392 <= (fillup_transition == 1'b1) ? i_input_data[992 % IN_WIDTH] : pong_storage_data_392 ^ i_input_data[992 % IN_WIDTH];
                default: pong_storage_data_392 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_392;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_392 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_392;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_392 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_392;
            end
        end
    end
end

logic ping_storage_data_393;
logic pong_storage_data_393;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_393 <= 1'b0;
        pong_storage_data_393 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                258 / IN_WIDTH: ping_storage_data_393 <= (fillup_transition == 1'b1) ? i_input_data[258 % IN_WIDTH] : ping_storage_data_393 ^ i_input_data[258 % IN_WIDTH];
                597 / IN_WIDTH: ping_storage_data_393 <= (fillup_transition == 1'b1) ? i_input_data[597 % IN_WIDTH] : ping_storage_data_393 ^ i_input_data[597 % IN_WIDTH];
                928 / IN_WIDTH: ping_storage_data_393 <= (fillup_transition == 1'b1) ? i_input_data[928 % IN_WIDTH] : ping_storage_data_393 ^ i_input_data[928 % IN_WIDTH];
                993 / IN_WIDTH: ping_storage_data_393 <= (fillup_transition == 1'b1) ? i_input_data[993 % IN_WIDTH] : ping_storage_data_393 ^ i_input_data[993 % IN_WIDTH];
                default: ping_storage_data_393 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_393;
                endcase
            end else begin
                case (input_count)
                258 / IN_WIDTH: pong_storage_data_393 <= (fillup_transition == 1'b1) ? i_input_data[258 % IN_WIDTH] : pong_storage_data_393 ^ i_input_data[258 % IN_WIDTH];
                597 / IN_WIDTH: pong_storage_data_393 <= (fillup_transition == 1'b1) ? i_input_data[597 % IN_WIDTH] : pong_storage_data_393 ^ i_input_data[597 % IN_WIDTH];
                928 / IN_WIDTH: pong_storage_data_393 <= (fillup_transition == 1'b1) ? i_input_data[928 % IN_WIDTH] : pong_storage_data_393 ^ i_input_data[928 % IN_WIDTH];
                993 / IN_WIDTH: pong_storage_data_393 <= (fillup_transition == 1'b1) ? i_input_data[993 % IN_WIDTH] : pong_storage_data_393 ^ i_input_data[993 % IN_WIDTH];
                default: pong_storage_data_393 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_393;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_393 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_393;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_393 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_393;
            end
        end
    end
end

logic ping_storage_data_394;
logic pong_storage_data_394;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_394 <= 1'b0;
        pong_storage_data_394 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                259 / IN_WIDTH: ping_storage_data_394 <= (fillup_transition == 1'b1) ? i_input_data[259 % IN_WIDTH] : ping_storage_data_394 ^ i_input_data[259 % IN_WIDTH];
                598 / IN_WIDTH: ping_storage_data_394 <= (fillup_transition == 1'b1) ? i_input_data[598 % IN_WIDTH] : ping_storage_data_394 ^ i_input_data[598 % IN_WIDTH];
                929 / IN_WIDTH: ping_storage_data_394 <= (fillup_transition == 1'b1) ? i_input_data[929 % IN_WIDTH] : ping_storage_data_394 ^ i_input_data[929 % IN_WIDTH];
                994 / IN_WIDTH: ping_storage_data_394 <= (fillup_transition == 1'b1) ? i_input_data[994 % IN_WIDTH] : ping_storage_data_394 ^ i_input_data[994 % IN_WIDTH];
                default: ping_storage_data_394 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_394;
                endcase
            end else begin
                case (input_count)
                259 / IN_WIDTH: pong_storage_data_394 <= (fillup_transition == 1'b1) ? i_input_data[259 % IN_WIDTH] : pong_storage_data_394 ^ i_input_data[259 % IN_WIDTH];
                598 / IN_WIDTH: pong_storage_data_394 <= (fillup_transition == 1'b1) ? i_input_data[598 % IN_WIDTH] : pong_storage_data_394 ^ i_input_data[598 % IN_WIDTH];
                929 / IN_WIDTH: pong_storage_data_394 <= (fillup_transition == 1'b1) ? i_input_data[929 % IN_WIDTH] : pong_storage_data_394 ^ i_input_data[929 % IN_WIDTH];
                994 / IN_WIDTH: pong_storage_data_394 <= (fillup_transition == 1'b1) ? i_input_data[994 % IN_WIDTH] : pong_storage_data_394 ^ i_input_data[994 % IN_WIDTH];
                default: pong_storage_data_394 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_394;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_394 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_394;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_394 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_394;
            end
        end
    end
end

logic ping_storage_data_395;
logic pong_storage_data_395;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_395 <= 1'b0;
        pong_storage_data_395 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                260 / IN_WIDTH: ping_storage_data_395 <= (fillup_transition == 1'b1) ? i_input_data[260 % IN_WIDTH] : ping_storage_data_395 ^ i_input_data[260 % IN_WIDTH];
                599 / IN_WIDTH: ping_storage_data_395 <= (fillup_transition == 1'b1) ? i_input_data[599 % IN_WIDTH] : ping_storage_data_395 ^ i_input_data[599 % IN_WIDTH];
                930 / IN_WIDTH: ping_storage_data_395 <= (fillup_transition == 1'b1) ? i_input_data[930 % IN_WIDTH] : ping_storage_data_395 ^ i_input_data[930 % IN_WIDTH];
                995 / IN_WIDTH: ping_storage_data_395 <= (fillup_transition == 1'b1) ? i_input_data[995 % IN_WIDTH] : ping_storage_data_395 ^ i_input_data[995 % IN_WIDTH];
                default: ping_storage_data_395 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_395;
                endcase
            end else begin
                case (input_count)
                260 / IN_WIDTH: pong_storage_data_395 <= (fillup_transition == 1'b1) ? i_input_data[260 % IN_WIDTH] : pong_storage_data_395 ^ i_input_data[260 % IN_WIDTH];
                599 / IN_WIDTH: pong_storage_data_395 <= (fillup_transition == 1'b1) ? i_input_data[599 % IN_WIDTH] : pong_storage_data_395 ^ i_input_data[599 % IN_WIDTH];
                930 / IN_WIDTH: pong_storage_data_395 <= (fillup_transition == 1'b1) ? i_input_data[930 % IN_WIDTH] : pong_storage_data_395 ^ i_input_data[930 % IN_WIDTH];
                995 / IN_WIDTH: pong_storage_data_395 <= (fillup_transition == 1'b1) ? i_input_data[995 % IN_WIDTH] : pong_storage_data_395 ^ i_input_data[995 % IN_WIDTH];
                default: pong_storage_data_395 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_395;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_395 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_395;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_395 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_395;
            end
        end
    end
end

logic ping_storage_data_396;
logic pong_storage_data_396;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_396 <= 1'b0;
        pong_storage_data_396 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                261 / IN_WIDTH: ping_storage_data_396 <= (fillup_transition == 1'b1) ? i_input_data[261 % IN_WIDTH] : ping_storage_data_396 ^ i_input_data[261 % IN_WIDTH];
                600 / IN_WIDTH: ping_storage_data_396 <= (fillup_transition == 1'b1) ? i_input_data[600 % IN_WIDTH] : ping_storage_data_396 ^ i_input_data[600 % IN_WIDTH];
                931 / IN_WIDTH: ping_storage_data_396 <= (fillup_transition == 1'b1) ? i_input_data[931 % IN_WIDTH] : ping_storage_data_396 ^ i_input_data[931 % IN_WIDTH];
                996 / IN_WIDTH: ping_storage_data_396 <= (fillup_transition == 1'b1) ? i_input_data[996 % IN_WIDTH] : ping_storage_data_396 ^ i_input_data[996 % IN_WIDTH];
                default: ping_storage_data_396 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_396;
                endcase
            end else begin
                case (input_count)
                261 / IN_WIDTH: pong_storage_data_396 <= (fillup_transition == 1'b1) ? i_input_data[261 % IN_WIDTH] : pong_storage_data_396 ^ i_input_data[261 % IN_WIDTH];
                600 / IN_WIDTH: pong_storage_data_396 <= (fillup_transition == 1'b1) ? i_input_data[600 % IN_WIDTH] : pong_storage_data_396 ^ i_input_data[600 % IN_WIDTH];
                931 / IN_WIDTH: pong_storage_data_396 <= (fillup_transition == 1'b1) ? i_input_data[931 % IN_WIDTH] : pong_storage_data_396 ^ i_input_data[931 % IN_WIDTH];
                996 / IN_WIDTH: pong_storage_data_396 <= (fillup_transition == 1'b1) ? i_input_data[996 % IN_WIDTH] : pong_storage_data_396 ^ i_input_data[996 % IN_WIDTH];
                default: pong_storage_data_396 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_396;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_396 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_396;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_396 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_396;
            end
        end
    end
end

logic ping_storage_data_397;
logic pong_storage_data_397;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_397 <= 1'b0;
        pong_storage_data_397 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                262 / IN_WIDTH: ping_storage_data_397 <= (fillup_transition == 1'b1) ? i_input_data[262 % IN_WIDTH] : ping_storage_data_397 ^ i_input_data[262 % IN_WIDTH];
                601 / IN_WIDTH: ping_storage_data_397 <= (fillup_transition == 1'b1) ? i_input_data[601 % IN_WIDTH] : ping_storage_data_397 ^ i_input_data[601 % IN_WIDTH];
                932 / IN_WIDTH: ping_storage_data_397 <= (fillup_transition == 1'b1) ? i_input_data[932 % IN_WIDTH] : ping_storage_data_397 ^ i_input_data[932 % IN_WIDTH];
                997 / IN_WIDTH: ping_storage_data_397 <= (fillup_transition == 1'b1) ? i_input_data[997 % IN_WIDTH] : ping_storage_data_397 ^ i_input_data[997 % IN_WIDTH];
                default: ping_storage_data_397 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_397;
                endcase
            end else begin
                case (input_count)
                262 / IN_WIDTH: pong_storage_data_397 <= (fillup_transition == 1'b1) ? i_input_data[262 % IN_WIDTH] : pong_storage_data_397 ^ i_input_data[262 % IN_WIDTH];
                601 / IN_WIDTH: pong_storage_data_397 <= (fillup_transition == 1'b1) ? i_input_data[601 % IN_WIDTH] : pong_storage_data_397 ^ i_input_data[601 % IN_WIDTH];
                932 / IN_WIDTH: pong_storage_data_397 <= (fillup_transition == 1'b1) ? i_input_data[932 % IN_WIDTH] : pong_storage_data_397 ^ i_input_data[932 % IN_WIDTH];
                997 / IN_WIDTH: pong_storage_data_397 <= (fillup_transition == 1'b1) ? i_input_data[997 % IN_WIDTH] : pong_storage_data_397 ^ i_input_data[997 % IN_WIDTH];
                default: pong_storage_data_397 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_397;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_397 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_397;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_397 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_397;
            end
        end
    end
end

logic ping_storage_data_398;
logic pong_storage_data_398;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_398 <= 1'b0;
        pong_storage_data_398 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                263 / IN_WIDTH: ping_storage_data_398 <= (fillup_transition == 1'b1) ? i_input_data[263 % IN_WIDTH] : ping_storage_data_398 ^ i_input_data[263 % IN_WIDTH];
                602 / IN_WIDTH: ping_storage_data_398 <= (fillup_transition == 1'b1) ? i_input_data[602 % IN_WIDTH] : ping_storage_data_398 ^ i_input_data[602 % IN_WIDTH];
                933 / IN_WIDTH: ping_storage_data_398 <= (fillup_transition == 1'b1) ? i_input_data[933 % IN_WIDTH] : ping_storage_data_398 ^ i_input_data[933 % IN_WIDTH];
                998 / IN_WIDTH: ping_storage_data_398 <= (fillup_transition == 1'b1) ? i_input_data[998 % IN_WIDTH] : ping_storage_data_398 ^ i_input_data[998 % IN_WIDTH];
                default: ping_storage_data_398 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_398;
                endcase
            end else begin
                case (input_count)
                263 / IN_WIDTH: pong_storage_data_398 <= (fillup_transition == 1'b1) ? i_input_data[263 % IN_WIDTH] : pong_storage_data_398 ^ i_input_data[263 % IN_WIDTH];
                602 / IN_WIDTH: pong_storage_data_398 <= (fillup_transition == 1'b1) ? i_input_data[602 % IN_WIDTH] : pong_storage_data_398 ^ i_input_data[602 % IN_WIDTH];
                933 / IN_WIDTH: pong_storage_data_398 <= (fillup_transition == 1'b1) ? i_input_data[933 % IN_WIDTH] : pong_storage_data_398 ^ i_input_data[933 % IN_WIDTH];
                998 / IN_WIDTH: pong_storage_data_398 <= (fillup_transition == 1'b1) ? i_input_data[998 % IN_WIDTH] : pong_storage_data_398 ^ i_input_data[998 % IN_WIDTH];
                default: pong_storage_data_398 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_398;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_398 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_398;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_398 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_398;
            end
        end
    end
end

logic ping_storage_data_399;
logic pong_storage_data_399;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_399 <= 1'b0;
        pong_storage_data_399 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                264 / IN_WIDTH: ping_storage_data_399 <= (fillup_transition == 1'b1) ? i_input_data[264 % IN_WIDTH] : ping_storage_data_399 ^ i_input_data[264 % IN_WIDTH];
                603 / IN_WIDTH: ping_storage_data_399 <= (fillup_transition == 1'b1) ? i_input_data[603 % IN_WIDTH] : ping_storage_data_399 ^ i_input_data[603 % IN_WIDTH];
                934 / IN_WIDTH: ping_storage_data_399 <= (fillup_transition == 1'b1) ? i_input_data[934 % IN_WIDTH] : ping_storage_data_399 ^ i_input_data[934 % IN_WIDTH];
                999 / IN_WIDTH: ping_storage_data_399 <= (fillup_transition == 1'b1) ? i_input_data[999 % IN_WIDTH] : ping_storage_data_399 ^ i_input_data[999 % IN_WIDTH];
                default: ping_storage_data_399 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_399;
                endcase
            end else begin
                case (input_count)
                264 / IN_WIDTH: pong_storage_data_399 <= (fillup_transition == 1'b1) ? i_input_data[264 % IN_WIDTH] : pong_storage_data_399 ^ i_input_data[264 % IN_WIDTH];
                603 / IN_WIDTH: pong_storage_data_399 <= (fillup_transition == 1'b1) ? i_input_data[603 % IN_WIDTH] : pong_storage_data_399 ^ i_input_data[603 % IN_WIDTH];
                934 / IN_WIDTH: pong_storage_data_399 <= (fillup_transition == 1'b1) ? i_input_data[934 % IN_WIDTH] : pong_storage_data_399 ^ i_input_data[934 % IN_WIDTH];
                999 / IN_WIDTH: pong_storage_data_399 <= (fillup_transition == 1'b1) ? i_input_data[999 % IN_WIDTH] : pong_storage_data_399 ^ i_input_data[999 % IN_WIDTH];
                default: pong_storage_data_399 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_399;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_399 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_399;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_399 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_399;
            end
        end
    end
end

logic ping_storage_data_400;
logic pong_storage_data_400;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_400 <= 1'b0;
        pong_storage_data_400 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                265 / IN_WIDTH: ping_storage_data_400 <= (fillup_transition == 1'b1) ? i_input_data[265 % IN_WIDTH] : ping_storage_data_400 ^ i_input_data[265 % IN_WIDTH];
                604 / IN_WIDTH: ping_storage_data_400 <= (fillup_transition == 1'b1) ? i_input_data[604 % IN_WIDTH] : ping_storage_data_400 ^ i_input_data[604 % IN_WIDTH];
                935 / IN_WIDTH: ping_storage_data_400 <= (fillup_transition == 1'b1) ? i_input_data[935 % IN_WIDTH] : ping_storage_data_400 ^ i_input_data[935 % IN_WIDTH];
                1000 / IN_WIDTH: ping_storage_data_400 <= (fillup_transition == 1'b1) ? i_input_data[1000 % IN_WIDTH] : ping_storage_data_400 ^ i_input_data[1000 % IN_WIDTH];
                default: ping_storage_data_400 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_400;
                endcase
            end else begin
                case (input_count)
                265 / IN_WIDTH: pong_storage_data_400 <= (fillup_transition == 1'b1) ? i_input_data[265 % IN_WIDTH] : pong_storage_data_400 ^ i_input_data[265 % IN_WIDTH];
                604 / IN_WIDTH: pong_storage_data_400 <= (fillup_transition == 1'b1) ? i_input_data[604 % IN_WIDTH] : pong_storage_data_400 ^ i_input_data[604 % IN_WIDTH];
                935 / IN_WIDTH: pong_storage_data_400 <= (fillup_transition == 1'b1) ? i_input_data[935 % IN_WIDTH] : pong_storage_data_400 ^ i_input_data[935 % IN_WIDTH];
                1000 / IN_WIDTH: pong_storage_data_400 <= (fillup_transition == 1'b1) ? i_input_data[1000 % IN_WIDTH] : pong_storage_data_400 ^ i_input_data[1000 % IN_WIDTH];
                default: pong_storage_data_400 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_400;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_400 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_400;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_400 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_400;
            end
        end
    end
end

logic ping_storage_data_401;
logic pong_storage_data_401;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_401 <= 1'b0;
        pong_storage_data_401 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                266 / IN_WIDTH: ping_storage_data_401 <= (fillup_transition == 1'b1) ? i_input_data[266 % IN_WIDTH] : ping_storage_data_401 ^ i_input_data[266 % IN_WIDTH];
                605 / IN_WIDTH: ping_storage_data_401 <= (fillup_transition == 1'b1) ? i_input_data[605 % IN_WIDTH] : ping_storage_data_401 ^ i_input_data[605 % IN_WIDTH];
                936 / IN_WIDTH: ping_storage_data_401 <= (fillup_transition == 1'b1) ? i_input_data[936 % IN_WIDTH] : ping_storage_data_401 ^ i_input_data[936 % IN_WIDTH];
                1001 / IN_WIDTH: ping_storage_data_401 <= (fillup_transition == 1'b1) ? i_input_data[1001 % IN_WIDTH] : ping_storage_data_401 ^ i_input_data[1001 % IN_WIDTH];
                default: ping_storage_data_401 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_401;
                endcase
            end else begin
                case (input_count)
                266 / IN_WIDTH: pong_storage_data_401 <= (fillup_transition == 1'b1) ? i_input_data[266 % IN_WIDTH] : pong_storage_data_401 ^ i_input_data[266 % IN_WIDTH];
                605 / IN_WIDTH: pong_storage_data_401 <= (fillup_transition == 1'b1) ? i_input_data[605 % IN_WIDTH] : pong_storage_data_401 ^ i_input_data[605 % IN_WIDTH];
                936 / IN_WIDTH: pong_storage_data_401 <= (fillup_transition == 1'b1) ? i_input_data[936 % IN_WIDTH] : pong_storage_data_401 ^ i_input_data[936 % IN_WIDTH];
                1001 / IN_WIDTH: pong_storage_data_401 <= (fillup_transition == 1'b1) ? i_input_data[1001 % IN_WIDTH] : pong_storage_data_401 ^ i_input_data[1001 % IN_WIDTH];
                default: pong_storage_data_401 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_401;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_401 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_401;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_401 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_401;
            end
        end
    end
end

logic ping_storage_data_402;
logic pong_storage_data_402;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_402 <= 1'b0;
        pong_storage_data_402 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                267 / IN_WIDTH: ping_storage_data_402 <= (fillup_transition == 1'b1) ? i_input_data[267 % IN_WIDTH] : ping_storage_data_402 ^ i_input_data[267 % IN_WIDTH];
                606 / IN_WIDTH: ping_storage_data_402 <= (fillup_transition == 1'b1) ? i_input_data[606 % IN_WIDTH] : ping_storage_data_402 ^ i_input_data[606 % IN_WIDTH];
                937 / IN_WIDTH: ping_storage_data_402 <= (fillup_transition == 1'b1) ? i_input_data[937 % IN_WIDTH] : ping_storage_data_402 ^ i_input_data[937 % IN_WIDTH];
                1002 / IN_WIDTH: ping_storage_data_402 <= (fillup_transition == 1'b1) ? i_input_data[1002 % IN_WIDTH] : ping_storage_data_402 ^ i_input_data[1002 % IN_WIDTH];
                default: ping_storage_data_402 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_402;
                endcase
            end else begin
                case (input_count)
                267 / IN_WIDTH: pong_storage_data_402 <= (fillup_transition == 1'b1) ? i_input_data[267 % IN_WIDTH] : pong_storage_data_402 ^ i_input_data[267 % IN_WIDTH];
                606 / IN_WIDTH: pong_storage_data_402 <= (fillup_transition == 1'b1) ? i_input_data[606 % IN_WIDTH] : pong_storage_data_402 ^ i_input_data[606 % IN_WIDTH];
                937 / IN_WIDTH: pong_storage_data_402 <= (fillup_transition == 1'b1) ? i_input_data[937 % IN_WIDTH] : pong_storage_data_402 ^ i_input_data[937 % IN_WIDTH];
                1002 / IN_WIDTH: pong_storage_data_402 <= (fillup_transition == 1'b1) ? i_input_data[1002 % IN_WIDTH] : pong_storage_data_402 ^ i_input_data[1002 % IN_WIDTH];
                default: pong_storage_data_402 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_402;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_402 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_402;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_402 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_402;
            end
        end
    end
end

logic ping_storage_data_403;
logic pong_storage_data_403;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_403 <= 1'b0;
        pong_storage_data_403 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                268 / IN_WIDTH: ping_storage_data_403 <= (fillup_transition == 1'b1) ? i_input_data[268 % IN_WIDTH] : ping_storage_data_403 ^ i_input_data[268 % IN_WIDTH];
                607 / IN_WIDTH: ping_storage_data_403 <= (fillup_transition == 1'b1) ? i_input_data[607 % IN_WIDTH] : ping_storage_data_403 ^ i_input_data[607 % IN_WIDTH];
                938 / IN_WIDTH: ping_storage_data_403 <= (fillup_transition == 1'b1) ? i_input_data[938 % IN_WIDTH] : ping_storage_data_403 ^ i_input_data[938 % IN_WIDTH];
                1003 / IN_WIDTH: ping_storage_data_403 <= (fillup_transition == 1'b1) ? i_input_data[1003 % IN_WIDTH] : ping_storage_data_403 ^ i_input_data[1003 % IN_WIDTH];
                default: ping_storage_data_403 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_403;
                endcase
            end else begin
                case (input_count)
                268 / IN_WIDTH: pong_storage_data_403 <= (fillup_transition == 1'b1) ? i_input_data[268 % IN_WIDTH] : pong_storage_data_403 ^ i_input_data[268 % IN_WIDTH];
                607 / IN_WIDTH: pong_storage_data_403 <= (fillup_transition == 1'b1) ? i_input_data[607 % IN_WIDTH] : pong_storage_data_403 ^ i_input_data[607 % IN_WIDTH];
                938 / IN_WIDTH: pong_storage_data_403 <= (fillup_transition == 1'b1) ? i_input_data[938 % IN_WIDTH] : pong_storage_data_403 ^ i_input_data[938 % IN_WIDTH];
                1003 / IN_WIDTH: pong_storage_data_403 <= (fillup_transition == 1'b1) ? i_input_data[1003 % IN_WIDTH] : pong_storage_data_403 ^ i_input_data[1003 % IN_WIDTH];
                default: pong_storage_data_403 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_403;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_403 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_403;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_403 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_403;
            end
        end
    end
end

logic ping_storage_data_404;
logic pong_storage_data_404;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_404 <= 1'b0;
        pong_storage_data_404 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                269 / IN_WIDTH: ping_storage_data_404 <= (fillup_transition == 1'b1) ? i_input_data[269 % IN_WIDTH] : ping_storage_data_404 ^ i_input_data[269 % IN_WIDTH];
                608 / IN_WIDTH: ping_storage_data_404 <= (fillup_transition == 1'b1) ? i_input_data[608 % IN_WIDTH] : ping_storage_data_404 ^ i_input_data[608 % IN_WIDTH];
                939 / IN_WIDTH: ping_storage_data_404 <= (fillup_transition == 1'b1) ? i_input_data[939 % IN_WIDTH] : ping_storage_data_404 ^ i_input_data[939 % IN_WIDTH];
                1004 / IN_WIDTH: ping_storage_data_404 <= (fillup_transition == 1'b1) ? i_input_data[1004 % IN_WIDTH] : ping_storage_data_404 ^ i_input_data[1004 % IN_WIDTH];
                default: ping_storage_data_404 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_404;
                endcase
            end else begin
                case (input_count)
                269 / IN_WIDTH: pong_storage_data_404 <= (fillup_transition == 1'b1) ? i_input_data[269 % IN_WIDTH] : pong_storage_data_404 ^ i_input_data[269 % IN_WIDTH];
                608 / IN_WIDTH: pong_storage_data_404 <= (fillup_transition == 1'b1) ? i_input_data[608 % IN_WIDTH] : pong_storage_data_404 ^ i_input_data[608 % IN_WIDTH];
                939 / IN_WIDTH: pong_storage_data_404 <= (fillup_transition == 1'b1) ? i_input_data[939 % IN_WIDTH] : pong_storage_data_404 ^ i_input_data[939 % IN_WIDTH];
                1004 / IN_WIDTH: pong_storage_data_404 <= (fillup_transition == 1'b1) ? i_input_data[1004 % IN_WIDTH] : pong_storage_data_404 ^ i_input_data[1004 % IN_WIDTH];
                default: pong_storage_data_404 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_404;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_404 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_404;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_404 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_404;
            end
        end
    end
end

logic ping_storage_data_405;
logic pong_storage_data_405;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_405 <= 1'b0;
        pong_storage_data_405 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                270 / IN_WIDTH: ping_storage_data_405 <= (fillup_transition == 1'b1) ? i_input_data[270 % IN_WIDTH] : ping_storage_data_405 ^ i_input_data[270 % IN_WIDTH];
                609 / IN_WIDTH: ping_storage_data_405 <= (fillup_transition == 1'b1) ? i_input_data[609 % IN_WIDTH] : ping_storage_data_405 ^ i_input_data[609 % IN_WIDTH];
                940 / IN_WIDTH: ping_storage_data_405 <= (fillup_transition == 1'b1) ? i_input_data[940 % IN_WIDTH] : ping_storage_data_405 ^ i_input_data[940 % IN_WIDTH];
                1005 / IN_WIDTH: ping_storage_data_405 <= (fillup_transition == 1'b1) ? i_input_data[1005 % IN_WIDTH] : ping_storage_data_405 ^ i_input_data[1005 % IN_WIDTH];
                default: ping_storage_data_405 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_405;
                endcase
            end else begin
                case (input_count)
                270 / IN_WIDTH: pong_storage_data_405 <= (fillup_transition == 1'b1) ? i_input_data[270 % IN_WIDTH] : pong_storage_data_405 ^ i_input_data[270 % IN_WIDTH];
                609 / IN_WIDTH: pong_storage_data_405 <= (fillup_transition == 1'b1) ? i_input_data[609 % IN_WIDTH] : pong_storage_data_405 ^ i_input_data[609 % IN_WIDTH];
                940 / IN_WIDTH: pong_storage_data_405 <= (fillup_transition == 1'b1) ? i_input_data[940 % IN_WIDTH] : pong_storage_data_405 ^ i_input_data[940 % IN_WIDTH];
                1005 / IN_WIDTH: pong_storage_data_405 <= (fillup_transition == 1'b1) ? i_input_data[1005 % IN_WIDTH] : pong_storage_data_405 ^ i_input_data[1005 % IN_WIDTH];
                default: pong_storage_data_405 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_405;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_405 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_405;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_405 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_405;
            end
        end
    end
end

logic ping_storage_data_406;
logic pong_storage_data_406;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_406 <= 1'b0;
        pong_storage_data_406 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                271 / IN_WIDTH: ping_storage_data_406 <= (fillup_transition == 1'b1) ? i_input_data[271 % IN_WIDTH] : ping_storage_data_406 ^ i_input_data[271 % IN_WIDTH];
                610 / IN_WIDTH: ping_storage_data_406 <= (fillup_transition == 1'b1) ? i_input_data[610 % IN_WIDTH] : ping_storage_data_406 ^ i_input_data[610 % IN_WIDTH];
                941 / IN_WIDTH: ping_storage_data_406 <= (fillup_transition == 1'b1) ? i_input_data[941 % IN_WIDTH] : ping_storage_data_406 ^ i_input_data[941 % IN_WIDTH];
                1006 / IN_WIDTH: ping_storage_data_406 <= (fillup_transition == 1'b1) ? i_input_data[1006 % IN_WIDTH] : ping_storage_data_406 ^ i_input_data[1006 % IN_WIDTH];
                default: ping_storage_data_406 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_406;
                endcase
            end else begin
                case (input_count)
                271 / IN_WIDTH: pong_storage_data_406 <= (fillup_transition == 1'b1) ? i_input_data[271 % IN_WIDTH] : pong_storage_data_406 ^ i_input_data[271 % IN_WIDTH];
                610 / IN_WIDTH: pong_storage_data_406 <= (fillup_transition == 1'b1) ? i_input_data[610 % IN_WIDTH] : pong_storage_data_406 ^ i_input_data[610 % IN_WIDTH];
                941 / IN_WIDTH: pong_storage_data_406 <= (fillup_transition == 1'b1) ? i_input_data[941 % IN_WIDTH] : pong_storage_data_406 ^ i_input_data[941 % IN_WIDTH];
                1006 / IN_WIDTH: pong_storage_data_406 <= (fillup_transition == 1'b1) ? i_input_data[1006 % IN_WIDTH] : pong_storage_data_406 ^ i_input_data[1006 % IN_WIDTH];
                default: pong_storage_data_406 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_406;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_406 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_406;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_406 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_406;
            end
        end
    end
end

logic ping_storage_data_407;
logic pong_storage_data_407;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_407 <= 1'b0;
        pong_storage_data_407 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                272 / IN_WIDTH: ping_storage_data_407 <= (fillup_transition == 1'b1) ? i_input_data[272 % IN_WIDTH] : ping_storage_data_407 ^ i_input_data[272 % IN_WIDTH];
                611 / IN_WIDTH: ping_storage_data_407 <= (fillup_transition == 1'b1) ? i_input_data[611 % IN_WIDTH] : ping_storage_data_407 ^ i_input_data[611 % IN_WIDTH];
                942 / IN_WIDTH: ping_storage_data_407 <= (fillup_transition == 1'b1) ? i_input_data[942 % IN_WIDTH] : ping_storage_data_407 ^ i_input_data[942 % IN_WIDTH];
                1007 / IN_WIDTH: ping_storage_data_407 <= (fillup_transition == 1'b1) ? i_input_data[1007 % IN_WIDTH] : ping_storage_data_407 ^ i_input_data[1007 % IN_WIDTH];
                default: ping_storage_data_407 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_407;
                endcase
            end else begin
                case (input_count)
                272 / IN_WIDTH: pong_storage_data_407 <= (fillup_transition == 1'b1) ? i_input_data[272 % IN_WIDTH] : pong_storage_data_407 ^ i_input_data[272 % IN_WIDTH];
                611 / IN_WIDTH: pong_storage_data_407 <= (fillup_transition == 1'b1) ? i_input_data[611 % IN_WIDTH] : pong_storage_data_407 ^ i_input_data[611 % IN_WIDTH];
                942 / IN_WIDTH: pong_storage_data_407 <= (fillup_transition == 1'b1) ? i_input_data[942 % IN_WIDTH] : pong_storage_data_407 ^ i_input_data[942 % IN_WIDTH];
                1007 / IN_WIDTH: pong_storage_data_407 <= (fillup_transition == 1'b1) ? i_input_data[1007 % IN_WIDTH] : pong_storage_data_407 ^ i_input_data[1007 % IN_WIDTH];
                default: pong_storage_data_407 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_407;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_407 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_407;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_407 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_407;
            end
        end
    end
end

logic ping_storage_data_408;
logic pong_storage_data_408;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_408 <= 1'b0;
        pong_storage_data_408 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                273 / IN_WIDTH: ping_storage_data_408 <= (fillup_transition == 1'b1) ? i_input_data[273 % IN_WIDTH] : ping_storage_data_408 ^ i_input_data[273 % IN_WIDTH];
                612 / IN_WIDTH: ping_storage_data_408 <= (fillup_transition == 1'b1) ? i_input_data[612 % IN_WIDTH] : ping_storage_data_408 ^ i_input_data[612 % IN_WIDTH];
                943 / IN_WIDTH: ping_storage_data_408 <= (fillup_transition == 1'b1) ? i_input_data[943 % IN_WIDTH] : ping_storage_data_408 ^ i_input_data[943 % IN_WIDTH];
                1008 / IN_WIDTH: ping_storage_data_408 <= (fillup_transition == 1'b1) ? i_input_data[1008 % IN_WIDTH] : ping_storage_data_408 ^ i_input_data[1008 % IN_WIDTH];
                default: ping_storage_data_408 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_408;
                endcase
            end else begin
                case (input_count)
                273 / IN_WIDTH: pong_storage_data_408 <= (fillup_transition == 1'b1) ? i_input_data[273 % IN_WIDTH] : pong_storage_data_408 ^ i_input_data[273 % IN_WIDTH];
                612 / IN_WIDTH: pong_storage_data_408 <= (fillup_transition == 1'b1) ? i_input_data[612 % IN_WIDTH] : pong_storage_data_408 ^ i_input_data[612 % IN_WIDTH];
                943 / IN_WIDTH: pong_storage_data_408 <= (fillup_transition == 1'b1) ? i_input_data[943 % IN_WIDTH] : pong_storage_data_408 ^ i_input_data[943 % IN_WIDTH];
                1008 / IN_WIDTH: pong_storage_data_408 <= (fillup_transition == 1'b1) ? i_input_data[1008 % IN_WIDTH] : pong_storage_data_408 ^ i_input_data[1008 % IN_WIDTH];
                default: pong_storage_data_408 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_408;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_408 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_408;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_408 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_408;
            end
        end
    end
end

logic ping_storage_data_409;
logic pong_storage_data_409;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_409 <= 1'b0;
        pong_storage_data_409 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                274 / IN_WIDTH: ping_storage_data_409 <= (fillup_transition == 1'b1) ? i_input_data[274 % IN_WIDTH] : ping_storage_data_409 ^ i_input_data[274 % IN_WIDTH];
                613 / IN_WIDTH: ping_storage_data_409 <= (fillup_transition == 1'b1) ? i_input_data[613 % IN_WIDTH] : ping_storage_data_409 ^ i_input_data[613 % IN_WIDTH];
                944 / IN_WIDTH: ping_storage_data_409 <= (fillup_transition == 1'b1) ? i_input_data[944 % IN_WIDTH] : ping_storage_data_409 ^ i_input_data[944 % IN_WIDTH];
                1009 / IN_WIDTH: ping_storage_data_409 <= (fillup_transition == 1'b1) ? i_input_data[1009 % IN_WIDTH] : ping_storage_data_409 ^ i_input_data[1009 % IN_WIDTH];
                default: ping_storage_data_409 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_409;
                endcase
            end else begin
                case (input_count)
                274 / IN_WIDTH: pong_storage_data_409 <= (fillup_transition == 1'b1) ? i_input_data[274 % IN_WIDTH] : pong_storage_data_409 ^ i_input_data[274 % IN_WIDTH];
                613 / IN_WIDTH: pong_storage_data_409 <= (fillup_transition == 1'b1) ? i_input_data[613 % IN_WIDTH] : pong_storage_data_409 ^ i_input_data[613 % IN_WIDTH];
                944 / IN_WIDTH: pong_storage_data_409 <= (fillup_transition == 1'b1) ? i_input_data[944 % IN_WIDTH] : pong_storage_data_409 ^ i_input_data[944 % IN_WIDTH];
                1009 / IN_WIDTH: pong_storage_data_409 <= (fillup_transition == 1'b1) ? i_input_data[1009 % IN_WIDTH] : pong_storage_data_409 ^ i_input_data[1009 % IN_WIDTH];
                default: pong_storage_data_409 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_409;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_409 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_409;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_409 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_409;
            end
        end
    end
end

logic ping_storage_data_410;
logic pong_storage_data_410;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_410 <= 1'b0;
        pong_storage_data_410 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                275 / IN_WIDTH: ping_storage_data_410 <= (fillup_transition == 1'b1) ? i_input_data[275 % IN_WIDTH] : ping_storage_data_410 ^ i_input_data[275 % IN_WIDTH];
                614 / IN_WIDTH: ping_storage_data_410 <= (fillup_transition == 1'b1) ? i_input_data[614 % IN_WIDTH] : ping_storage_data_410 ^ i_input_data[614 % IN_WIDTH];
                945 / IN_WIDTH: ping_storage_data_410 <= (fillup_transition == 1'b1) ? i_input_data[945 % IN_WIDTH] : ping_storage_data_410 ^ i_input_data[945 % IN_WIDTH];
                1010 / IN_WIDTH: ping_storage_data_410 <= (fillup_transition == 1'b1) ? i_input_data[1010 % IN_WIDTH] : ping_storage_data_410 ^ i_input_data[1010 % IN_WIDTH];
                default: ping_storage_data_410 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_410;
                endcase
            end else begin
                case (input_count)
                275 / IN_WIDTH: pong_storage_data_410 <= (fillup_transition == 1'b1) ? i_input_data[275 % IN_WIDTH] : pong_storage_data_410 ^ i_input_data[275 % IN_WIDTH];
                614 / IN_WIDTH: pong_storage_data_410 <= (fillup_transition == 1'b1) ? i_input_data[614 % IN_WIDTH] : pong_storage_data_410 ^ i_input_data[614 % IN_WIDTH];
                945 / IN_WIDTH: pong_storage_data_410 <= (fillup_transition == 1'b1) ? i_input_data[945 % IN_WIDTH] : pong_storage_data_410 ^ i_input_data[945 % IN_WIDTH];
                1010 / IN_WIDTH: pong_storage_data_410 <= (fillup_transition == 1'b1) ? i_input_data[1010 % IN_WIDTH] : pong_storage_data_410 ^ i_input_data[1010 % IN_WIDTH];
                default: pong_storage_data_410 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_410;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_410 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_410;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_410 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_410;
            end
        end
    end
end

logic ping_storage_data_411;
logic pong_storage_data_411;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_411 <= 1'b0;
        pong_storage_data_411 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                276 / IN_WIDTH: ping_storage_data_411 <= (fillup_transition == 1'b1) ? i_input_data[276 % IN_WIDTH] : ping_storage_data_411 ^ i_input_data[276 % IN_WIDTH];
                615 / IN_WIDTH: ping_storage_data_411 <= (fillup_transition == 1'b1) ? i_input_data[615 % IN_WIDTH] : ping_storage_data_411 ^ i_input_data[615 % IN_WIDTH];
                946 / IN_WIDTH: ping_storage_data_411 <= (fillup_transition == 1'b1) ? i_input_data[946 % IN_WIDTH] : ping_storage_data_411 ^ i_input_data[946 % IN_WIDTH];
                1011 / IN_WIDTH: ping_storage_data_411 <= (fillup_transition == 1'b1) ? i_input_data[1011 % IN_WIDTH] : ping_storage_data_411 ^ i_input_data[1011 % IN_WIDTH];
                default: ping_storage_data_411 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_411;
                endcase
            end else begin
                case (input_count)
                276 / IN_WIDTH: pong_storage_data_411 <= (fillup_transition == 1'b1) ? i_input_data[276 % IN_WIDTH] : pong_storage_data_411 ^ i_input_data[276 % IN_WIDTH];
                615 / IN_WIDTH: pong_storage_data_411 <= (fillup_transition == 1'b1) ? i_input_data[615 % IN_WIDTH] : pong_storage_data_411 ^ i_input_data[615 % IN_WIDTH];
                946 / IN_WIDTH: pong_storage_data_411 <= (fillup_transition == 1'b1) ? i_input_data[946 % IN_WIDTH] : pong_storage_data_411 ^ i_input_data[946 % IN_WIDTH];
                1011 / IN_WIDTH: pong_storage_data_411 <= (fillup_transition == 1'b1) ? i_input_data[1011 % IN_WIDTH] : pong_storage_data_411 ^ i_input_data[1011 % IN_WIDTH];
                default: pong_storage_data_411 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_411;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_411 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_411;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_411 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_411;
            end
        end
    end
end

logic ping_storage_data_412;
logic pong_storage_data_412;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_412 <= 1'b0;
        pong_storage_data_412 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                277 / IN_WIDTH: ping_storage_data_412 <= (fillup_transition == 1'b1) ? i_input_data[277 % IN_WIDTH] : ping_storage_data_412 ^ i_input_data[277 % IN_WIDTH];
                616 / IN_WIDTH: ping_storage_data_412 <= (fillup_transition == 1'b1) ? i_input_data[616 % IN_WIDTH] : ping_storage_data_412 ^ i_input_data[616 % IN_WIDTH];
                947 / IN_WIDTH: ping_storage_data_412 <= (fillup_transition == 1'b1) ? i_input_data[947 % IN_WIDTH] : ping_storage_data_412 ^ i_input_data[947 % IN_WIDTH];
                1012 / IN_WIDTH: ping_storage_data_412 <= (fillup_transition == 1'b1) ? i_input_data[1012 % IN_WIDTH] : ping_storage_data_412 ^ i_input_data[1012 % IN_WIDTH];
                default: ping_storage_data_412 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_412;
                endcase
            end else begin
                case (input_count)
                277 / IN_WIDTH: pong_storage_data_412 <= (fillup_transition == 1'b1) ? i_input_data[277 % IN_WIDTH] : pong_storage_data_412 ^ i_input_data[277 % IN_WIDTH];
                616 / IN_WIDTH: pong_storage_data_412 <= (fillup_transition == 1'b1) ? i_input_data[616 % IN_WIDTH] : pong_storage_data_412 ^ i_input_data[616 % IN_WIDTH];
                947 / IN_WIDTH: pong_storage_data_412 <= (fillup_transition == 1'b1) ? i_input_data[947 % IN_WIDTH] : pong_storage_data_412 ^ i_input_data[947 % IN_WIDTH];
                1012 / IN_WIDTH: pong_storage_data_412 <= (fillup_transition == 1'b1) ? i_input_data[1012 % IN_WIDTH] : pong_storage_data_412 ^ i_input_data[1012 % IN_WIDTH];
                default: pong_storage_data_412 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_412;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_412 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_412;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_412 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_412;
            end
        end
    end
end

logic ping_storage_data_413;
logic pong_storage_data_413;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_413 <= 1'b0;
        pong_storage_data_413 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                278 / IN_WIDTH: ping_storage_data_413 <= (fillup_transition == 1'b1) ? i_input_data[278 % IN_WIDTH] : ping_storage_data_413 ^ i_input_data[278 % IN_WIDTH];
                617 / IN_WIDTH: ping_storage_data_413 <= (fillup_transition == 1'b1) ? i_input_data[617 % IN_WIDTH] : ping_storage_data_413 ^ i_input_data[617 % IN_WIDTH];
                948 / IN_WIDTH: ping_storage_data_413 <= (fillup_transition == 1'b1) ? i_input_data[948 % IN_WIDTH] : ping_storage_data_413 ^ i_input_data[948 % IN_WIDTH];
                1013 / IN_WIDTH: ping_storage_data_413 <= (fillup_transition == 1'b1) ? i_input_data[1013 % IN_WIDTH] : ping_storage_data_413 ^ i_input_data[1013 % IN_WIDTH];
                default: ping_storage_data_413 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_413;
                endcase
            end else begin
                case (input_count)
                278 / IN_WIDTH: pong_storage_data_413 <= (fillup_transition == 1'b1) ? i_input_data[278 % IN_WIDTH] : pong_storage_data_413 ^ i_input_data[278 % IN_WIDTH];
                617 / IN_WIDTH: pong_storage_data_413 <= (fillup_transition == 1'b1) ? i_input_data[617 % IN_WIDTH] : pong_storage_data_413 ^ i_input_data[617 % IN_WIDTH];
                948 / IN_WIDTH: pong_storage_data_413 <= (fillup_transition == 1'b1) ? i_input_data[948 % IN_WIDTH] : pong_storage_data_413 ^ i_input_data[948 % IN_WIDTH];
                1013 / IN_WIDTH: pong_storage_data_413 <= (fillup_transition == 1'b1) ? i_input_data[1013 % IN_WIDTH] : pong_storage_data_413 ^ i_input_data[1013 % IN_WIDTH];
                default: pong_storage_data_413 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_413;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_413 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_413;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_413 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_413;
            end
        end
    end
end

logic ping_storage_data_414;
logic pong_storage_data_414;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_414 <= 1'b0;
        pong_storage_data_414 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                279 / IN_WIDTH: ping_storage_data_414 <= (fillup_transition == 1'b1) ? i_input_data[279 % IN_WIDTH] : ping_storage_data_414 ^ i_input_data[279 % IN_WIDTH];
                618 / IN_WIDTH: ping_storage_data_414 <= (fillup_transition == 1'b1) ? i_input_data[618 % IN_WIDTH] : ping_storage_data_414 ^ i_input_data[618 % IN_WIDTH];
                949 / IN_WIDTH: ping_storage_data_414 <= (fillup_transition == 1'b1) ? i_input_data[949 % IN_WIDTH] : ping_storage_data_414 ^ i_input_data[949 % IN_WIDTH];
                1014 / IN_WIDTH: ping_storage_data_414 <= (fillup_transition == 1'b1) ? i_input_data[1014 % IN_WIDTH] : ping_storage_data_414 ^ i_input_data[1014 % IN_WIDTH];
                default: ping_storage_data_414 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_414;
                endcase
            end else begin
                case (input_count)
                279 / IN_WIDTH: pong_storage_data_414 <= (fillup_transition == 1'b1) ? i_input_data[279 % IN_WIDTH] : pong_storage_data_414 ^ i_input_data[279 % IN_WIDTH];
                618 / IN_WIDTH: pong_storage_data_414 <= (fillup_transition == 1'b1) ? i_input_data[618 % IN_WIDTH] : pong_storage_data_414 ^ i_input_data[618 % IN_WIDTH];
                949 / IN_WIDTH: pong_storage_data_414 <= (fillup_transition == 1'b1) ? i_input_data[949 % IN_WIDTH] : pong_storage_data_414 ^ i_input_data[949 % IN_WIDTH];
                1014 / IN_WIDTH: pong_storage_data_414 <= (fillup_transition == 1'b1) ? i_input_data[1014 % IN_WIDTH] : pong_storage_data_414 ^ i_input_data[1014 % IN_WIDTH];
                default: pong_storage_data_414 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_414;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_414 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_414;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_414 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_414;
            end
        end
    end
end

logic ping_storage_data_415;
logic pong_storage_data_415;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_415 <= 1'b0;
        pong_storage_data_415 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                280 / IN_WIDTH: ping_storage_data_415 <= (fillup_transition == 1'b1) ? i_input_data[280 % IN_WIDTH] : ping_storage_data_415 ^ i_input_data[280 % IN_WIDTH];
                619 / IN_WIDTH: ping_storage_data_415 <= (fillup_transition == 1'b1) ? i_input_data[619 % IN_WIDTH] : ping_storage_data_415 ^ i_input_data[619 % IN_WIDTH];
                950 / IN_WIDTH: ping_storage_data_415 <= (fillup_transition == 1'b1) ? i_input_data[950 % IN_WIDTH] : ping_storage_data_415 ^ i_input_data[950 % IN_WIDTH];
                1015 / IN_WIDTH: ping_storage_data_415 <= (fillup_transition == 1'b1) ? i_input_data[1015 % IN_WIDTH] : ping_storage_data_415 ^ i_input_data[1015 % IN_WIDTH];
                default: ping_storage_data_415 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_415;
                endcase
            end else begin
                case (input_count)
                280 / IN_WIDTH: pong_storage_data_415 <= (fillup_transition == 1'b1) ? i_input_data[280 % IN_WIDTH] : pong_storage_data_415 ^ i_input_data[280 % IN_WIDTH];
                619 / IN_WIDTH: pong_storage_data_415 <= (fillup_transition == 1'b1) ? i_input_data[619 % IN_WIDTH] : pong_storage_data_415 ^ i_input_data[619 % IN_WIDTH];
                950 / IN_WIDTH: pong_storage_data_415 <= (fillup_transition == 1'b1) ? i_input_data[950 % IN_WIDTH] : pong_storage_data_415 ^ i_input_data[950 % IN_WIDTH];
                1015 / IN_WIDTH: pong_storage_data_415 <= (fillup_transition == 1'b1) ? i_input_data[1015 % IN_WIDTH] : pong_storage_data_415 ^ i_input_data[1015 % IN_WIDTH];
                default: pong_storage_data_415 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_415;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_415 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_415;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_415 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_415;
            end
        end
    end
end

logic ping_storage_data_416;
logic pong_storage_data_416;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_416 <= 1'b0;
        pong_storage_data_416 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                281 / IN_WIDTH: ping_storage_data_416 <= (fillup_transition == 1'b1) ? i_input_data[281 % IN_WIDTH] : ping_storage_data_416 ^ i_input_data[281 % IN_WIDTH];
                620 / IN_WIDTH: ping_storage_data_416 <= (fillup_transition == 1'b1) ? i_input_data[620 % IN_WIDTH] : ping_storage_data_416 ^ i_input_data[620 % IN_WIDTH];
                951 / IN_WIDTH: ping_storage_data_416 <= (fillup_transition == 1'b1) ? i_input_data[951 % IN_WIDTH] : ping_storage_data_416 ^ i_input_data[951 % IN_WIDTH];
                1016 / IN_WIDTH: ping_storage_data_416 <= (fillup_transition == 1'b1) ? i_input_data[1016 % IN_WIDTH] : ping_storage_data_416 ^ i_input_data[1016 % IN_WIDTH];
                default: ping_storage_data_416 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_416;
                endcase
            end else begin
                case (input_count)
                281 / IN_WIDTH: pong_storage_data_416 <= (fillup_transition == 1'b1) ? i_input_data[281 % IN_WIDTH] : pong_storage_data_416 ^ i_input_data[281 % IN_WIDTH];
                620 / IN_WIDTH: pong_storage_data_416 <= (fillup_transition == 1'b1) ? i_input_data[620 % IN_WIDTH] : pong_storage_data_416 ^ i_input_data[620 % IN_WIDTH];
                951 / IN_WIDTH: pong_storage_data_416 <= (fillup_transition == 1'b1) ? i_input_data[951 % IN_WIDTH] : pong_storage_data_416 ^ i_input_data[951 % IN_WIDTH];
                1016 / IN_WIDTH: pong_storage_data_416 <= (fillup_transition == 1'b1) ? i_input_data[1016 % IN_WIDTH] : pong_storage_data_416 ^ i_input_data[1016 % IN_WIDTH];
                default: pong_storage_data_416 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_416;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_416 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_416;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_416 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_416;
            end
        end
    end
end

logic ping_storage_data_417;
logic pong_storage_data_417;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_417 <= 1'b0;
        pong_storage_data_417 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                282 / IN_WIDTH: ping_storage_data_417 <= (fillup_transition == 1'b1) ? i_input_data[282 % IN_WIDTH] : ping_storage_data_417 ^ i_input_data[282 % IN_WIDTH];
                621 / IN_WIDTH: ping_storage_data_417 <= (fillup_transition == 1'b1) ? i_input_data[621 % IN_WIDTH] : ping_storage_data_417 ^ i_input_data[621 % IN_WIDTH];
                952 / IN_WIDTH: ping_storage_data_417 <= (fillup_transition == 1'b1) ? i_input_data[952 % IN_WIDTH] : ping_storage_data_417 ^ i_input_data[952 % IN_WIDTH];
                1017 / IN_WIDTH: ping_storage_data_417 <= (fillup_transition == 1'b1) ? i_input_data[1017 % IN_WIDTH] : ping_storage_data_417 ^ i_input_data[1017 % IN_WIDTH];
                default: ping_storage_data_417 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_417;
                endcase
            end else begin
                case (input_count)
                282 / IN_WIDTH: pong_storage_data_417 <= (fillup_transition == 1'b1) ? i_input_data[282 % IN_WIDTH] : pong_storage_data_417 ^ i_input_data[282 % IN_WIDTH];
                621 / IN_WIDTH: pong_storage_data_417 <= (fillup_transition == 1'b1) ? i_input_data[621 % IN_WIDTH] : pong_storage_data_417 ^ i_input_data[621 % IN_WIDTH];
                952 / IN_WIDTH: pong_storage_data_417 <= (fillup_transition == 1'b1) ? i_input_data[952 % IN_WIDTH] : pong_storage_data_417 ^ i_input_data[952 % IN_WIDTH];
                1017 / IN_WIDTH: pong_storage_data_417 <= (fillup_transition == 1'b1) ? i_input_data[1017 % IN_WIDTH] : pong_storage_data_417 ^ i_input_data[1017 % IN_WIDTH];
                default: pong_storage_data_417 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_417;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_417 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_417;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_417 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_417;
            end
        end
    end
end

logic ping_storage_data_418;
logic pong_storage_data_418;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_418 <= 1'b0;
        pong_storage_data_418 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                283 / IN_WIDTH: ping_storage_data_418 <= (fillup_transition == 1'b1) ? i_input_data[283 % IN_WIDTH] : ping_storage_data_418 ^ i_input_data[283 % IN_WIDTH];
                622 / IN_WIDTH: ping_storage_data_418 <= (fillup_transition == 1'b1) ? i_input_data[622 % IN_WIDTH] : ping_storage_data_418 ^ i_input_data[622 % IN_WIDTH];
                953 / IN_WIDTH: ping_storage_data_418 <= (fillup_transition == 1'b1) ? i_input_data[953 % IN_WIDTH] : ping_storage_data_418 ^ i_input_data[953 % IN_WIDTH];
                1018 / IN_WIDTH: ping_storage_data_418 <= (fillup_transition == 1'b1) ? i_input_data[1018 % IN_WIDTH] : ping_storage_data_418 ^ i_input_data[1018 % IN_WIDTH];
                default: ping_storage_data_418 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_418;
                endcase
            end else begin
                case (input_count)
                283 / IN_WIDTH: pong_storage_data_418 <= (fillup_transition == 1'b1) ? i_input_data[283 % IN_WIDTH] : pong_storage_data_418 ^ i_input_data[283 % IN_WIDTH];
                622 / IN_WIDTH: pong_storage_data_418 <= (fillup_transition == 1'b1) ? i_input_data[622 % IN_WIDTH] : pong_storage_data_418 ^ i_input_data[622 % IN_WIDTH];
                953 / IN_WIDTH: pong_storage_data_418 <= (fillup_transition == 1'b1) ? i_input_data[953 % IN_WIDTH] : pong_storage_data_418 ^ i_input_data[953 % IN_WIDTH];
                1018 / IN_WIDTH: pong_storage_data_418 <= (fillup_transition == 1'b1) ? i_input_data[1018 % IN_WIDTH] : pong_storage_data_418 ^ i_input_data[1018 % IN_WIDTH];
                default: pong_storage_data_418 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_418;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_418 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_418;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_418 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_418;
            end
        end
    end
end

logic ping_storage_data_419;
logic pong_storage_data_419;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_419 <= 1'b0;
        pong_storage_data_419 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                284 / IN_WIDTH: ping_storage_data_419 <= (fillup_transition == 1'b1) ? i_input_data[284 % IN_WIDTH] : ping_storage_data_419 ^ i_input_data[284 % IN_WIDTH];
                623 / IN_WIDTH: ping_storage_data_419 <= (fillup_transition == 1'b1) ? i_input_data[623 % IN_WIDTH] : ping_storage_data_419 ^ i_input_data[623 % IN_WIDTH];
                954 / IN_WIDTH: ping_storage_data_419 <= (fillup_transition == 1'b1) ? i_input_data[954 % IN_WIDTH] : ping_storage_data_419 ^ i_input_data[954 % IN_WIDTH];
                1019 / IN_WIDTH: ping_storage_data_419 <= (fillup_transition == 1'b1) ? i_input_data[1019 % IN_WIDTH] : ping_storage_data_419 ^ i_input_data[1019 % IN_WIDTH];
                default: ping_storage_data_419 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_419;
                endcase
            end else begin
                case (input_count)
                284 / IN_WIDTH: pong_storage_data_419 <= (fillup_transition == 1'b1) ? i_input_data[284 % IN_WIDTH] : pong_storage_data_419 ^ i_input_data[284 % IN_WIDTH];
                623 / IN_WIDTH: pong_storage_data_419 <= (fillup_transition == 1'b1) ? i_input_data[623 % IN_WIDTH] : pong_storage_data_419 ^ i_input_data[623 % IN_WIDTH];
                954 / IN_WIDTH: pong_storage_data_419 <= (fillup_transition == 1'b1) ? i_input_data[954 % IN_WIDTH] : pong_storage_data_419 ^ i_input_data[954 % IN_WIDTH];
                1019 / IN_WIDTH: pong_storage_data_419 <= (fillup_transition == 1'b1) ? i_input_data[1019 % IN_WIDTH] : pong_storage_data_419 ^ i_input_data[1019 % IN_WIDTH];
                default: pong_storage_data_419 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_419;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_419 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_419;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_419 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_419;
            end
        end
    end
end

logic ping_storage_data_420;
logic pong_storage_data_420;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_420 <= 1'b0;
        pong_storage_data_420 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                285 / IN_WIDTH: ping_storage_data_420 <= (fillup_transition == 1'b1) ? i_input_data[285 % IN_WIDTH] : ping_storage_data_420 ^ i_input_data[285 % IN_WIDTH];
                624 / IN_WIDTH: ping_storage_data_420 <= (fillup_transition == 1'b1) ? i_input_data[624 % IN_WIDTH] : ping_storage_data_420 ^ i_input_data[624 % IN_WIDTH];
                955 / IN_WIDTH: ping_storage_data_420 <= (fillup_transition == 1'b1) ? i_input_data[955 % IN_WIDTH] : ping_storage_data_420 ^ i_input_data[955 % IN_WIDTH];
                1020 / IN_WIDTH: ping_storage_data_420 <= (fillup_transition == 1'b1) ? i_input_data[1020 % IN_WIDTH] : ping_storage_data_420 ^ i_input_data[1020 % IN_WIDTH];
                default: ping_storage_data_420 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_420;
                endcase
            end else begin
                case (input_count)
                285 / IN_WIDTH: pong_storage_data_420 <= (fillup_transition == 1'b1) ? i_input_data[285 % IN_WIDTH] : pong_storage_data_420 ^ i_input_data[285 % IN_WIDTH];
                624 / IN_WIDTH: pong_storage_data_420 <= (fillup_transition == 1'b1) ? i_input_data[624 % IN_WIDTH] : pong_storage_data_420 ^ i_input_data[624 % IN_WIDTH];
                955 / IN_WIDTH: pong_storage_data_420 <= (fillup_transition == 1'b1) ? i_input_data[955 % IN_WIDTH] : pong_storage_data_420 ^ i_input_data[955 % IN_WIDTH];
                1020 / IN_WIDTH: pong_storage_data_420 <= (fillup_transition == 1'b1) ? i_input_data[1020 % IN_WIDTH] : pong_storage_data_420 ^ i_input_data[1020 % IN_WIDTH];
                default: pong_storage_data_420 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_420;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_420 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_420;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_420 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_420;
            end
        end
    end
end

logic ping_storage_data_421;
logic pong_storage_data_421;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_421 <= 1'b0;
        pong_storage_data_421 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                286 / IN_WIDTH: ping_storage_data_421 <= (fillup_transition == 1'b1) ? i_input_data[286 % IN_WIDTH] : ping_storage_data_421 ^ i_input_data[286 % IN_WIDTH];
                625 / IN_WIDTH: ping_storage_data_421 <= (fillup_transition == 1'b1) ? i_input_data[625 % IN_WIDTH] : ping_storage_data_421 ^ i_input_data[625 % IN_WIDTH];
                956 / IN_WIDTH: ping_storage_data_421 <= (fillup_transition == 1'b1) ? i_input_data[956 % IN_WIDTH] : ping_storage_data_421 ^ i_input_data[956 % IN_WIDTH];
                1021 / IN_WIDTH: ping_storage_data_421 <= (fillup_transition == 1'b1) ? i_input_data[1021 % IN_WIDTH] : ping_storage_data_421 ^ i_input_data[1021 % IN_WIDTH];
                default: ping_storage_data_421 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_421;
                endcase
            end else begin
                case (input_count)
                286 / IN_WIDTH: pong_storage_data_421 <= (fillup_transition == 1'b1) ? i_input_data[286 % IN_WIDTH] : pong_storage_data_421 ^ i_input_data[286 % IN_WIDTH];
                625 / IN_WIDTH: pong_storage_data_421 <= (fillup_transition == 1'b1) ? i_input_data[625 % IN_WIDTH] : pong_storage_data_421 ^ i_input_data[625 % IN_WIDTH];
                956 / IN_WIDTH: pong_storage_data_421 <= (fillup_transition == 1'b1) ? i_input_data[956 % IN_WIDTH] : pong_storage_data_421 ^ i_input_data[956 % IN_WIDTH];
                1021 / IN_WIDTH: pong_storage_data_421 <= (fillup_transition == 1'b1) ? i_input_data[1021 % IN_WIDTH] : pong_storage_data_421 ^ i_input_data[1021 % IN_WIDTH];
                default: pong_storage_data_421 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_421;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_421 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_421;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_421 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_421;
            end
        end
    end
end

logic ping_storage_data_422;
logic pong_storage_data_422;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_422 <= 1'b0;
        pong_storage_data_422 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                287 / IN_WIDTH: ping_storage_data_422 <= (fillup_transition == 1'b1) ? i_input_data[287 % IN_WIDTH] : ping_storage_data_422 ^ i_input_data[287 % IN_WIDTH];
                626 / IN_WIDTH: ping_storage_data_422 <= (fillup_transition == 1'b1) ? i_input_data[626 % IN_WIDTH] : ping_storage_data_422 ^ i_input_data[626 % IN_WIDTH];
                957 / IN_WIDTH: ping_storage_data_422 <= (fillup_transition == 1'b1) ? i_input_data[957 % IN_WIDTH] : ping_storage_data_422 ^ i_input_data[957 % IN_WIDTH];
                1022 / IN_WIDTH: ping_storage_data_422 <= (fillup_transition == 1'b1) ? i_input_data[1022 % IN_WIDTH] : ping_storage_data_422 ^ i_input_data[1022 % IN_WIDTH];
                default: ping_storage_data_422 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_422;
                endcase
            end else begin
                case (input_count)
                287 / IN_WIDTH: pong_storage_data_422 <= (fillup_transition == 1'b1) ? i_input_data[287 % IN_WIDTH] : pong_storage_data_422 ^ i_input_data[287 % IN_WIDTH];
                626 / IN_WIDTH: pong_storage_data_422 <= (fillup_transition == 1'b1) ? i_input_data[626 % IN_WIDTH] : pong_storage_data_422 ^ i_input_data[626 % IN_WIDTH];
                957 / IN_WIDTH: pong_storage_data_422 <= (fillup_transition == 1'b1) ? i_input_data[957 % IN_WIDTH] : pong_storage_data_422 ^ i_input_data[957 % IN_WIDTH];
                1022 / IN_WIDTH: pong_storage_data_422 <= (fillup_transition == 1'b1) ? i_input_data[1022 % IN_WIDTH] : pong_storage_data_422 ^ i_input_data[1022 % IN_WIDTH];
                default: pong_storage_data_422 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_422;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_422 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_422;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_422 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_422;
            end
        end
    end
end

logic ping_storage_data_423;
logic pong_storage_data_423;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_423 <= 1'b0;
        pong_storage_data_423 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                192 / IN_WIDTH: ping_storage_data_423 <= (fillup_transition == 1'b1) ? i_input_data[192 % IN_WIDTH] : ping_storage_data_423 ^ i_input_data[192 % IN_WIDTH];
                627 / IN_WIDTH: ping_storage_data_423 <= (fillup_transition == 1'b1) ? i_input_data[627 % IN_WIDTH] : ping_storage_data_423 ^ i_input_data[627 % IN_WIDTH];
                958 / IN_WIDTH: ping_storage_data_423 <= (fillup_transition == 1'b1) ? i_input_data[958 % IN_WIDTH] : ping_storage_data_423 ^ i_input_data[958 % IN_WIDTH];
                1023 / IN_WIDTH: ping_storage_data_423 <= (fillup_transition == 1'b1) ? i_input_data[1023 % IN_WIDTH] : ping_storage_data_423 ^ i_input_data[1023 % IN_WIDTH];
                default: ping_storage_data_423 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_423;
                endcase
            end else begin
                case (input_count)
                192 / IN_WIDTH: pong_storage_data_423 <= (fillup_transition == 1'b1) ? i_input_data[192 % IN_WIDTH] : pong_storage_data_423 ^ i_input_data[192 % IN_WIDTH];
                627 / IN_WIDTH: pong_storage_data_423 <= (fillup_transition == 1'b1) ? i_input_data[627 % IN_WIDTH] : pong_storage_data_423 ^ i_input_data[627 % IN_WIDTH];
                958 / IN_WIDTH: pong_storage_data_423 <= (fillup_transition == 1'b1) ? i_input_data[958 % IN_WIDTH] : pong_storage_data_423 ^ i_input_data[958 % IN_WIDTH];
                1023 / IN_WIDTH: pong_storage_data_423 <= (fillup_transition == 1'b1) ? i_input_data[1023 % IN_WIDTH] : pong_storage_data_423 ^ i_input_data[1023 % IN_WIDTH];
                default: pong_storage_data_423 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_423;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_423 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_423;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_423 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_423;
            end
        end
    end
end

logic ping_storage_data_424;
logic pong_storage_data_424;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_424 <= 1'b0;
        pong_storage_data_424 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                193 / IN_WIDTH: ping_storage_data_424 <= (fillup_transition == 1'b1) ? i_input_data[193 % IN_WIDTH] : ping_storage_data_424 ^ i_input_data[193 % IN_WIDTH];
                628 / IN_WIDTH: ping_storage_data_424 <= (fillup_transition == 1'b1) ? i_input_data[628 % IN_WIDTH] : ping_storage_data_424 ^ i_input_data[628 % IN_WIDTH];
                959 / IN_WIDTH: ping_storage_data_424 <= (fillup_transition == 1'b1) ? i_input_data[959 % IN_WIDTH] : ping_storage_data_424 ^ i_input_data[959 % IN_WIDTH];
                1024 / IN_WIDTH: ping_storage_data_424 <= (fillup_transition == 1'b1) ? i_input_data[1024 % IN_WIDTH] : ping_storage_data_424 ^ i_input_data[1024 % IN_WIDTH];
                default: ping_storage_data_424 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_424;
                endcase
            end else begin
                case (input_count)
                193 / IN_WIDTH: pong_storage_data_424 <= (fillup_transition == 1'b1) ? i_input_data[193 % IN_WIDTH] : pong_storage_data_424 ^ i_input_data[193 % IN_WIDTH];
                628 / IN_WIDTH: pong_storage_data_424 <= (fillup_transition == 1'b1) ? i_input_data[628 % IN_WIDTH] : pong_storage_data_424 ^ i_input_data[628 % IN_WIDTH];
                959 / IN_WIDTH: pong_storage_data_424 <= (fillup_transition == 1'b1) ? i_input_data[959 % IN_WIDTH] : pong_storage_data_424 ^ i_input_data[959 % IN_WIDTH];
                1024 / IN_WIDTH: pong_storage_data_424 <= (fillup_transition == 1'b1) ? i_input_data[1024 % IN_WIDTH] : pong_storage_data_424 ^ i_input_data[1024 % IN_WIDTH];
                default: pong_storage_data_424 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_424;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_424 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_424;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_424 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_424;
            end
        end
    end
end

logic ping_storage_data_425;
logic pong_storage_data_425;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_425 <= 1'b0;
        pong_storage_data_425 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                194 / IN_WIDTH: ping_storage_data_425 <= (fillup_transition == 1'b1) ? i_input_data[194 % IN_WIDTH] : ping_storage_data_425 ^ i_input_data[194 % IN_WIDTH];
                629 / IN_WIDTH: ping_storage_data_425 <= (fillup_transition == 1'b1) ? i_input_data[629 % IN_WIDTH] : ping_storage_data_425 ^ i_input_data[629 % IN_WIDTH];
                864 / IN_WIDTH: ping_storage_data_425 <= (fillup_transition == 1'b1) ? i_input_data[864 % IN_WIDTH] : ping_storage_data_425 ^ i_input_data[864 % IN_WIDTH];
                1025 / IN_WIDTH: ping_storage_data_425 <= (fillup_transition == 1'b1) ? i_input_data[1025 % IN_WIDTH] : ping_storage_data_425 ^ i_input_data[1025 % IN_WIDTH];
                default: ping_storage_data_425 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_425;
                endcase
            end else begin
                case (input_count)
                194 / IN_WIDTH: pong_storage_data_425 <= (fillup_transition == 1'b1) ? i_input_data[194 % IN_WIDTH] : pong_storage_data_425 ^ i_input_data[194 % IN_WIDTH];
                629 / IN_WIDTH: pong_storage_data_425 <= (fillup_transition == 1'b1) ? i_input_data[629 % IN_WIDTH] : pong_storage_data_425 ^ i_input_data[629 % IN_WIDTH];
                864 / IN_WIDTH: pong_storage_data_425 <= (fillup_transition == 1'b1) ? i_input_data[864 % IN_WIDTH] : pong_storage_data_425 ^ i_input_data[864 % IN_WIDTH];
                1025 / IN_WIDTH: pong_storage_data_425 <= (fillup_transition == 1'b1) ? i_input_data[1025 % IN_WIDTH] : pong_storage_data_425 ^ i_input_data[1025 % IN_WIDTH];
                default: pong_storage_data_425 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_425;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_425 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_425;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_425 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_425;
            end
        end
    end
end

logic ping_storage_data_426;
logic pong_storage_data_426;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_426 <= 1'b0;
        pong_storage_data_426 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                195 / IN_WIDTH: ping_storage_data_426 <= (fillup_transition == 1'b1) ? i_input_data[195 % IN_WIDTH] : ping_storage_data_426 ^ i_input_data[195 % IN_WIDTH];
                630 / IN_WIDTH: ping_storage_data_426 <= (fillup_transition == 1'b1) ? i_input_data[630 % IN_WIDTH] : ping_storage_data_426 ^ i_input_data[630 % IN_WIDTH];
                865 / IN_WIDTH: ping_storage_data_426 <= (fillup_transition == 1'b1) ? i_input_data[865 % IN_WIDTH] : ping_storage_data_426 ^ i_input_data[865 % IN_WIDTH];
                1026 / IN_WIDTH: ping_storage_data_426 <= (fillup_transition == 1'b1) ? i_input_data[1026 % IN_WIDTH] : ping_storage_data_426 ^ i_input_data[1026 % IN_WIDTH];
                default: ping_storage_data_426 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_426;
                endcase
            end else begin
                case (input_count)
                195 / IN_WIDTH: pong_storage_data_426 <= (fillup_transition == 1'b1) ? i_input_data[195 % IN_WIDTH] : pong_storage_data_426 ^ i_input_data[195 % IN_WIDTH];
                630 / IN_WIDTH: pong_storage_data_426 <= (fillup_transition == 1'b1) ? i_input_data[630 % IN_WIDTH] : pong_storage_data_426 ^ i_input_data[630 % IN_WIDTH];
                865 / IN_WIDTH: pong_storage_data_426 <= (fillup_transition == 1'b1) ? i_input_data[865 % IN_WIDTH] : pong_storage_data_426 ^ i_input_data[865 % IN_WIDTH];
                1026 / IN_WIDTH: pong_storage_data_426 <= (fillup_transition == 1'b1) ? i_input_data[1026 % IN_WIDTH] : pong_storage_data_426 ^ i_input_data[1026 % IN_WIDTH];
                default: pong_storage_data_426 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_426;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_426 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_426;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_426 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_426;
            end
        end
    end
end

logic ping_storage_data_427;
logic pong_storage_data_427;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_427 <= 1'b0;
        pong_storage_data_427 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                196 / IN_WIDTH: ping_storage_data_427 <= (fillup_transition == 1'b1) ? i_input_data[196 % IN_WIDTH] : ping_storage_data_427 ^ i_input_data[196 % IN_WIDTH];
                631 / IN_WIDTH: ping_storage_data_427 <= (fillup_transition == 1'b1) ? i_input_data[631 % IN_WIDTH] : ping_storage_data_427 ^ i_input_data[631 % IN_WIDTH];
                866 / IN_WIDTH: ping_storage_data_427 <= (fillup_transition == 1'b1) ? i_input_data[866 % IN_WIDTH] : ping_storage_data_427 ^ i_input_data[866 % IN_WIDTH];
                1027 / IN_WIDTH: ping_storage_data_427 <= (fillup_transition == 1'b1) ? i_input_data[1027 % IN_WIDTH] : ping_storage_data_427 ^ i_input_data[1027 % IN_WIDTH];
                default: ping_storage_data_427 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_427;
                endcase
            end else begin
                case (input_count)
                196 / IN_WIDTH: pong_storage_data_427 <= (fillup_transition == 1'b1) ? i_input_data[196 % IN_WIDTH] : pong_storage_data_427 ^ i_input_data[196 % IN_WIDTH];
                631 / IN_WIDTH: pong_storage_data_427 <= (fillup_transition == 1'b1) ? i_input_data[631 % IN_WIDTH] : pong_storage_data_427 ^ i_input_data[631 % IN_WIDTH];
                866 / IN_WIDTH: pong_storage_data_427 <= (fillup_transition == 1'b1) ? i_input_data[866 % IN_WIDTH] : pong_storage_data_427 ^ i_input_data[866 % IN_WIDTH];
                1027 / IN_WIDTH: pong_storage_data_427 <= (fillup_transition == 1'b1) ? i_input_data[1027 % IN_WIDTH] : pong_storage_data_427 ^ i_input_data[1027 % IN_WIDTH];
                default: pong_storage_data_427 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_427;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_427 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_427;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_427 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_427;
            end
        end
    end
end

logic ping_storage_data_428;
logic pong_storage_data_428;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_428 <= 1'b0;
        pong_storage_data_428 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                197 / IN_WIDTH: ping_storage_data_428 <= (fillup_transition == 1'b1) ? i_input_data[197 % IN_WIDTH] : ping_storage_data_428 ^ i_input_data[197 % IN_WIDTH];
                632 / IN_WIDTH: ping_storage_data_428 <= (fillup_transition == 1'b1) ? i_input_data[632 % IN_WIDTH] : ping_storage_data_428 ^ i_input_data[632 % IN_WIDTH];
                867 / IN_WIDTH: ping_storage_data_428 <= (fillup_transition == 1'b1) ? i_input_data[867 % IN_WIDTH] : ping_storage_data_428 ^ i_input_data[867 % IN_WIDTH];
                1028 / IN_WIDTH: ping_storage_data_428 <= (fillup_transition == 1'b1) ? i_input_data[1028 % IN_WIDTH] : ping_storage_data_428 ^ i_input_data[1028 % IN_WIDTH];
                default: ping_storage_data_428 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_428;
                endcase
            end else begin
                case (input_count)
                197 / IN_WIDTH: pong_storage_data_428 <= (fillup_transition == 1'b1) ? i_input_data[197 % IN_WIDTH] : pong_storage_data_428 ^ i_input_data[197 % IN_WIDTH];
                632 / IN_WIDTH: pong_storage_data_428 <= (fillup_transition == 1'b1) ? i_input_data[632 % IN_WIDTH] : pong_storage_data_428 ^ i_input_data[632 % IN_WIDTH];
                867 / IN_WIDTH: pong_storage_data_428 <= (fillup_transition == 1'b1) ? i_input_data[867 % IN_WIDTH] : pong_storage_data_428 ^ i_input_data[867 % IN_WIDTH];
                1028 / IN_WIDTH: pong_storage_data_428 <= (fillup_transition == 1'b1) ? i_input_data[1028 % IN_WIDTH] : pong_storage_data_428 ^ i_input_data[1028 % IN_WIDTH];
                default: pong_storage_data_428 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_428;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_428 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_428;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_428 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_428;
            end
        end
    end
end

logic ping_storage_data_429;
logic pong_storage_data_429;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_429 <= 1'b0;
        pong_storage_data_429 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                198 / IN_WIDTH: ping_storage_data_429 <= (fillup_transition == 1'b1) ? i_input_data[198 % IN_WIDTH] : ping_storage_data_429 ^ i_input_data[198 % IN_WIDTH];
                633 / IN_WIDTH: ping_storage_data_429 <= (fillup_transition == 1'b1) ? i_input_data[633 % IN_WIDTH] : ping_storage_data_429 ^ i_input_data[633 % IN_WIDTH];
                868 / IN_WIDTH: ping_storage_data_429 <= (fillup_transition == 1'b1) ? i_input_data[868 % IN_WIDTH] : ping_storage_data_429 ^ i_input_data[868 % IN_WIDTH];
                1029 / IN_WIDTH: ping_storage_data_429 <= (fillup_transition == 1'b1) ? i_input_data[1029 % IN_WIDTH] : ping_storage_data_429 ^ i_input_data[1029 % IN_WIDTH];
                default: ping_storage_data_429 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_429;
                endcase
            end else begin
                case (input_count)
                198 / IN_WIDTH: pong_storage_data_429 <= (fillup_transition == 1'b1) ? i_input_data[198 % IN_WIDTH] : pong_storage_data_429 ^ i_input_data[198 % IN_WIDTH];
                633 / IN_WIDTH: pong_storage_data_429 <= (fillup_transition == 1'b1) ? i_input_data[633 % IN_WIDTH] : pong_storage_data_429 ^ i_input_data[633 % IN_WIDTH];
                868 / IN_WIDTH: pong_storage_data_429 <= (fillup_transition == 1'b1) ? i_input_data[868 % IN_WIDTH] : pong_storage_data_429 ^ i_input_data[868 % IN_WIDTH];
                1029 / IN_WIDTH: pong_storage_data_429 <= (fillup_transition == 1'b1) ? i_input_data[1029 % IN_WIDTH] : pong_storage_data_429 ^ i_input_data[1029 % IN_WIDTH];
                default: pong_storage_data_429 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_429;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_429 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_429;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_429 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_429;
            end
        end
    end
end

logic ping_storage_data_430;
logic pong_storage_data_430;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_430 <= 1'b0;
        pong_storage_data_430 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                199 / IN_WIDTH: ping_storage_data_430 <= (fillup_transition == 1'b1) ? i_input_data[199 % IN_WIDTH] : ping_storage_data_430 ^ i_input_data[199 % IN_WIDTH];
                634 / IN_WIDTH: ping_storage_data_430 <= (fillup_transition == 1'b1) ? i_input_data[634 % IN_WIDTH] : ping_storage_data_430 ^ i_input_data[634 % IN_WIDTH];
                869 / IN_WIDTH: ping_storage_data_430 <= (fillup_transition == 1'b1) ? i_input_data[869 % IN_WIDTH] : ping_storage_data_430 ^ i_input_data[869 % IN_WIDTH];
                1030 / IN_WIDTH: ping_storage_data_430 <= (fillup_transition == 1'b1) ? i_input_data[1030 % IN_WIDTH] : ping_storage_data_430 ^ i_input_data[1030 % IN_WIDTH];
                default: ping_storage_data_430 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_430;
                endcase
            end else begin
                case (input_count)
                199 / IN_WIDTH: pong_storage_data_430 <= (fillup_transition == 1'b1) ? i_input_data[199 % IN_WIDTH] : pong_storage_data_430 ^ i_input_data[199 % IN_WIDTH];
                634 / IN_WIDTH: pong_storage_data_430 <= (fillup_transition == 1'b1) ? i_input_data[634 % IN_WIDTH] : pong_storage_data_430 ^ i_input_data[634 % IN_WIDTH];
                869 / IN_WIDTH: pong_storage_data_430 <= (fillup_transition == 1'b1) ? i_input_data[869 % IN_WIDTH] : pong_storage_data_430 ^ i_input_data[869 % IN_WIDTH];
                1030 / IN_WIDTH: pong_storage_data_430 <= (fillup_transition == 1'b1) ? i_input_data[1030 % IN_WIDTH] : pong_storage_data_430 ^ i_input_data[1030 % IN_WIDTH];
                default: pong_storage_data_430 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_430;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_430 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_430;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_430 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_430;
            end
        end
    end
end

logic ping_storage_data_431;
logic pong_storage_data_431;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_431 <= 1'b0;
        pong_storage_data_431 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                200 / IN_WIDTH: ping_storage_data_431 <= (fillup_transition == 1'b1) ? i_input_data[200 % IN_WIDTH] : ping_storage_data_431 ^ i_input_data[200 % IN_WIDTH];
                635 / IN_WIDTH: ping_storage_data_431 <= (fillup_transition == 1'b1) ? i_input_data[635 % IN_WIDTH] : ping_storage_data_431 ^ i_input_data[635 % IN_WIDTH];
                870 / IN_WIDTH: ping_storage_data_431 <= (fillup_transition == 1'b1) ? i_input_data[870 % IN_WIDTH] : ping_storage_data_431 ^ i_input_data[870 % IN_WIDTH];
                1031 / IN_WIDTH: ping_storage_data_431 <= (fillup_transition == 1'b1) ? i_input_data[1031 % IN_WIDTH] : ping_storage_data_431 ^ i_input_data[1031 % IN_WIDTH];
                default: ping_storage_data_431 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_431;
                endcase
            end else begin
                case (input_count)
                200 / IN_WIDTH: pong_storage_data_431 <= (fillup_transition == 1'b1) ? i_input_data[200 % IN_WIDTH] : pong_storage_data_431 ^ i_input_data[200 % IN_WIDTH];
                635 / IN_WIDTH: pong_storage_data_431 <= (fillup_transition == 1'b1) ? i_input_data[635 % IN_WIDTH] : pong_storage_data_431 ^ i_input_data[635 % IN_WIDTH];
                870 / IN_WIDTH: pong_storage_data_431 <= (fillup_transition == 1'b1) ? i_input_data[870 % IN_WIDTH] : pong_storage_data_431 ^ i_input_data[870 % IN_WIDTH];
                1031 / IN_WIDTH: pong_storage_data_431 <= (fillup_transition == 1'b1) ? i_input_data[1031 % IN_WIDTH] : pong_storage_data_431 ^ i_input_data[1031 % IN_WIDTH];
                default: pong_storage_data_431 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_431;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_431 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_431;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_431 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_431;
            end
        end
    end
end

logic ping_storage_data_432;
logic pong_storage_data_432;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_432 <= 1'b0;
        pong_storage_data_432 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                201 / IN_WIDTH: ping_storage_data_432 <= (fillup_transition == 1'b1) ? i_input_data[201 % IN_WIDTH] : ping_storage_data_432 ^ i_input_data[201 % IN_WIDTH];
                636 / IN_WIDTH: ping_storage_data_432 <= (fillup_transition == 1'b1) ? i_input_data[636 % IN_WIDTH] : ping_storage_data_432 ^ i_input_data[636 % IN_WIDTH];
                871 / IN_WIDTH: ping_storage_data_432 <= (fillup_transition == 1'b1) ? i_input_data[871 % IN_WIDTH] : ping_storage_data_432 ^ i_input_data[871 % IN_WIDTH];
                1032 / IN_WIDTH: ping_storage_data_432 <= (fillup_transition == 1'b1) ? i_input_data[1032 % IN_WIDTH] : ping_storage_data_432 ^ i_input_data[1032 % IN_WIDTH];
                default: ping_storage_data_432 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_432;
                endcase
            end else begin
                case (input_count)
                201 / IN_WIDTH: pong_storage_data_432 <= (fillup_transition == 1'b1) ? i_input_data[201 % IN_WIDTH] : pong_storage_data_432 ^ i_input_data[201 % IN_WIDTH];
                636 / IN_WIDTH: pong_storage_data_432 <= (fillup_transition == 1'b1) ? i_input_data[636 % IN_WIDTH] : pong_storage_data_432 ^ i_input_data[636 % IN_WIDTH];
                871 / IN_WIDTH: pong_storage_data_432 <= (fillup_transition == 1'b1) ? i_input_data[871 % IN_WIDTH] : pong_storage_data_432 ^ i_input_data[871 % IN_WIDTH];
                1032 / IN_WIDTH: pong_storage_data_432 <= (fillup_transition == 1'b1) ? i_input_data[1032 % IN_WIDTH] : pong_storage_data_432 ^ i_input_data[1032 % IN_WIDTH];
                default: pong_storage_data_432 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_432;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_432 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_432;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_432 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_432;
            end
        end
    end
end

logic ping_storage_data_433;
logic pong_storage_data_433;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_433 <= 1'b0;
        pong_storage_data_433 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                202 / IN_WIDTH: ping_storage_data_433 <= (fillup_transition == 1'b1) ? i_input_data[202 % IN_WIDTH] : ping_storage_data_433 ^ i_input_data[202 % IN_WIDTH];
                637 / IN_WIDTH: ping_storage_data_433 <= (fillup_transition == 1'b1) ? i_input_data[637 % IN_WIDTH] : ping_storage_data_433 ^ i_input_data[637 % IN_WIDTH];
                872 / IN_WIDTH: ping_storage_data_433 <= (fillup_transition == 1'b1) ? i_input_data[872 % IN_WIDTH] : ping_storage_data_433 ^ i_input_data[872 % IN_WIDTH];
                1033 / IN_WIDTH: ping_storage_data_433 <= (fillup_transition == 1'b1) ? i_input_data[1033 % IN_WIDTH] : ping_storage_data_433 ^ i_input_data[1033 % IN_WIDTH];
                default: ping_storage_data_433 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_433;
                endcase
            end else begin
                case (input_count)
                202 / IN_WIDTH: pong_storage_data_433 <= (fillup_transition == 1'b1) ? i_input_data[202 % IN_WIDTH] : pong_storage_data_433 ^ i_input_data[202 % IN_WIDTH];
                637 / IN_WIDTH: pong_storage_data_433 <= (fillup_transition == 1'b1) ? i_input_data[637 % IN_WIDTH] : pong_storage_data_433 ^ i_input_data[637 % IN_WIDTH];
                872 / IN_WIDTH: pong_storage_data_433 <= (fillup_transition == 1'b1) ? i_input_data[872 % IN_WIDTH] : pong_storage_data_433 ^ i_input_data[872 % IN_WIDTH];
                1033 / IN_WIDTH: pong_storage_data_433 <= (fillup_transition == 1'b1) ? i_input_data[1033 % IN_WIDTH] : pong_storage_data_433 ^ i_input_data[1033 % IN_WIDTH];
                default: pong_storage_data_433 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_433;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_433 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_433;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_433 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_433;
            end
        end
    end
end

logic ping_storage_data_434;
logic pong_storage_data_434;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_434 <= 1'b0;
        pong_storage_data_434 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                203 / IN_WIDTH: ping_storage_data_434 <= (fillup_transition == 1'b1) ? i_input_data[203 % IN_WIDTH] : ping_storage_data_434 ^ i_input_data[203 % IN_WIDTH];
                638 / IN_WIDTH: ping_storage_data_434 <= (fillup_transition == 1'b1) ? i_input_data[638 % IN_WIDTH] : ping_storage_data_434 ^ i_input_data[638 % IN_WIDTH];
                873 / IN_WIDTH: ping_storage_data_434 <= (fillup_transition == 1'b1) ? i_input_data[873 % IN_WIDTH] : ping_storage_data_434 ^ i_input_data[873 % IN_WIDTH];
                1034 / IN_WIDTH: ping_storage_data_434 <= (fillup_transition == 1'b1) ? i_input_data[1034 % IN_WIDTH] : ping_storage_data_434 ^ i_input_data[1034 % IN_WIDTH];
                default: ping_storage_data_434 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_434;
                endcase
            end else begin
                case (input_count)
                203 / IN_WIDTH: pong_storage_data_434 <= (fillup_transition == 1'b1) ? i_input_data[203 % IN_WIDTH] : pong_storage_data_434 ^ i_input_data[203 % IN_WIDTH];
                638 / IN_WIDTH: pong_storage_data_434 <= (fillup_transition == 1'b1) ? i_input_data[638 % IN_WIDTH] : pong_storage_data_434 ^ i_input_data[638 % IN_WIDTH];
                873 / IN_WIDTH: pong_storage_data_434 <= (fillup_transition == 1'b1) ? i_input_data[873 % IN_WIDTH] : pong_storage_data_434 ^ i_input_data[873 % IN_WIDTH];
                1034 / IN_WIDTH: pong_storage_data_434 <= (fillup_transition == 1'b1) ? i_input_data[1034 % IN_WIDTH] : pong_storage_data_434 ^ i_input_data[1034 % IN_WIDTH];
                default: pong_storage_data_434 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_434;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_434 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_434;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_434 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_434;
            end
        end
    end
end

logic ping_storage_data_435;
logic pong_storage_data_435;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_435 <= 1'b0;
        pong_storage_data_435 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                204 / IN_WIDTH: ping_storage_data_435 <= (fillup_transition == 1'b1) ? i_input_data[204 % IN_WIDTH] : ping_storage_data_435 ^ i_input_data[204 % IN_WIDTH];
                639 / IN_WIDTH: ping_storage_data_435 <= (fillup_transition == 1'b1) ? i_input_data[639 % IN_WIDTH] : ping_storage_data_435 ^ i_input_data[639 % IN_WIDTH];
                874 / IN_WIDTH: ping_storage_data_435 <= (fillup_transition == 1'b1) ? i_input_data[874 % IN_WIDTH] : ping_storage_data_435 ^ i_input_data[874 % IN_WIDTH];
                1035 / IN_WIDTH: ping_storage_data_435 <= (fillup_transition == 1'b1) ? i_input_data[1035 % IN_WIDTH] : ping_storage_data_435 ^ i_input_data[1035 % IN_WIDTH];
                default: ping_storage_data_435 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_435;
                endcase
            end else begin
                case (input_count)
                204 / IN_WIDTH: pong_storage_data_435 <= (fillup_transition == 1'b1) ? i_input_data[204 % IN_WIDTH] : pong_storage_data_435 ^ i_input_data[204 % IN_WIDTH];
                639 / IN_WIDTH: pong_storage_data_435 <= (fillup_transition == 1'b1) ? i_input_data[639 % IN_WIDTH] : pong_storage_data_435 ^ i_input_data[639 % IN_WIDTH];
                874 / IN_WIDTH: pong_storage_data_435 <= (fillup_transition == 1'b1) ? i_input_data[874 % IN_WIDTH] : pong_storage_data_435 ^ i_input_data[874 % IN_WIDTH];
                1035 / IN_WIDTH: pong_storage_data_435 <= (fillup_transition == 1'b1) ? i_input_data[1035 % IN_WIDTH] : pong_storage_data_435 ^ i_input_data[1035 % IN_WIDTH];
                default: pong_storage_data_435 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_435;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_435 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_435;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_435 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_435;
            end
        end
    end
end

logic ping_storage_data_436;
logic pong_storage_data_436;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_436 <= 1'b0;
        pong_storage_data_436 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                205 / IN_WIDTH: ping_storage_data_436 <= (fillup_transition == 1'b1) ? i_input_data[205 % IN_WIDTH] : ping_storage_data_436 ^ i_input_data[205 % IN_WIDTH];
                640 / IN_WIDTH: ping_storage_data_436 <= (fillup_transition == 1'b1) ? i_input_data[640 % IN_WIDTH] : ping_storage_data_436 ^ i_input_data[640 % IN_WIDTH];
                875 / IN_WIDTH: ping_storage_data_436 <= (fillup_transition == 1'b1) ? i_input_data[875 % IN_WIDTH] : ping_storage_data_436 ^ i_input_data[875 % IN_WIDTH];
                1036 / IN_WIDTH: ping_storage_data_436 <= (fillup_transition == 1'b1) ? i_input_data[1036 % IN_WIDTH] : ping_storage_data_436 ^ i_input_data[1036 % IN_WIDTH];
                default: ping_storage_data_436 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_436;
                endcase
            end else begin
                case (input_count)
                205 / IN_WIDTH: pong_storage_data_436 <= (fillup_transition == 1'b1) ? i_input_data[205 % IN_WIDTH] : pong_storage_data_436 ^ i_input_data[205 % IN_WIDTH];
                640 / IN_WIDTH: pong_storage_data_436 <= (fillup_transition == 1'b1) ? i_input_data[640 % IN_WIDTH] : pong_storage_data_436 ^ i_input_data[640 % IN_WIDTH];
                875 / IN_WIDTH: pong_storage_data_436 <= (fillup_transition == 1'b1) ? i_input_data[875 % IN_WIDTH] : pong_storage_data_436 ^ i_input_data[875 % IN_WIDTH];
                1036 / IN_WIDTH: pong_storage_data_436 <= (fillup_transition == 1'b1) ? i_input_data[1036 % IN_WIDTH] : pong_storage_data_436 ^ i_input_data[1036 % IN_WIDTH];
                default: pong_storage_data_436 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_436;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_436 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_436;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_436 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_436;
            end
        end
    end
end

logic ping_storage_data_437;
logic pong_storage_data_437;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_437 <= 1'b0;
        pong_storage_data_437 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                206 / IN_WIDTH: ping_storage_data_437 <= (fillup_transition == 1'b1) ? i_input_data[206 % IN_WIDTH] : ping_storage_data_437 ^ i_input_data[206 % IN_WIDTH];
                641 / IN_WIDTH: ping_storage_data_437 <= (fillup_transition == 1'b1) ? i_input_data[641 % IN_WIDTH] : ping_storage_data_437 ^ i_input_data[641 % IN_WIDTH];
                876 / IN_WIDTH: ping_storage_data_437 <= (fillup_transition == 1'b1) ? i_input_data[876 % IN_WIDTH] : ping_storage_data_437 ^ i_input_data[876 % IN_WIDTH];
                1037 / IN_WIDTH: ping_storage_data_437 <= (fillup_transition == 1'b1) ? i_input_data[1037 % IN_WIDTH] : ping_storage_data_437 ^ i_input_data[1037 % IN_WIDTH];
                default: ping_storage_data_437 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_437;
                endcase
            end else begin
                case (input_count)
                206 / IN_WIDTH: pong_storage_data_437 <= (fillup_transition == 1'b1) ? i_input_data[206 % IN_WIDTH] : pong_storage_data_437 ^ i_input_data[206 % IN_WIDTH];
                641 / IN_WIDTH: pong_storage_data_437 <= (fillup_transition == 1'b1) ? i_input_data[641 % IN_WIDTH] : pong_storage_data_437 ^ i_input_data[641 % IN_WIDTH];
                876 / IN_WIDTH: pong_storage_data_437 <= (fillup_transition == 1'b1) ? i_input_data[876 % IN_WIDTH] : pong_storage_data_437 ^ i_input_data[876 % IN_WIDTH];
                1037 / IN_WIDTH: pong_storage_data_437 <= (fillup_transition == 1'b1) ? i_input_data[1037 % IN_WIDTH] : pong_storage_data_437 ^ i_input_data[1037 % IN_WIDTH];
                default: pong_storage_data_437 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_437;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_437 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_437;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_437 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_437;
            end
        end
    end
end

logic ping_storage_data_438;
logic pong_storage_data_438;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_438 <= 1'b0;
        pong_storage_data_438 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                207 / IN_WIDTH: ping_storage_data_438 <= (fillup_transition == 1'b1) ? i_input_data[207 % IN_WIDTH] : ping_storage_data_438 ^ i_input_data[207 % IN_WIDTH];
                642 / IN_WIDTH: ping_storage_data_438 <= (fillup_transition == 1'b1) ? i_input_data[642 % IN_WIDTH] : ping_storage_data_438 ^ i_input_data[642 % IN_WIDTH];
                877 / IN_WIDTH: ping_storage_data_438 <= (fillup_transition == 1'b1) ? i_input_data[877 % IN_WIDTH] : ping_storage_data_438 ^ i_input_data[877 % IN_WIDTH];
                1038 / IN_WIDTH: ping_storage_data_438 <= (fillup_transition == 1'b1) ? i_input_data[1038 % IN_WIDTH] : ping_storage_data_438 ^ i_input_data[1038 % IN_WIDTH];
                default: ping_storage_data_438 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_438;
                endcase
            end else begin
                case (input_count)
                207 / IN_WIDTH: pong_storage_data_438 <= (fillup_transition == 1'b1) ? i_input_data[207 % IN_WIDTH] : pong_storage_data_438 ^ i_input_data[207 % IN_WIDTH];
                642 / IN_WIDTH: pong_storage_data_438 <= (fillup_transition == 1'b1) ? i_input_data[642 % IN_WIDTH] : pong_storage_data_438 ^ i_input_data[642 % IN_WIDTH];
                877 / IN_WIDTH: pong_storage_data_438 <= (fillup_transition == 1'b1) ? i_input_data[877 % IN_WIDTH] : pong_storage_data_438 ^ i_input_data[877 % IN_WIDTH];
                1038 / IN_WIDTH: pong_storage_data_438 <= (fillup_transition == 1'b1) ? i_input_data[1038 % IN_WIDTH] : pong_storage_data_438 ^ i_input_data[1038 % IN_WIDTH];
                default: pong_storage_data_438 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_438;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_438 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_438;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_438 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_438;
            end
        end
    end
end

logic ping_storage_data_439;
logic pong_storage_data_439;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_439 <= 1'b0;
        pong_storage_data_439 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                208 / IN_WIDTH: ping_storage_data_439 <= (fillup_transition == 1'b1) ? i_input_data[208 % IN_WIDTH] : ping_storage_data_439 ^ i_input_data[208 % IN_WIDTH];
                643 / IN_WIDTH: ping_storage_data_439 <= (fillup_transition == 1'b1) ? i_input_data[643 % IN_WIDTH] : ping_storage_data_439 ^ i_input_data[643 % IN_WIDTH];
                878 / IN_WIDTH: ping_storage_data_439 <= (fillup_transition == 1'b1) ? i_input_data[878 % IN_WIDTH] : ping_storage_data_439 ^ i_input_data[878 % IN_WIDTH];
                1039 / IN_WIDTH: ping_storage_data_439 <= (fillup_transition == 1'b1) ? i_input_data[1039 % IN_WIDTH] : ping_storage_data_439 ^ i_input_data[1039 % IN_WIDTH];
                default: ping_storage_data_439 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_439;
                endcase
            end else begin
                case (input_count)
                208 / IN_WIDTH: pong_storage_data_439 <= (fillup_transition == 1'b1) ? i_input_data[208 % IN_WIDTH] : pong_storage_data_439 ^ i_input_data[208 % IN_WIDTH];
                643 / IN_WIDTH: pong_storage_data_439 <= (fillup_transition == 1'b1) ? i_input_data[643 % IN_WIDTH] : pong_storage_data_439 ^ i_input_data[643 % IN_WIDTH];
                878 / IN_WIDTH: pong_storage_data_439 <= (fillup_transition == 1'b1) ? i_input_data[878 % IN_WIDTH] : pong_storage_data_439 ^ i_input_data[878 % IN_WIDTH];
                1039 / IN_WIDTH: pong_storage_data_439 <= (fillup_transition == 1'b1) ? i_input_data[1039 % IN_WIDTH] : pong_storage_data_439 ^ i_input_data[1039 % IN_WIDTH];
                default: pong_storage_data_439 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_439;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_439 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_439;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_439 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_439;
            end
        end
    end
end

logic ping_storage_data_440;
logic pong_storage_data_440;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_440 <= 1'b0;
        pong_storage_data_440 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                209 / IN_WIDTH: ping_storage_data_440 <= (fillup_transition == 1'b1) ? i_input_data[209 % IN_WIDTH] : ping_storage_data_440 ^ i_input_data[209 % IN_WIDTH];
                644 / IN_WIDTH: ping_storage_data_440 <= (fillup_transition == 1'b1) ? i_input_data[644 % IN_WIDTH] : ping_storage_data_440 ^ i_input_data[644 % IN_WIDTH];
                879 / IN_WIDTH: ping_storage_data_440 <= (fillup_transition == 1'b1) ? i_input_data[879 % IN_WIDTH] : ping_storage_data_440 ^ i_input_data[879 % IN_WIDTH];
                1040 / IN_WIDTH: ping_storage_data_440 <= (fillup_transition == 1'b1) ? i_input_data[1040 % IN_WIDTH] : ping_storage_data_440 ^ i_input_data[1040 % IN_WIDTH];
                default: ping_storage_data_440 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_440;
                endcase
            end else begin
                case (input_count)
                209 / IN_WIDTH: pong_storage_data_440 <= (fillup_transition == 1'b1) ? i_input_data[209 % IN_WIDTH] : pong_storage_data_440 ^ i_input_data[209 % IN_WIDTH];
                644 / IN_WIDTH: pong_storage_data_440 <= (fillup_transition == 1'b1) ? i_input_data[644 % IN_WIDTH] : pong_storage_data_440 ^ i_input_data[644 % IN_WIDTH];
                879 / IN_WIDTH: pong_storage_data_440 <= (fillup_transition == 1'b1) ? i_input_data[879 % IN_WIDTH] : pong_storage_data_440 ^ i_input_data[879 % IN_WIDTH];
                1040 / IN_WIDTH: pong_storage_data_440 <= (fillup_transition == 1'b1) ? i_input_data[1040 % IN_WIDTH] : pong_storage_data_440 ^ i_input_data[1040 % IN_WIDTH];
                default: pong_storage_data_440 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_440;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_440 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_440;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_440 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_440;
            end
        end
    end
end

logic ping_storage_data_441;
logic pong_storage_data_441;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_441 <= 1'b0;
        pong_storage_data_441 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                210 / IN_WIDTH: ping_storage_data_441 <= (fillup_transition == 1'b1) ? i_input_data[210 % IN_WIDTH] : ping_storage_data_441 ^ i_input_data[210 % IN_WIDTH];
                645 / IN_WIDTH: ping_storage_data_441 <= (fillup_transition == 1'b1) ? i_input_data[645 % IN_WIDTH] : ping_storage_data_441 ^ i_input_data[645 % IN_WIDTH];
                880 / IN_WIDTH: ping_storage_data_441 <= (fillup_transition == 1'b1) ? i_input_data[880 % IN_WIDTH] : ping_storage_data_441 ^ i_input_data[880 % IN_WIDTH];
                1041 / IN_WIDTH: ping_storage_data_441 <= (fillup_transition == 1'b1) ? i_input_data[1041 % IN_WIDTH] : ping_storage_data_441 ^ i_input_data[1041 % IN_WIDTH];
                default: ping_storage_data_441 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_441;
                endcase
            end else begin
                case (input_count)
                210 / IN_WIDTH: pong_storage_data_441 <= (fillup_transition == 1'b1) ? i_input_data[210 % IN_WIDTH] : pong_storage_data_441 ^ i_input_data[210 % IN_WIDTH];
                645 / IN_WIDTH: pong_storage_data_441 <= (fillup_transition == 1'b1) ? i_input_data[645 % IN_WIDTH] : pong_storage_data_441 ^ i_input_data[645 % IN_WIDTH];
                880 / IN_WIDTH: pong_storage_data_441 <= (fillup_transition == 1'b1) ? i_input_data[880 % IN_WIDTH] : pong_storage_data_441 ^ i_input_data[880 % IN_WIDTH];
                1041 / IN_WIDTH: pong_storage_data_441 <= (fillup_transition == 1'b1) ? i_input_data[1041 % IN_WIDTH] : pong_storage_data_441 ^ i_input_data[1041 % IN_WIDTH];
                default: pong_storage_data_441 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_441;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_441 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_441;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_441 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_441;
            end
        end
    end
end

logic ping_storage_data_442;
logic pong_storage_data_442;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_442 <= 1'b0;
        pong_storage_data_442 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                211 / IN_WIDTH: ping_storage_data_442 <= (fillup_transition == 1'b1) ? i_input_data[211 % IN_WIDTH] : ping_storage_data_442 ^ i_input_data[211 % IN_WIDTH];
                646 / IN_WIDTH: ping_storage_data_442 <= (fillup_transition == 1'b1) ? i_input_data[646 % IN_WIDTH] : ping_storage_data_442 ^ i_input_data[646 % IN_WIDTH];
                881 / IN_WIDTH: ping_storage_data_442 <= (fillup_transition == 1'b1) ? i_input_data[881 % IN_WIDTH] : ping_storage_data_442 ^ i_input_data[881 % IN_WIDTH];
                1042 / IN_WIDTH: ping_storage_data_442 <= (fillup_transition == 1'b1) ? i_input_data[1042 % IN_WIDTH] : ping_storage_data_442 ^ i_input_data[1042 % IN_WIDTH];
                default: ping_storage_data_442 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_442;
                endcase
            end else begin
                case (input_count)
                211 / IN_WIDTH: pong_storage_data_442 <= (fillup_transition == 1'b1) ? i_input_data[211 % IN_WIDTH] : pong_storage_data_442 ^ i_input_data[211 % IN_WIDTH];
                646 / IN_WIDTH: pong_storage_data_442 <= (fillup_transition == 1'b1) ? i_input_data[646 % IN_WIDTH] : pong_storage_data_442 ^ i_input_data[646 % IN_WIDTH];
                881 / IN_WIDTH: pong_storage_data_442 <= (fillup_transition == 1'b1) ? i_input_data[881 % IN_WIDTH] : pong_storage_data_442 ^ i_input_data[881 % IN_WIDTH];
                1042 / IN_WIDTH: pong_storage_data_442 <= (fillup_transition == 1'b1) ? i_input_data[1042 % IN_WIDTH] : pong_storage_data_442 ^ i_input_data[1042 % IN_WIDTH];
                default: pong_storage_data_442 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_442;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_442 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_442;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_442 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_442;
            end
        end
    end
end

logic ping_storage_data_443;
logic pong_storage_data_443;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_443 <= 1'b0;
        pong_storage_data_443 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                212 / IN_WIDTH: ping_storage_data_443 <= (fillup_transition == 1'b1) ? i_input_data[212 % IN_WIDTH] : ping_storage_data_443 ^ i_input_data[212 % IN_WIDTH];
                647 / IN_WIDTH: ping_storage_data_443 <= (fillup_transition == 1'b1) ? i_input_data[647 % IN_WIDTH] : ping_storage_data_443 ^ i_input_data[647 % IN_WIDTH];
                882 / IN_WIDTH: ping_storage_data_443 <= (fillup_transition == 1'b1) ? i_input_data[882 % IN_WIDTH] : ping_storage_data_443 ^ i_input_data[882 % IN_WIDTH];
                1043 / IN_WIDTH: ping_storage_data_443 <= (fillup_transition == 1'b1) ? i_input_data[1043 % IN_WIDTH] : ping_storage_data_443 ^ i_input_data[1043 % IN_WIDTH];
                default: ping_storage_data_443 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_443;
                endcase
            end else begin
                case (input_count)
                212 / IN_WIDTH: pong_storage_data_443 <= (fillup_transition == 1'b1) ? i_input_data[212 % IN_WIDTH] : pong_storage_data_443 ^ i_input_data[212 % IN_WIDTH];
                647 / IN_WIDTH: pong_storage_data_443 <= (fillup_transition == 1'b1) ? i_input_data[647 % IN_WIDTH] : pong_storage_data_443 ^ i_input_data[647 % IN_WIDTH];
                882 / IN_WIDTH: pong_storage_data_443 <= (fillup_transition == 1'b1) ? i_input_data[882 % IN_WIDTH] : pong_storage_data_443 ^ i_input_data[882 % IN_WIDTH];
                1043 / IN_WIDTH: pong_storage_data_443 <= (fillup_transition == 1'b1) ? i_input_data[1043 % IN_WIDTH] : pong_storage_data_443 ^ i_input_data[1043 % IN_WIDTH];
                default: pong_storage_data_443 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_443;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_443 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_443;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_443 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_443;
            end
        end
    end
end

logic ping_storage_data_444;
logic pong_storage_data_444;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_444 <= 1'b0;
        pong_storage_data_444 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                213 / IN_WIDTH: ping_storage_data_444 <= (fillup_transition == 1'b1) ? i_input_data[213 % IN_WIDTH] : ping_storage_data_444 ^ i_input_data[213 % IN_WIDTH];
                648 / IN_WIDTH: ping_storage_data_444 <= (fillup_transition == 1'b1) ? i_input_data[648 % IN_WIDTH] : ping_storage_data_444 ^ i_input_data[648 % IN_WIDTH];
                883 / IN_WIDTH: ping_storage_data_444 <= (fillup_transition == 1'b1) ? i_input_data[883 % IN_WIDTH] : ping_storage_data_444 ^ i_input_data[883 % IN_WIDTH];
                1044 / IN_WIDTH: ping_storage_data_444 <= (fillup_transition == 1'b1) ? i_input_data[1044 % IN_WIDTH] : ping_storage_data_444 ^ i_input_data[1044 % IN_WIDTH];
                default: ping_storage_data_444 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_444;
                endcase
            end else begin
                case (input_count)
                213 / IN_WIDTH: pong_storage_data_444 <= (fillup_transition == 1'b1) ? i_input_data[213 % IN_WIDTH] : pong_storage_data_444 ^ i_input_data[213 % IN_WIDTH];
                648 / IN_WIDTH: pong_storage_data_444 <= (fillup_transition == 1'b1) ? i_input_data[648 % IN_WIDTH] : pong_storage_data_444 ^ i_input_data[648 % IN_WIDTH];
                883 / IN_WIDTH: pong_storage_data_444 <= (fillup_transition == 1'b1) ? i_input_data[883 % IN_WIDTH] : pong_storage_data_444 ^ i_input_data[883 % IN_WIDTH];
                1044 / IN_WIDTH: pong_storage_data_444 <= (fillup_transition == 1'b1) ? i_input_data[1044 % IN_WIDTH] : pong_storage_data_444 ^ i_input_data[1044 % IN_WIDTH];
                default: pong_storage_data_444 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_444;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_444 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_444;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_444 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_444;
            end
        end
    end
end

logic ping_storage_data_445;
logic pong_storage_data_445;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_445 <= 1'b0;
        pong_storage_data_445 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                214 / IN_WIDTH: ping_storage_data_445 <= (fillup_transition == 1'b1) ? i_input_data[214 % IN_WIDTH] : ping_storage_data_445 ^ i_input_data[214 % IN_WIDTH];
                649 / IN_WIDTH: ping_storage_data_445 <= (fillup_transition == 1'b1) ? i_input_data[649 % IN_WIDTH] : ping_storage_data_445 ^ i_input_data[649 % IN_WIDTH];
                884 / IN_WIDTH: ping_storage_data_445 <= (fillup_transition == 1'b1) ? i_input_data[884 % IN_WIDTH] : ping_storage_data_445 ^ i_input_data[884 % IN_WIDTH];
                1045 / IN_WIDTH: ping_storage_data_445 <= (fillup_transition == 1'b1) ? i_input_data[1045 % IN_WIDTH] : ping_storage_data_445 ^ i_input_data[1045 % IN_WIDTH];
                default: ping_storage_data_445 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_445;
                endcase
            end else begin
                case (input_count)
                214 / IN_WIDTH: pong_storage_data_445 <= (fillup_transition == 1'b1) ? i_input_data[214 % IN_WIDTH] : pong_storage_data_445 ^ i_input_data[214 % IN_WIDTH];
                649 / IN_WIDTH: pong_storage_data_445 <= (fillup_transition == 1'b1) ? i_input_data[649 % IN_WIDTH] : pong_storage_data_445 ^ i_input_data[649 % IN_WIDTH];
                884 / IN_WIDTH: pong_storage_data_445 <= (fillup_transition == 1'b1) ? i_input_data[884 % IN_WIDTH] : pong_storage_data_445 ^ i_input_data[884 % IN_WIDTH];
                1045 / IN_WIDTH: pong_storage_data_445 <= (fillup_transition == 1'b1) ? i_input_data[1045 % IN_WIDTH] : pong_storage_data_445 ^ i_input_data[1045 % IN_WIDTH];
                default: pong_storage_data_445 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_445;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_445 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_445;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_445 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_445;
            end
        end
    end
end

logic ping_storage_data_446;
logic pong_storage_data_446;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_446 <= 1'b0;
        pong_storage_data_446 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                215 / IN_WIDTH: ping_storage_data_446 <= (fillup_transition == 1'b1) ? i_input_data[215 % IN_WIDTH] : ping_storage_data_446 ^ i_input_data[215 % IN_WIDTH];
                650 / IN_WIDTH: ping_storage_data_446 <= (fillup_transition == 1'b1) ? i_input_data[650 % IN_WIDTH] : ping_storage_data_446 ^ i_input_data[650 % IN_WIDTH];
                885 / IN_WIDTH: ping_storage_data_446 <= (fillup_transition == 1'b1) ? i_input_data[885 % IN_WIDTH] : ping_storage_data_446 ^ i_input_data[885 % IN_WIDTH];
                1046 / IN_WIDTH: ping_storage_data_446 <= (fillup_transition == 1'b1) ? i_input_data[1046 % IN_WIDTH] : ping_storage_data_446 ^ i_input_data[1046 % IN_WIDTH];
                default: ping_storage_data_446 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_446;
                endcase
            end else begin
                case (input_count)
                215 / IN_WIDTH: pong_storage_data_446 <= (fillup_transition == 1'b1) ? i_input_data[215 % IN_WIDTH] : pong_storage_data_446 ^ i_input_data[215 % IN_WIDTH];
                650 / IN_WIDTH: pong_storage_data_446 <= (fillup_transition == 1'b1) ? i_input_data[650 % IN_WIDTH] : pong_storage_data_446 ^ i_input_data[650 % IN_WIDTH];
                885 / IN_WIDTH: pong_storage_data_446 <= (fillup_transition == 1'b1) ? i_input_data[885 % IN_WIDTH] : pong_storage_data_446 ^ i_input_data[885 % IN_WIDTH];
                1046 / IN_WIDTH: pong_storage_data_446 <= (fillup_transition == 1'b1) ? i_input_data[1046 % IN_WIDTH] : pong_storage_data_446 ^ i_input_data[1046 % IN_WIDTH];
                default: pong_storage_data_446 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_446;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_446 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_446;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_446 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_446;
            end
        end
    end
end

logic ping_storage_data_447;
logic pong_storage_data_447;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_447 <= 1'b0;
        pong_storage_data_447 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                216 / IN_WIDTH: ping_storage_data_447 <= (fillup_transition == 1'b1) ? i_input_data[216 % IN_WIDTH] : ping_storage_data_447 ^ i_input_data[216 % IN_WIDTH];
                651 / IN_WIDTH: ping_storage_data_447 <= (fillup_transition == 1'b1) ? i_input_data[651 % IN_WIDTH] : ping_storage_data_447 ^ i_input_data[651 % IN_WIDTH];
                886 / IN_WIDTH: ping_storage_data_447 <= (fillup_transition == 1'b1) ? i_input_data[886 % IN_WIDTH] : ping_storage_data_447 ^ i_input_data[886 % IN_WIDTH];
                1047 / IN_WIDTH: ping_storage_data_447 <= (fillup_transition == 1'b1) ? i_input_data[1047 % IN_WIDTH] : ping_storage_data_447 ^ i_input_data[1047 % IN_WIDTH];
                default: ping_storage_data_447 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_447;
                endcase
            end else begin
                case (input_count)
                216 / IN_WIDTH: pong_storage_data_447 <= (fillup_transition == 1'b1) ? i_input_data[216 % IN_WIDTH] : pong_storage_data_447 ^ i_input_data[216 % IN_WIDTH];
                651 / IN_WIDTH: pong_storage_data_447 <= (fillup_transition == 1'b1) ? i_input_data[651 % IN_WIDTH] : pong_storage_data_447 ^ i_input_data[651 % IN_WIDTH];
                886 / IN_WIDTH: pong_storage_data_447 <= (fillup_transition == 1'b1) ? i_input_data[886 % IN_WIDTH] : pong_storage_data_447 ^ i_input_data[886 % IN_WIDTH];
                1047 / IN_WIDTH: pong_storage_data_447 <= (fillup_transition == 1'b1) ? i_input_data[1047 % IN_WIDTH] : pong_storage_data_447 ^ i_input_data[1047 % IN_WIDTH];
                default: pong_storage_data_447 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_447;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_447 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_447;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_447 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_447;
            end
        end
    end
end

logic ping_storage_data_448;
logic pong_storage_data_448;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_448 <= 1'b0;
        pong_storage_data_448 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                217 / IN_WIDTH: ping_storage_data_448 <= (fillup_transition == 1'b1) ? i_input_data[217 % IN_WIDTH] : ping_storage_data_448 ^ i_input_data[217 % IN_WIDTH];
                652 / IN_WIDTH: ping_storage_data_448 <= (fillup_transition == 1'b1) ? i_input_data[652 % IN_WIDTH] : ping_storage_data_448 ^ i_input_data[652 % IN_WIDTH];
                887 / IN_WIDTH: ping_storage_data_448 <= (fillup_transition == 1'b1) ? i_input_data[887 % IN_WIDTH] : ping_storage_data_448 ^ i_input_data[887 % IN_WIDTH];
                1048 / IN_WIDTH: ping_storage_data_448 <= (fillup_transition == 1'b1) ? i_input_data[1048 % IN_WIDTH] : ping_storage_data_448 ^ i_input_data[1048 % IN_WIDTH];
                default: ping_storage_data_448 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_448;
                endcase
            end else begin
                case (input_count)
                217 / IN_WIDTH: pong_storage_data_448 <= (fillup_transition == 1'b1) ? i_input_data[217 % IN_WIDTH] : pong_storage_data_448 ^ i_input_data[217 % IN_WIDTH];
                652 / IN_WIDTH: pong_storage_data_448 <= (fillup_transition == 1'b1) ? i_input_data[652 % IN_WIDTH] : pong_storage_data_448 ^ i_input_data[652 % IN_WIDTH];
                887 / IN_WIDTH: pong_storage_data_448 <= (fillup_transition == 1'b1) ? i_input_data[887 % IN_WIDTH] : pong_storage_data_448 ^ i_input_data[887 % IN_WIDTH];
                1048 / IN_WIDTH: pong_storage_data_448 <= (fillup_transition == 1'b1) ? i_input_data[1048 % IN_WIDTH] : pong_storage_data_448 ^ i_input_data[1048 % IN_WIDTH];
                default: pong_storage_data_448 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_448;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_448 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_448;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_448 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_448;
            end
        end
    end
end

logic ping_storage_data_449;
logic pong_storage_data_449;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_449 <= 1'b0;
        pong_storage_data_449 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                218 / IN_WIDTH: ping_storage_data_449 <= (fillup_transition == 1'b1) ? i_input_data[218 % IN_WIDTH] : ping_storage_data_449 ^ i_input_data[218 % IN_WIDTH];
                653 / IN_WIDTH: ping_storage_data_449 <= (fillup_transition == 1'b1) ? i_input_data[653 % IN_WIDTH] : ping_storage_data_449 ^ i_input_data[653 % IN_WIDTH];
                888 / IN_WIDTH: ping_storage_data_449 <= (fillup_transition == 1'b1) ? i_input_data[888 % IN_WIDTH] : ping_storage_data_449 ^ i_input_data[888 % IN_WIDTH];
                1049 / IN_WIDTH: ping_storage_data_449 <= (fillup_transition == 1'b1) ? i_input_data[1049 % IN_WIDTH] : ping_storage_data_449 ^ i_input_data[1049 % IN_WIDTH];
                default: ping_storage_data_449 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_449;
                endcase
            end else begin
                case (input_count)
                218 / IN_WIDTH: pong_storage_data_449 <= (fillup_transition == 1'b1) ? i_input_data[218 % IN_WIDTH] : pong_storage_data_449 ^ i_input_data[218 % IN_WIDTH];
                653 / IN_WIDTH: pong_storage_data_449 <= (fillup_transition == 1'b1) ? i_input_data[653 % IN_WIDTH] : pong_storage_data_449 ^ i_input_data[653 % IN_WIDTH];
                888 / IN_WIDTH: pong_storage_data_449 <= (fillup_transition == 1'b1) ? i_input_data[888 % IN_WIDTH] : pong_storage_data_449 ^ i_input_data[888 % IN_WIDTH];
                1049 / IN_WIDTH: pong_storage_data_449 <= (fillup_transition == 1'b1) ? i_input_data[1049 % IN_WIDTH] : pong_storage_data_449 ^ i_input_data[1049 % IN_WIDTH];
                default: pong_storage_data_449 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_449;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_449 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_449;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_449 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_449;
            end
        end
    end
end

logic ping_storage_data_450;
logic pong_storage_data_450;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_450 <= 1'b0;
        pong_storage_data_450 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                219 / IN_WIDTH: ping_storage_data_450 <= (fillup_transition == 1'b1) ? i_input_data[219 % IN_WIDTH] : ping_storage_data_450 ^ i_input_data[219 % IN_WIDTH];
                654 / IN_WIDTH: ping_storage_data_450 <= (fillup_transition == 1'b1) ? i_input_data[654 % IN_WIDTH] : ping_storage_data_450 ^ i_input_data[654 % IN_WIDTH];
                889 / IN_WIDTH: ping_storage_data_450 <= (fillup_transition == 1'b1) ? i_input_data[889 % IN_WIDTH] : ping_storage_data_450 ^ i_input_data[889 % IN_WIDTH];
                1050 / IN_WIDTH: ping_storage_data_450 <= (fillup_transition == 1'b1) ? i_input_data[1050 % IN_WIDTH] : ping_storage_data_450 ^ i_input_data[1050 % IN_WIDTH];
                default: ping_storage_data_450 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_450;
                endcase
            end else begin
                case (input_count)
                219 / IN_WIDTH: pong_storage_data_450 <= (fillup_transition == 1'b1) ? i_input_data[219 % IN_WIDTH] : pong_storage_data_450 ^ i_input_data[219 % IN_WIDTH];
                654 / IN_WIDTH: pong_storage_data_450 <= (fillup_transition == 1'b1) ? i_input_data[654 % IN_WIDTH] : pong_storage_data_450 ^ i_input_data[654 % IN_WIDTH];
                889 / IN_WIDTH: pong_storage_data_450 <= (fillup_transition == 1'b1) ? i_input_data[889 % IN_WIDTH] : pong_storage_data_450 ^ i_input_data[889 % IN_WIDTH];
                1050 / IN_WIDTH: pong_storage_data_450 <= (fillup_transition == 1'b1) ? i_input_data[1050 % IN_WIDTH] : pong_storage_data_450 ^ i_input_data[1050 % IN_WIDTH];
                default: pong_storage_data_450 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_450;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_450 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_450;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_450 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_450;
            end
        end
    end
end

logic ping_storage_data_451;
logic pong_storage_data_451;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_451 <= 1'b0;
        pong_storage_data_451 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                220 / IN_WIDTH: ping_storage_data_451 <= (fillup_transition == 1'b1) ? i_input_data[220 % IN_WIDTH] : ping_storage_data_451 ^ i_input_data[220 % IN_WIDTH];
                655 / IN_WIDTH: ping_storage_data_451 <= (fillup_transition == 1'b1) ? i_input_data[655 % IN_WIDTH] : ping_storage_data_451 ^ i_input_data[655 % IN_WIDTH];
                890 / IN_WIDTH: ping_storage_data_451 <= (fillup_transition == 1'b1) ? i_input_data[890 % IN_WIDTH] : ping_storage_data_451 ^ i_input_data[890 % IN_WIDTH];
                1051 / IN_WIDTH: ping_storage_data_451 <= (fillup_transition == 1'b1) ? i_input_data[1051 % IN_WIDTH] : ping_storage_data_451 ^ i_input_data[1051 % IN_WIDTH];
                default: ping_storage_data_451 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_451;
                endcase
            end else begin
                case (input_count)
                220 / IN_WIDTH: pong_storage_data_451 <= (fillup_transition == 1'b1) ? i_input_data[220 % IN_WIDTH] : pong_storage_data_451 ^ i_input_data[220 % IN_WIDTH];
                655 / IN_WIDTH: pong_storage_data_451 <= (fillup_transition == 1'b1) ? i_input_data[655 % IN_WIDTH] : pong_storage_data_451 ^ i_input_data[655 % IN_WIDTH];
                890 / IN_WIDTH: pong_storage_data_451 <= (fillup_transition == 1'b1) ? i_input_data[890 % IN_WIDTH] : pong_storage_data_451 ^ i_input_data[890 % IN_WIDTH];
                1051 / IN_WIDTH: pong_storage_data_451 <= (fillup_transition == 1'b1) ? i_input_data[1051 % IN_WIDTH] : pong_storage_data_451 ^ i_input_data[1051 % IN_WIDTH];
                default: pong_storage_data_451 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_451;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_451 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_451;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_451 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_451;
            end
        end
    end
end

logic ping_storage_data_452;
logic pong_storage_data_452;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_452 <= 1'b0;
        pong_storage_data_452 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                221 / IN_WIDTH: ping_storage_data_452 <= (fillup_transition == 1'b1) ? i_input_data[221 % IN_WIDTH] : ping_storage_data_452 ^ i_input_data[221 % IN_WIDTH];
                656 / IN_WIDTH: ping_storage_data_452 <= (fillup_transition == 1'b1) ? i_input_data[656 % IN_WIDTH] : ping_storage_data_452 ^ i_input_data[656 % IN_WIDTH];
                891 / IN_WIDTH: ping_storage_data_452 <= (fillup_transition == 1'b1) ? i_input_data[891 % IN_WIDTH] : ping_storage_data_452 ^ i_input_data[891 % IN_WIDTH];
                1052 / IN_WIDTH: ping_storage_data_452 <= (fillup_transition == 1'b1) ? i_input_data[1052 % IN_WIDTH] : ping_storage_data_452 ^ i_input_data[1052 % IN_WIDTH];
                default: ping_storage_data_452 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_452;
                endcase
            end else begin
                case (input_count)
                221 / IN_WIDTH: pong_storage_data_452 <= (fillup_transition == 1'b1) ? i_input_data[221 % IN_WIDTH] : pong_storage_data_452 ^ i_input_data[221 % IN_WIDTH];
                656 / IN_WIDTH: pong_storage_data_452 <= (fillup_transition == 1'b1) ? i_input_data[656 % IN_WIDTH] : pong_storage_data_452 ^ i_input_data[656 % IN_WIDTH];
                891 / IN_WIDTH: pong_storage_data_452 <= (fillup_transition == 1'b1) ? i_input_data[891 % IN_WIDTH] : pong_storage_data_452 ^ i_input_data[891 % IN_WIDTH];
                1052 / IN_WIDTH: pong_storage_data_452 <= (fillup_transition == 1'b1) ? i_input_data[1052 % IN_WIDTH] : pong_storage_data_452 ^ i_input_data[1052 % IN_WIDTH];
                default: pong_storage_data_452 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_452;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_452 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_452;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_452 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_452;
            end
        end
    end
end

logic ping_storage_data_453;
logic pong_storage_data_453;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_453 <= 1'b0;
        pong_storage_data_453 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                222 / IN_WIDTH: ping_storage_data_453 <= (fillup_transition == 1'b1) ? i_input_data[222 % IN_WIDTH] : ping_storage_data_453 ^ i_input_data[222 % IN_WIDTH];
                657 / IN_WIDTH: ping_storage_data_453 <= (fillup_transition == 1'b1) ? i_input_data[657 % IN_WIDTH] : ping_storage_data_453 ^ i_input_data[657 % IN_WIDTH];
                892 / IN_WIDTH: ping_storage_data_453 <= (fillup_transition == 1'b1) ? i_input_data[892 % IN_WIDTH] : ping_storage_data_453 ^ i_input_data[892 % IN_WIDTH];
                1053 / IN_WIDTH: ping_storage_data_453 <= (fillup_transition == 1'b1) ? i_input_data[1053 % IN_WIDTH] : ping_storage_data_453 ^ i_input_data[1053 % IN_WIDTH];
                default: ping_storage_data_453 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_453;
                endcase
            end else begin
                case (input_count)
                222 / IN_WIDTH: pong_storage_data_453 <= (fillup_transition == 1'b1) ? i_input_data[222 % IN_WIDTH] : pong_storage_data_453 ^ i_input_data[222 % IN_WIDTH];
                657 / IN_WIDTH: pong_storage_data_453 <= (fillup_transition == 1'b1) ? i_input_data[657 % IN_WIDTH] : pong_storage_data_453 ^ i_input_data[657 % IN_WIDTH];
                892 / IN_WIDTH: pong_storage_data_453 <= (fillup_transition == 1'b1) ? i_input_data[892 % IN_WIDTH] : pong_storage_data_453 ^ i_input_data[892 % IN_WIDTH];
                1053 / IN_WIDTH: pong_storage_data_453 <= (fillup_transition == 1'b1) ? i_input_data[1053 % IN_WIDTH] : pong_storage_data_453 ^ i_input_data[1053 % IN_WIDTH];
                default: pong_storage_data_453 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_453;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_453 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_453;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_453 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_453;
            end
        end
    end
end

logic ping_storage_data_454;
logic pong_storage_data_454;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_454 <= 1'b0;
        pong_storage_data_454 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                223 / IN_WIDTH: ping_storage_data_454 <= (fillup_transition == 1'b1) ? i_input_data[223 % IN_WIDTH] : ping_storage_data_454 ^ i_input_data[223 % IN_WIDTH];
                658 / IN_WIDTH: ping_storage_data_454 <= (fillup_transition == 1'b1) ? i_input_data[658 % IN_WIDTH] : ping_storage_data_454 ^ i_input_data[658 % IN_WIDTH];
                893 / IN_WIDTH: ping_storage_data_454 <= (fillup_transition == 1'b1) ? i_input_data[893 % IN_WIDTH] : ping_storage_data_454 ^ i_input_data[893 % IN_WIDTH];
                1054 / IN_WIDTH: ping_storage_data_454 <= (fillup_transition == 1'b1) ? i_input_data[1054 % IN_WIDTH] : ping_storage_data_454 ^ i_input_data[1054 % IN_WIDTH];
                default: ping_storage_data_454 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_454;
                endcase
            end else begin
                case (input_count)
                223 / IN_WIDTH: pong_storage_data_454 <= (fillup_transition == 1'b1) ? i_input_data[223 % IN_WIDTH] : pong_storage_data_454 ^ i_input_data[223 % IN_WIDTH];
                658 / IN_WIDTH: pong_storage_data_454 <= (fillup_transition == 1'b1) ? i_input_data[658 % IN_WIDTH] : pong_storage_data_454 ^ i_input_data[658 % IN_WIDTH];
                893 / IN_WIDTH: pong_storage_data_454 <= (fillup_transition == 1'b1) ? i_input_data[893 % IN_WIDTH] : pong_storage_data_454 ^ i_input_data[893 % IN_WIDTH];
                1054 / IN_WIDTH: pong_storage_data_454 <= (fillup_transition == 1'b1) ? i_input_data[1054 % IN_WIDTH] : pong_storage_data_454 ^ i_input_data[1054 % IN_WIDTH];
                default: pong_storage_data_454 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_454;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_454 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_454;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_454 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_454;
            end
        end
    end
end

logic ping_storage_data_455;
logic pong_storage_data_455;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_455 <= 1'b0;
        pong_storage_data_455 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                224 / IN_WIDTH: ping_storage_data_455 <= (fillup_transition == 1'b1) ? i_input_data[224 % IN_WIDTH] : ping_storage_data_455 ^ i_input_data[224 % IN_WIDTH];
                659 / IN_WIDTH: ping_storage_data_455 <= (fillup_transition == 1'b1) ? i_input_data[659 % IN_WIDTH] : ping_storage_data_455 ^ i_input_data[659 % IN_WIDTH];
                894 / IN_WIDTH: ping_storage_data_455 <= (fillup_transition == 1'b1) ? i_input_data[894 % IN_WIDTH] : ping_storage_data_455 ^ i_input_data[894 % IN_WIDTH];
                1055 / IN_WIDTH: ping_storage_data_455 <= (fillup_transition == 1'b1) ? i_input_data[1055 % IN_WIDTH] : ping_storage_data_455 ^ i_input_data[1055 % IN_WIDTH];
                default: ping_storage_data_455 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_455;
                endcase
            end else begin
                case (input_count)
                224 / IN_WIDTH: pong_storage_data_455 <= (fillup_transition == 1'b1) ? i_input_data[224 % IN_WIDTH] : pong_storage_data_455 ^ i_input_data[224 % IN_WIDTH];
                659 / IN_WIDTH: pong_storage_data_455 <= (fillup_transition == 1'b1) ? i_input_data[659 % IN_WIDTH] : pong_storage_data_455 ^ i_input_data[659 % IN_WIDTH];
                894 / IN_WIDTH: pong_storage_data_455 <= (fillup_transition == 1'b1) ? i_input_data[894 % IN_WIDTH] : pong_storage_data_455 ^ i_input_data[894 % IN_WIDTH];
                1055 / IN_WIDTH: pong_storage_data_455 <= (fillup_transition == 1'b1) ? i_input_data[1055 % IN_WIDTH] : pong_storage_data_455 ^ i_input_data[1055 % IN_WIDTH];
                default: pong_storage_data_455 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_455;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_455 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_455;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_455 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_455;
            end
        end
    end
end

logic ping_storage_data_456;
logic pong_storage_data_456;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_456 <= 1'b0;
        pong_storage_data_456 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                225 / IN_WIDTH: ping_storage_data_456 <= (fillup_transition == 1'b1) ? i_input_data[225 % IN_WIDTH] : ping_storage_data_456 ^ i_input_data[225 % IN_WIDTH];
                660 / IN_WIDTH: ping_storage_data_456 <= (fillup_transition == 1'b1) ? i_input_data[660 % IN_WIDTH] : ping_storage_data_456 ^ i_input_data[660 % IN_WIDTH];
                895 / IN_WIDTH: ping_storage_data_456 <= (fillup_transition == 1'b1) ? i_input_data[895 % IN_WIDTH] : ping_storage_data_456 ^ i_input_data[895 % IN_WIDTH];
                960 / IN_WIDTH: ping_storage_data_456 <= (fillup_transition == 1'b1) ? i_input_data[960 % IN_WIDTH] : ping_storage_data_456 ^ i_input_data[960 % IN_WIDTH];
                default: ping_storage_data_456 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_456;
                endcase
            end else begin
                case (input_count)
                225 / IN_WIDTH: pong_storage_data_456 <= (fillup_transition == 1'b1) ? i_input_data[225 % IN_WIDTH] : pong_storage_data_456 ^ i_input_data[225 % IN_WIDTH];
                660 / IN_WIDTH: pong_storage_data_456 <= (fillup_transition == 1'b1) ? i_input_data[660 % IN_WIDTH] : pong_storage_data_456 ^ i_input_data[660 % IN_WIDTH];
                895 / IN_WIDTH: pong_storage_data_456 <= (fillup_transition == 1'b1) ? i_input_data[895 % IN_WIDTH] : pong_storage_data_456 ^ i_input_data[895 % IN_WIDTH];
                960 / IN_WIDTH: pong_storage_data_456 <= (fillup_transition == 1'b1) ? i_input_data[960 % IN_WIDTH] : pong_storage_data_456 ^ i_input_data[960 % IN_WIDTH];
                default: pong_storage_data_456 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_456;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_456 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_456;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_456 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_456;
            end
        end
    end
end

logic ping_storage_data_457;
logic pong_storage_data_457;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_457 <= 1'b0;
        pong_storage_data_457 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                226 / IN_WIDTH: ping_storage_data_457 <= (fillup_transition == 1'b1) ? i_input_data[226 % IN_WIDTH] : ping_storage_data_457 ^ i_input_data[226 % IN_WIDTH];
                661 / IN_WIDTH: ping_storage_data_457 <= (fillup_transition == 1'b1) ? i_input_data[661 % IN_WIDTH] : ping_storage_data_457 ^ i_input_data[661 % IN_WIDTH];
                896 / IN_WIDTH: ping_storage_data_457 <= (fillup_transition == 1'b1) ? i_input_data[896 % IN_WIDTH] : ping_storage_data_457 ^ i_input_data[896 % IN_WIDTH];
                961 / IN_WIDTH: ping_storage_data_457 <= (fillup_transition == 1'b1) ? i_input_data[961 % IN_WIDTH] : ping_storage_data_457 ^ i_input_data[961 % IN_WIDTH];
                default: ping_storage_data_457 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_457;
                endcase
            end else begin
                case (input_count)
                226 / IN_WIDTH: pong_storage_data_457 <= (fillup_transition == 1'b1) ? i_input_data[226 % IN_WIDTH] : pong_storage_data_457 ^ i_input_data[226 % IN_WIDTH];
                661 / IN_WIDTH: pong_storage_data_457 <= (fillup_transition == 1'b1) ? i_input_data[661 % IN_WIDTH] : pong_storage_data_457 ^ i_input_data[661 % IN_WIDTH];
                896 / IN_WIDTH: pong_storage_data_457 <= (fillup_transition == 1'b1) ? i_input_data[896 % IN_WIDTH] : pong_storage_data_457 ^ i_input_data[896 % IN_WIDTH];
                961 / IN_WIDTH: pong_storage_data_457 <= (fillup_transition == 1'b1) ? i_input_data[961 % IN_WIDTH] : pong_storage_data_457 ^ i_input_data[961 % IN_WIDTH];
                default: pong_storage_data_457 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_457;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_457 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_457;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_457 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_457;
            end
        end
    end
end

logic ping_storage_data_458;
logic pong_storage_data_458;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_458 <= 1'b0;
        pong_storage_data_458 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                227 / IN_WIDTH: ping_storage_data_458 <= (fillup_transition == 1'b1) ? i_input_data[227 % IN_WIDTH] : ping_storage_data_458 ^ i_input_data[227 % IN_WIDTH];
                662 / IN_WIDTH: ping_storage_data_458 <= (fillup_transition == 1'b1) ? i_input_data[662 % IN_WIDTH] : ping_storage_data_458 ^ i_input_data[662 % IN_WIDTH];
                897 / IN_WIDTH: ping_storage_data_458 <= (fillup_transition == 1'b1) ? i_input_data[897 % IN_WIDTH] : ping_storage_data_458 ^ i_input_data[897 % IN_WIDTH];
                962 / IN_WIDTH: ping_storage_data_458 <= (fillup_transition == 1'b1) ? i_input_data[962 % IN_WIDTH] : ping_storage_data_458 ^ i_input_data[962 % IN_WIDTH];
                default: ping_storage_data_458 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_458;
                endcase
            end else begin
                case (input_count)
                227 / IN_WIDTH: pong_storage_data_458 <= (fillup_transition == 1'b1) ? i_input_data[227 % IN_WIDTH] : pong_storage_data_458 ^ i_input_data[227 % IN_WIDTH];
                662 / IN_WIDTH: pong_storage_data_458 <= (fillup_transition == 1'b1) ? i_input_data[662 % IN_WIDTH] : pong_storage_data_458 ^ i_input_data[662 % IN_WIDTH];
                897 / IN_WIDTH: pong_storage_data_458 <= (fillup_transition == 1'b1) ? i_input_data[897 % IN_WIDTH] : pong_storage_data_458 ^ i_input_data[897 % IN_WIDTH];
                962 / IN_WIDTH: pong_storage_data_458 <= (fillup_transition == 1'b1) ? i_input_data[962 % IN_WIDTH] : pong_storage_data_458 ^ i_input_data[962 % IN_WIDTH];
                default: pong_storage_data_458 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_458;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_458 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_458;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_458 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_458;
            end
        end
    end
end

logic ping_storage_data_459;
logic pong_storage_data_459;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_459 <= 1'b0;
        pong_storage_data_459 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                228 / IN_WIDTH: ping_storage_data_459 <= (fillup_transition == 1'b1) ? i_input_data[228 % IN_WIDTH] : ping_storage_data_459 ^ i_input_data[228 % IN_WIDTH];
                663 / IN_WIDTH: ping_storage_data_459 <= (fillup_transition == 1'b1) ? i_input_data[663 % IN_WIDTH] : ping_storage_data_459 ^ i_input_data[663 % IN_WIDTH];
                898 / IN_WIDTH: ping_storage_data_459 <= (fillup_transition == 1'b1) ? i_input_data[898 % IN_WIDTH] : ping_storage_data_459 ^ i_input_data[898 % IN_WIDTH];
                963 / IN_WIDTH: ping_storage_data_459 <= (fillup_transition == 1'b1) ? i_input_data[963 % IN_WIDTH] : ping_storage_data_459 ^ i_input_data[963 % IN_WIDTH];
                default: ping_storage_data_459 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_459;
                endcase
            end else begin
                case (input_count)
                228 / IN_WIDTH: pong_storage_data_459 <= (fillup_transition == 1'b1) ? i_input_data[228 % IN_WIDTH] : pong_storage_data_459 ^ i_input_data[228 % IN_WIDTH];
                663 / IN_WIDTH: pong_storage_data_459 <= (fillup_transition == 1'b1) ? i_input_data[663 % IN_WIDTH] : pong_storage_data_459 ^ i_input_data[663 % IN_WIDTH];
                898 / IN_WIDTH: pong_storage_data_459 <= (fillup_transition == 1'b1) ? i_input_data[898 % IN_WIDTH] : pong_storage_data_459 ^ i_input_data[898 % IN_WIDTH];
                963 / IN_WIDTH: pong_storage_data_459 <= (fillup_transition == 1'b1) ? i_input_data[963 % IN_WIDTH] : pong_storage_data_459 ^ i_input_data[963 % IN_WIDTH];
                default: pong_storage_data_459 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_459;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_459 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_459;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_459 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_459;
            end
        end
    end
end

logic ping_storage_data_460;
logic pong_storage_data_460;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_460 <= 1'b0;
        pong_storage_data_460 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                229 / IN_WIDTH: ping_storage_data_460 <= (fillup_transition == 1'b1) ? i_input_data[229 % IN_WIDTH] : ping_storage_data_460 ^ i_input_data[229 % IN_WIDTH];
                664 / IN_WIDTH: ping_storage_data_460 <= (fillup_transition == 1'b1) ? i_input_data[664 % IN_WIDTH] : ping_storage_data_460 ^ i_input_data[664 % IN_WIDTH];
                899 / IN_WIDTH: ping_storage_data_460 <= (fillup_transition == 1'b1) ? i_input_data[899 % IN_WIDTH] : ping_storage_data_460 ^ i_input_data[899 % IN_WIDTH];
                964 / IN_WIDTH: ping_storage_data_460 <= (fillup_transition == 1'b1) ? i_input_data[964 % IN_WIDTH] : ping_storage_data_460 ^ i_input_data[964 % IN_WIDTH];
                default: ping_storage_data_460 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_460;
                endcase
            end else begin
                case (input_count)
                229 / IN_WIDTH: pong_storage_data_460 <= (fillup_transition == 1'b1) ? i_input_data[229 % IN_WIDTH] : pong_storage_data_460 ^ i_input_data[229 % IN_WIDTH];
                664 / IN_WIDTH: pong_storage_data_460 <= (fillup_transition == 1'b1) ? i_input_data[664 % IN_WIDTH] : pong_storage_data_460 ^ i_input_data[664 % IN_WIDTH];
                899 / IN_WIDTH: pong_storage_data_460 <= (fillup_transition == 1'b1) ? i_input_data[899 % IN_WIDTH] : pong_storage_data_460 ^ i_input_data[899 % IN_WIDTH];
                964 / IN_WIDTH: pong_storage_data_460 <= (fillup_transition == 1'b1) ? i_input_data[964 % IN_WIDTH] : pong_storage_data_460 ^ i_input_data[964 % IN_WIDTH];
                default: pong_storage_data_460 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_460;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_460 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_460;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_460 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_460;
            end
        end
    end
end

logic ping_storage_data_461;
logic pong_storage_data_461;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_461 <= 1'b0;
        pong_storage_data_461 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                230 / IN_WIDTH: ping_storage_data_461 <= (fillup_transition == 1'b1) ? i_input_data[230 % IN_WIDTH] : ping_storage_data_461 ^ i_input_data[230 % IN_WIDTH];
                665 / IN_WIDTH: ping_storage_data_461 <= (fillup_transition == 1'b1) ? i_input_data[665 % IN_WIDTH] : ping_storage_data_461 ^ i_input_data[665 % IN_WIDTH];
                900 / IN_WIDTH: ping_storage_data_461 <= (fillup_transition == 1'b1) ? i_input_data[900 % IN_WIDTH] : ping_storage_data_461 ^ i_input_data[900 % IN_WIDTH];
                965 / IN_WIDTH: ping_storage_data_461 <= (fillup_transition == 1'b1) ? i_input_data[965 % IN_WIDTH] : ping_storage_data_461 ^ i_input_data[965 % IN_WIDTH];
                default: ping_storage_data_461 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_461;
                endcase
            end else begin
                case (input_count)
                230 / IN_WIDTH: pong_storage_data_461 <= (fillup_transition == 1'b1) ? i_input_data[230 % IN_WIDTH] : pong_storage_data_461 ^ i_input_data[230 % IN_WIDTH];
                665 / IN_WIDTH: pong_storage_data_461 <= (fillup_transition == 1'b1) ? i_input_data[665 % IN_WIDTH] : pong_storage_data_461 ^ i_input_data[665 % IN_WIDTH];
                900 / IN_WIDTH: pong_storage_data_461 <= (fillup_transition == 1'b1) ? i_input_data[900 % IN_WIDTH] : pong_storage_data_461 ^ i_input_data[900 % IN_WIDTH];
                965 / IN_WIDTH: pong_storage_data_461 <= (fillup_transition == 1'b1) ? i_input_data[965 % IN_WIDTH] : pong_storage_data_461 ^ i_input_data[965 % IN_WIDTH];
                default: pong_storage_data_461 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_461;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_461 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_461;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_461 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_461;
            end
        end
    end
end

logic ping_storage_data_462;
logic pong_storage_data_462;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_462 <= 1'b0;
        pong_storage_data_462 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                231 / IN_WIDTH: ping_storage_data_462 <= (fillup_transition == 1'b1) ? i_input_data[231 % IN_WIDTH] : ping_storage_data_462 ^ i_input_data[231 % IN_WIDTH];
                666 / IN_WIDTH: ping_storage_data_462 <= (fillup_transition == 1'b1) ? i_input_data[666 % IN_WIDTH] : ping_storage_data_462 ^ i_input_data[666 % IN_WIDTH];
                901 / IN_WIDTH: ping_storage_data_462 <= (fillup_transition == 1'b1) ? i_input_data[901 % IN_WIDTH] : ping_storage_data_462 ^ i_input_data[901 % IN_WIDTH];
                966 / IN_WIDTH: ping_storage_data_462 <= (fillup_transition == 1'b1) ? i_input_data[966 % IN_WIDTH] : ping_storage_data_462 ^ i_input_data[966 % IN_WIDTH];
                default: ping_storage_data_462 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_462;
                endcase
            end else begin
                case (input_count)
                231 / IN_WIDTH: pong_storage_data_462 <= (fillup_transition == 1'b1) ? i_input_data[231 % IN_WIDTH] : pong_storage_data_462 ^ i_input_data[231 % IN_WIDTH];
                666 / IN_WIDTH: pong_storage_data_462 <= (fillup_transition == 1'b1) ? i_input_data[666 % IN_WIDTH] : pong_storage_data_462 ^ i_input_data[666 % IN_WIDTH];
                901 / IN_WIDTH: pong_storage_data_462 <= (fillup_transition == 1'b1) ? i_input_data[901 % IN_WIDTH] : pong_storage_data_462 ^ i_input_data[901 % IN_WIDTH];
                966 / IN_WIDTH: pong_storage_data_462 <= (fillup_transition == 1'b1) ? i_input_data[966 % IN_WIDTH] : pong_storage_data_462 ^ i_input_data[966 % IN_WIDTH];
                default: pong_storage_data_462 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_462;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_462 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_462;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_462 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_462;
            end
        end
    end
end

logic ping_storage_data_463;
logic pong_storage_data_463;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_463 <= 1'b0;
        pong_storage_data_463 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                232 / IN_WIDTH: ping_storage_data_463 <= (fillup_transition == 1'b1) ? i_input_data[232 % IN_WIDTH] : ping_storage_data_463 ^ i_input_data[232 % IN_WIDTH];
                667 / IN_WIDTH: ping_storage_data_463 <= (fillup_transition == 1'b1) ? i_input_data[667 % IN_WIDTH] : ping_storage_data_463 ^ i_input_data[667 % IN_WIDTH];
                902 / IN_WIDTH: ping_storage_data_463 <= (fillup_transition == 1'b1) ? i_input_data[902 % IN_WIDTH] : ping_storage_data_463 ^ i_input_data[902 % IN_WIDTH];
                967 / IN_WIDTH: ping_storage_data_463 <= (fillup_transition == 1'b1) ? i_input_data[967 % IN_WIDTH] : ping_storage_data_463 ^ i_input_data[967 % IN_WIDTH];
                default: ping_storage_data_463 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_463;
                endcase
            end else begin
                case (input_count)
                232 / IN_WIDTH: pong_storage_data_463 <= (fillup_transition == 1'b1) ? i_input_data[232 % IN_WIDTH] : pong_storage_data_463 ^ i_input_data[232 % IN_WIDTH];
                667 / IN_WIDTH: pong_storage_data_463 <= (fillup_transition == 1'b1) ? i_input_data[667 % IN_WIDTH] : pong_storage_data_463 ^ i_input_data[667 % IN_WIDTH];
                902 / IN_WIDTH: pong_storage_data_463 <= (fillup_transition == 1'b1) ? i_input_data[902 % IN_WIDTH] : pong_storage_data_463 ^ i_input_data[902 % IN_WIDTH];
                967 / IN_WIDTH: pong_storage_data_463 <= (fillup_transition == 1'b1) ? i_input_data[967 % IN_WIDTH] : pong_storage_data_463 ^ i_input_data[967 % IN_WIDTH];
                default: pong_storage_data_463 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_463;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_463 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_463;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_463 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_463;
            end
        end
    end
end

logic ping_storage_data_464;
logic pong_storage_data_464;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_464 <= 1'b0;
        pong_storage_data_464 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                233 / IN_WIDTH: ping_storage_data_464 <= (fillup_transition == 1'b1) ? i_input_data[233 % IN_WIDTH] : ping_storage_data_464 ^ i_input_data[233 % IN_WIDTH];
                668 / IN_WIDTH: ping_storage_data_464 <= (fillup_transition == 1'b1) ? i_input_data[668 % IN_WIDTH] : ping_storage_data_464 ^ i_input_data[668 % IN_WIDTH];
                903 / IN_WIDTH: ping_storage_data_464 <= (fillup_transition == 1'b1) ? i_input_data[903 % IN_WIDTH] : ping_storage_data_464 ^ i_input_data[903 % IN_WIDTH];
                968 / IN_WIDTH: ping_storage_data_464 <= (fillup_transition == 1'b1) ? i_input_data[968 % IN_WIDTH] : ping_storage_data_464 ^ i_input_data[968 % IN_WIDTH];
                default: ping_storage_data_464 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_464;
                endcase
            end else begin
                case (input_count)
                233 / IN_WIDTH: pong_storage_data_464 <= (fillup_transition == 1'b1) ? i_input_data[233 % IN_WIDTH] : pong_storage_data_464 ^ i_input_data[233 % IN_WIDTH];
                668 / IN_WIDTH: pong_storage_data_464 <= (fillup_transition == 1'b1) ? i_input_data[668 % IN_WIDTH] : pong_storage_data_464 ^ i_input_data[668 % IN_WIDTH];
                903 / IN_WIDTH: pong_storage_data_464 <= (fillup_transition == 1'b1) ? i_input_data[903 % IN_WIDTH] : pong_storage_data_464 ^ i_input_data[903 % IN_WIDTH];
                968 / IN_WIDTH: pong_storage_data_464 <= (fillup_transition == 1'b1) ? i_input_data[968 % IN_WIDTH] : pong_storage_data_464 ^ i_input_data[968 % IN_WIDTH];
                default: pong_storage_data_464 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_464;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_464 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_464;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_464 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_464;
            end
        end
    end
end

logic ping_storage_data_465;
logic pong_storage_data_465;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_465 <= 1'b0;
        pong_storage_data_465 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                234 / IN_WIDTH: ping_storage_data_465 <= (fillup_transition == 1'b1) ? i_input_data[234 % IN_WIDTH] : ping_storage_data_465 ^ i_input_data[234 % IN_WIDTH];
                669 / IN_WIDTH: ping_storage_data_465 <= (fillup_transition == 1'b1) ? i_input_data[669 % IN_WIDTH] : ping_storage_data_465 ^ i_input_data[669 % IN_WIDTH];
                904 / IN_WIDTH: ping_storage_data_465 <= (fillup_transition == 1'b1) ? i_input_data[904 % IN_WIDTH] : ping_storage_data_465 ^ i_input_data[904 % IN_WIDTH];
                969 / IN_WIDTH: ping_storage_data_465 <= (fillup_transition == 1'b1) ? i_input_data[969 % IN_WIDTH] : ping_storage_data_465 ^ i_input_data[969 % IN_WIDTH];
                default: ping_storage_data_465 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_465;
                endcase
            end else begin
                case (input_count)
                234 / IN_WIDTH: pong_storage_data_465 <= (fillup_transition == 1'b1) ? i_input_data[234 % IN_WIDTH] : pong_storage_data_465 ^ i_input_data[234 % IN_WIDTH];
                669 / IN_WIDTH: pong_storage_data_465 <= (fillup_transition == 1'b1) ? i_input_data[669 % IN_WIDTH] : pong_storage_data_465 ^ i_input_data[669 % IN_WIDTH];
                904 / IN_WIDTH: pong_storage_data_465 <= (fillup_transition == 1'b1) ? i_input_data[904 % IN_WIDTH] : pong_storage_data_465 ^ i_input_data[904 % IN_WIDTH];
                969 / IN_WIDTH: pong_storage_data_465 <= (fillup_transition == 1'b1) ? i_input_data[969 % IN_WIDTH] : pong_storage_data_465 ^ i_input_data[969 % IN_WIDTH];
                default: pong_storage_data_465 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_465;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_465 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_465;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_465 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_465;
            end
        end
    end
end

logic ping_storage_data_466;
logic pong_storage_data_466;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_466 <= 1'b0;
        pong_storage_data_466 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                235 / IN_WIDTH: ping_storage_data_466 <= (fillup_transition == 1'b1) ? i_input_data[235 % IN_WIDTH] : ping_storage_data_466 ^ i_input_data[235 % IN_WIDTH];
                670 / IN_WIDTH: ping_storage_data_466 <= (fillup_transition == 1'b1) ? i_input_data[670 % IN_WIDTH] : ping_storage_data_466 ^ i_input_data[670 % IN_WIDTH];
                905 / IN_WIDTH: ping_storage_data_466 <= (fillup_transition == 1'b1) ? i_input_data[905 % IN_WIDTH] : ping_storage_data_466 ^ i_input_data[905 % IN_WIDTH];
                970 / IN_WIDTH: ping_storage_data_466 <= (fillup_transition == 1'b1) ? i_input_data[970 % IN_WIDTH] : ping_storage_data_466 ^ i_input_data[970 % IN_WIDTH];
                default: ping_storage_data_466 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_466;
                endcase
            end else begin
                case (input_count)
                235 / IN_WIDTH: pong_storage_data_466 <= (fillup_transition == 1'b1) ? i_input_data[235 % IN_WIDTH] : pong_storage_data_466 ^ i_input_data[235 % IN_WIDTH];
                670 / IN_WIDTH: pong_storage_data_466 <= (fillup_transition == 1'b1) ? i_input_data[670 % IN_WIDTH] : pong_storage_data_466 ^ i_input_data[670 % IN_WIDTH];
                905 / IN_WIDTH: pong_storage_data_466 <= (fillup_transition == 1'b1) ? i_input_data[905 % IN_WIDTH] : pong_storage_data_466 ^ i_input_data[905 % IN_WIDTH];
                970 / IN_WIDTH: pong_storage_data_466 <= (fillup_transition == 1'b1) ? i_input_data[970 % IN_WIDTH] : pong_storage_data_466 ^ i_input_data[970 % IN_WIDTH];
                default: pong_storage_data_466 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_466;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_466 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_466;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_466 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_466;
            end
        end
    end
end

logic ping_storage_data_467;
logic pong_storage_data_467;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_467 <= 1'b0;
        pong_storage_data_467 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                236 / IN_WIDTH: ping_storage_data_467 <= (fillup_transition == 1'b1) ? i_input_data[236 % IN_WIDTH] : ping_storage_data_467 ^ i_input_data[236 % IN_WIDTH];
                671 / IN_WIDTH: ping_storage_data_467 <= (fillup_transition == 1'b1) ? i_input_data[671 % IN_WIDTH] : ping_storage_data_467 ^ i_input_data[671 % IN_WIDTH];
                906 / IN_WIDTH: ping_storage_data_467 <= (fillup_transition == 1'b1) ? i_input_data[906 % IN_WIDTH] : ping_storage_data_467 ^ i_input_data[906 % IN_WIDTH];
                971 / IN_WIDTH: ping_storage_data_467 <= (fillup_transition == 1'b1) ? i_input_data[971 % IN_WIDTH] : ping_storage_data_467 ^ i_input_data[971 % IN_WIDTH];
                default: ping_storage_data_467 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_467;
                endcase
            end else begin
                case (input_count)
                236 / IN_WIDTH: pong_storage_data_467 <= (fillup_transition == 1'b1) ? i_input_data[236 % IN_WIDTH] : pong_storage_data_467 ^ i_input_data[236 % IN_WIDTH];
                671 / IN_WIDTH: pong_storage_data_467 <= (fillup_transition == 1'b1) ? i_input_data[671 % IN_WIDTH] : pong_storage_data_467 ^ i_input_data[671 % IN_WIDTH];
                906 / IN_WIDTH: pong_storage_data_467 <= (fillup_transition == 1'b1) ? i_input_data[906 % IN_WIDTH] : pong_storage_data_467 ^ i_input_data[906 % IN_WIDTH];
                971 / IN_WIDTH: pong_storage_data_467 <= (fillup_transition == 1'b1) ? i_input_data[971 % IN_WIDTH] : pong_storage_data_467 ^ i_input_data[971 % IN_WIDTH];
                default: pong_storage_data_467 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_467;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_467 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_467;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_467 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_467;
            end
        end
    end
end

logic ping_storage_data_468;
logic pong_storage_data_468;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_468 <= 1'b0;
        pong_storage_data_468 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                237 / IN_WIDTH: ping_storage_data_468 <= (fillup_transition == 1'b1) ? i_input_data[237 % IN_WIDTH] : ping_storage_data_468 ^ i_input_data[237 % IN_WIDTH];
                576 / IN_WIDTH: ping_storage_data_468 <= (fillup_transition == 1'b1) ? i_input_data[576 % IN_WIDTH] : ping_storage_data_468 ^ i_input_data[576 % IN_WIDTH];
                907 / IN_WIDTH: ping_storage_data_468 <= (fillup_transition == 1'b1) ? i_input_data[907 % IN_WIDTH] : ping_storage_data_468 ^ i_input_data[907 % IN_WIDTH];
                972 / IN_WIDTH: ping_storage_data_468 <= (fillup_transition == 1'b1) ? i_input_data[972 % IN_WIDTH] : ping_storage_data_468 ^ i_input_data[972 % IN_WIDTH];
                default: ping_storage_data_468 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_468;
                endcase
            end else begin
                case (input_count)
                237 / IN_WIDTH: pong_storage_data_468 <= (fillup_transition == 1'b1) ? i_input_data[237 % IN_WIDTH] : pong_storage_data_468 ^ i_input_data[237 % IN_WIDTH];
                576 / IN_WIDTH: pong_storage_data_468 <= (fillup_transition == 1'b1) ? i_input_data[576 % IN_WIDTH] : pong_storage_data_468 ^ i_input_data[576 % IN_WIDTH];
                907 / IN_WIDTH: pong_storage_data_468 <= (fillup_transition == 1'b1) ? i_input_data[907 % IN_WIDTH] : pong_storage_data_468 ^ i_input_data[907 % IN_WIDTH];
                972 / IN_WIDTH: pong_storage_data_468 <= (fillup_transition == 1'b1) ? i_input_data[972 % IN_WIDTH] : pong_storage_data_468 ^ i_input_data[972 % IN_WIDTH];
                default: pong_storage_data_468 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_468;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_468 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_468;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_468 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_468;
            end
        end
    end
end

logic ping_storage_data_469;
logic pong_storage_data_469;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_469 <= 1'b0;
        pong_storage_data_469 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                238 / IN_WIDTH: ping_storage_data_469 <= (fillup_transition == 1'b1) ? i_input_data[238 % IN_WIDTH] : ping_storage_data_469 ^ i_input_data[238 % IN_WIDTH];
                577 / IN_WIDTH: ping_storage_data_469 <= (fillup_transition == 1'b1) ? i_input_data[577 % IN_WIDTH] : ping_storage_data_469 ^ i_input_data[577 % IN_WIDTH];
                908 / IN_WIDTH: ping_storage_data_469 <= (fillup_transition == 1'b1) ? i_input_data[908 % IN_WIDTH] : ping_storage_data_469 ^ i_input_data[908 % IN_WIDTH];
                973 / IN_WIDTH: ping_storage_data_469 <= (fillup_transition == 1'b1) ? i_input_data[973 % IN_WIDTH] : ping_storage_data_469 ^ i_input_data[973 % IN_WIDTH];
                default: ping_storage_data_469 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_469;
                endcase
            end else begin
                case (input_count)
                238 / IN_WIDTH: pong_storage_data_469 <= (fillup_transition == 1'b1) ? i_input_data[238 % IN_WIDTH] : pong_storage_data_469 ^ i_input_data[238 % IN_WIDTH];
                577 / IN_WIDTH: pong_storage_data_469 <= (fillup_transition == 1'b1) ? i_input_data[577 % IN_WIDTH] : pong_storage_data_469 ^ i_input_data[577 % IN_WIDTH];
                908 / IN_WIDTH: pong_storage_data_469 <= (fillup_transition == 1'b1) ? i_input_data[908 % IN_WIDTH] : pong_storage_data_469 ^ i_input_data[908 % IN_WIDTH];
                973 / IN_WIDTH: pong_storage_data_469 <= (fillup_transition == 1'b1) ? i_input_data[973 % IN_WIDTH] : pong_storage_data_469 ^ i_input_data[973 % IN_WIDTH];
                default: pong_storage_data_469 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_469;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_469 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_469;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_469 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_469;
            end
        end
    end
end

logic ping_storage_data_470;
logic pong_storage_data_470;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_470 <= 1'b0;
        pong_storage_data_470 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                239 / IN_WIDTH: ping_storage_data_470 <= (fillup_transition == 1'b1) ? i_input_data[239 % IN_WIDTH] : ping_storage_data_470 ^ i_input_data[239 % IN_WIDTH];
                578 / IN_WIDTH: ping_storage_data_470 <= (fillup_transition == 1'b1) ? i_input_data[578 % IN_WIDTH] : ping_storage_data_470 ^ i_input_data[578 % IN_WIDTH];
                909 / IN_WIDTH: ping_storage_data_470 <= (fillup_transition == 1'b1) ? i_input_data[909 % IN_WIDTH] : ping_storage_data_470 ^ i_input_data[909 % IN_WIDTH];
                974 / IN_WIDTH: ping_storage_data_470 <= (fillup_transition == 1'b1) ? i_input_data[974 % IN_WIDTH] : ping_storage_data_470 ^ i_input_data[974 % IN_WIDTH];
                default: ping_storage_data_470 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_470;
                endcase
            end else begin
                case (input_count)
                239 / IN_WIDTH: pong_storage_data_470 <= (fillup_transition == 1'b1) ? i_input_data[239 % IN_WIDTH] : pong_storage_data_470 ^ i_input_data[239 % IN_WIDTH];
                578 / IN_WIDTH: pong_storage_data_470 <= (fillup_transition == 1'b1) ? i_input_data[578 % IN_WIDTH] : pong_storage_data_470 ^ i_input_data[578 % IN_WIDTH];
                909 / IN_WIDTH: pong_storage_data_470 <= (fillup_transition == 1'b1) ? i_input_data[909 % IN_WIDTH] : pong_storage_data_470 ^ i_input_data[909 % IN_WIDTH];
                974 / IN_WIDTH: pong_storage_data_470 <= (fillup_transition == 1'b1) ? i_input_data[974 % IN_WIDTH] : pong_storage_data_470 ^ i_input_data[974 % IN_WIDTH];
                default: pong_storage_data_470 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_470;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_470 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_470;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_470 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_470;
            end
        end
    end
end

logic ping_storage_data_471;
logic pong_storage_data_471;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_471 <= 1'b0;
        pong_storage_data_471 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                240 / IN_WIDTH: ping_storage_data_471 <= (fillup_transition == 1'b1) ? i_input_data[240 % IN_WIDTH] : ping_storage_data_471 ^ i_input_data[240 % IN_WIDTH];
                579 / IN_WIDTH: ping_storage_data_471 <= (fillup_transition == 1'b1) ? i_input_data[579 % IN_WIDTH] : ping_storage_data_471 ^ i_input_data[579 % IN_WIDTH];
                910 / IN_WIDTH: ping_storage_data_471 <= (fillup_transition == 1'b1) ? i_input_data[910 % IN_WIDTH] : ping_storage_data_471 ^ i_input_data[910 % IN_WIDTH];
                975 / IN_WIDTH: ping_storage_data_471 <= (fillup_transition == 1'b1) ? i_input_data[975 % IN_WIDTH] : ping_storage_data_471 ^ i_input_data[975 % IN_WIDTH];
                default: ping_storage_data_471 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_471;
                endcase
            end else begin
                case (input_count)
                240 / IN_WIDTH: pong_storage_data_471 <= (fillup_transition == 1'b1) ? i_input_data[240 % IN_WIDTH] : pong_storage_data_471 ^ i_input_data[240 % IN_WIDTH];
                579 / IN_WIDTH: pong_storage_data_471 <= (fillup_transition == 1'b1) ? i_input_data[579 % IN_WIDTH] : pong_storage_data_471 ^ i_input_data[579 % IN_WIDTH];
                910 / IN_WIDTH: pong_storage_data_471 <= (fillup_transition == 1'b1) ? i_input_data[910 % IN_WIDTH] : pong_storage_data_471 ^ i_input_data[910 % IN_WIDTH];
                975 / IN_WIDTH: pong_storage_data_471 <= (fillup_transition == 1'b1) ? i_input_data[975 % IN_WIDTH] : pong_storage_data_471 ^ i_input_data[975 % IN_WIDTH];
                default: pong_storage_data_471 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_471;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_471 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_471;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_471 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_471;
            end
        end
    end
end

logic ping_storage_data_472;
logic pong_storage_data_472;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_472 <= 1'b0;
        pong_storage_data_472 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                241 / IN_WIDTH: ping_storage_data_472 <= (fillup_transition == 1'b1) ? i_input_data[241 % IN_WIDTH] : ping_storage_data_472 ^ i_input_data[241 % IN_WIDTH];
                580 / IN_WIDTH: ping_storage_data_472 <= (fillup_transition == 1'b1) ? i_input_data[580 % IN_WIDTH] : ping_storage_data_472 ^ i_input_data[580 % IN_WIDTH];
                911 / IN_WIDTH: ping_storage_data_472 <= (fillup_transition == 1'b1) ? i_input_data[911 % IN_WIDTH] : ping_storage_data_472 ^ i_input_data[911 % IN_WIDTH];
                976 / IN_WIDTH: ping_storage_data_472 <= (fillup_transition == 1'b1) ? i_input_data[976 % IN_WIDTH] : ping_storage_data_472 ^ i_input_data[976 % IN_WIDTH];
                default: ping_storage_data_472 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_472;
                endcase
            end else begin
                case (input_count)
                241 / IN_WIDTH: pong_storage_data_472 <= (fillup_transition == 1'b1) ? i_input_data[241 % IN_WIDTH] : pong_storage_data_472 ^ i_input_data[241 % IN_WIDTH];
                580 / IN_WIDTH: pong_storage_data_472 <= (fillup_transition == 1'b1) ? i_input_data[580 % IN_WIDTH] : pong_storage_data_472 ^ i_input_data[580 % IN_WIDTH];
                911 / IN_WIDTH: pong_storage_data_472 <= (fillup_transition == 1'b1) ? i_input_data[911 % IN_WIDTH] : pong_storage_data_472 ^ i_input_data[911 % IN_WIDTH];
                976 / IN_WIDTH: pong_storage_data_472 <= (fillup_transition == 1'b1) ? i_input_data[976 % IN_WIDTH] : pong_storage_data_472 ^ i_input_data[976 % IN_WIDTH];
                default: pong_storage_data_472 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_472;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_472 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_472;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_472 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_472;
            end
        end
    end
end

logic ping_storage_data_473;
logic pong_storage_data_473;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_473 <= 1'b0;
        pong_storage_data_473 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                242 / IN_WIDTH: ping_storage_data_473 <= (fillup_transition == 1'b1) ? i_input_data[242 % IN_WIDTH] : ping_storage_data_473 ^ i_input_data[242 % IN_WIDTH];
                581 / IN_WIDTH: ping_storage_data_473 <= (fillup_transition == 1'b1) ? i_input_data[581 % IN_WIDTH] : ping_storage_data_473 ^ i_input_data[581 % IN_WIDTH];
                912 / IN_WIDTH: ping_storage_data_473 <= (fillup_transition == 1'b1) ? i_input_data[912 % IN_WIDTH] : ping_storage_data_473 ^ i_input_data[912 % IN_WIDTH];
                977 / IN_WIDTH: ping_storage_data_473 <= (fillup_transition == 1'b1) ? i_input_data[977 % IN_WIDTH] : ping_storage_data_473 ^ i_input_data[977 % IN_WIDTH];
                default: ping_storage_data_473 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_473;
                endcase
            end else begin
                case (input_count)
                242 / IN_WIDTH: pong_storage_data_473 <= (fillup_transition == 1'b1) ? i_input_data[242 % IN_WIDTH] : pong_storage_data_473 ^ i_input_data[242 % IN_WIDTH];
                581 / IN_WIDTH: pong_storage_data_473 <= (fillup_transition == 1'b1) ? i_input_data[581 % IN_WIDTH] : pong_storage_data_473 ^ i_input_data[581 % IN_WIDTH];
                912 / IN_WIDTH: pong_storage_data_473 <= (fillup_transition == 1'b1) ? i_input_data[912 % IN_WIDTH] : pong_storage_data_473 ^ i_input_data[912 % IN_WIDTH];
                977 / IN_WIDTH: pong_storage_data_473 <= (fillup_transition == 1'b1) ? i_input_data[977 % IN_WIDTH] : pong_storage_data_473 ^ i_input_data[977 % IN_WIDTH];
                default: pong_storage_data_473 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_473;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_473 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_473;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_473 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_473;
            end
        end
    end
end

logic ping_storage_data_474;
logic pong_storage_data_474;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_474 <= 1'b0;
        pong_storage_data_474 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                243 / IN_WIDTH: ping_storage_data_474 <= (fillup_transition == 1'b1) ? i_input_data[243 % IN_WIDTH] : ping_storage_data_474 ^ i_input_data[243 % IN_WIDTH];
                582 / IN_WIDTH: ping_storage_data_474 <= (fillup_transition == 1'b1) ? i_input_data[582 % IN_WIDTH] : ping_storage_data_474 ^ i_input_data[582 % IN_WIDTH];
                913 / IN_WIDTH: ping_storage_data_474 <= (fillup_transition == 1'b1) ? i_input_data[913 % IN_WIDTH] : ping_storage_data_474 ^ i_input_data[913 % IN_WIDTH];
                978 / IN_WIDTH: ping_storage_data_474 <= (fillup_transition == 1'b1) ? i_input_data[978 % IN_WIDTH] : ping_storage_data_474 ^ i_input_data[978 % IN_WIDTH];
                default: ping_storage_data_474 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_474;
                endcase
            end else begin
                case (input_count)
                243 / IN_WIDTH: pong_storage_data_474 <= (fillup_transition == 1'b1) ? i_input_data[243 % IN_WIDTH] : pong_storage_data_474 ^ i_input_data[243 % IN_WIDTH];
                582 / IN_WIDTH: pong_storage_data_474 <= (fillup_transition == 1'b1) ? i_input_data[582 % IN_WIDTH] : pong_storage_data_474 ^ i_input_data[582 % IN_WIDTH];
                913 / IN_WIDTH: pong_storage_data_474 <= (fillup_transition == 1'b1) ? i_input_data[913 % IN_WIDTH] : pong_storage_data_474 ^ i_input_data[913 % IN_WIDTH];
                978 / IN_WIDTH: pong_storage_data_474 <= (fillup_transition == 1'b1) ? i_input_data[978 % IN_WIDTH] : pong_storage_data_474 ^ i_input_data[978 % IN_WIDTH];
                default: pong_storage_data_474 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_474;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_474 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_474;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_474 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_474;
            end
        end
    end
end

logic ping_storage_data_475;
logic pong_storage_data_475;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_475 <= 1'b0;
        pong_storage_data_475 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                244 / IN_WIDTH: ping_storage_data_475 <= (fillup_transition == 1'b1) ? i_input_data[244 % IN_WIDTH] : ping_storage_data_475 ^ i_input_data[244 % IN_WIDTH];
                583 / IN_WIDTH: ping_storage_data_475 <= (fillup_transition == 1'b1) ? i_input_data[583 % IN_WIDTH] : ping_storage_data_475 ^ i_input_data[583 % IN_WIDTH];
                914 / IN_WIDTH: ping_storage_data_475 <= (fillup_transition == 1'b1) ? i_input_data[914 % IN_WIDTH] : ping_storage_data_475 ^ i_input_data[914 % IN_WIDTH];
                979 / IN_WIDTH: ping_storage_data_475 <= (fillup_transition == 1'b1) ? i_input_data[979 % IN_WIDTH] : ping_storage_data_475 ^ i_input_data[979 % IN_WIDTH];
                default: ping_storage_data_475 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_475;
                endcase
            end else begin
                case (input_count)
                244 / IN_WIDTH: pong_storage_data_475 <= (fillup_transition == 1'b1) ? i_input_data[244 % IN_WIDTH] : pong_storage_data_475 ^ i_input_data[244 % IN_WIDTH];
                583 / IN_WIDTH: pong_storage_data_475 <= (fillup_transition == 1'b1) ? i_input_data[583 % IN_WIDTH] : pong_storage_data_475 ^ i_input_data[583 % IN_WIDTH];
                914 / IN_WIDTH: pong_storage_data_475 <= (fillup_transition == 1'b1) ? i_input_data[914 % IN_WIDTH] : pong_storage_data_475 ^ i_input_data[914 % IN_WIDTH];
                979 / IN_WIDTH: pong_storage_data_475 <= (fillup_transition == 1'b1) ? i_input_data[979 % IN_WIDTH] : pong_storage_data_475 ^ i_input_data[979 % IN_WIDTH];
                default: pong_storage_data_475 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_475;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_475 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_475;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_475 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_475;
            end
        end
    end
end

logic ping_storage_data_476;
logic pong_storage_data_476;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_476 <= 1'b0;
        pong_storage_data_476 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                245 / IN_WIDTH: ping_storage_data_476 <= (fillup_transition == 1'b1) ? i_input_data[245 % IN_WIDTH] : ping_storage_data_476 ^ i_input_data[245 % IN_WIDTH];
                584 / IN_WIDTH: ping_storage_data_476 <= (fillup_transition == 1'b1) ? i_input_data[584 % IN_WIDTH] : ping_storage_data_476 ^ i_input_data[584 % IN_WIDTH];
                915 / IN_WIDTH: ping_storage_data_476 <= (fillup_transition == 1'b1) ? i_input_data[915 % IN_WIDTH] : ping_storage_data_476 ^ i_input_data[915 % IN_WIDTH];
                980 / IN_WIDTH: ping_storage_data_476 <= (fillup_transition == 1'b1) ? i_input_data[980 % IN_WIDTH] : ping_storage_data_476 ^ i_input_data[980 % IN_WIDTH];
                default: ping_storage_data_476 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_476;
                endcase
            end else begin
                case (input_count)
                245 / IN_WIDTH: pong_storage_data_476 <= (fillup_transition == 1'b1) ? i_input_data[245 % IN_WIDTH] : pong_storage_data_476 ^ i_input_data[245 % IN_WIDTH];
                584 / IN_WIDTH: pong_storage_data_476 <= (fillup_transition == 1'b1) ? i_input_data[584 % IN_WIDTH] : pong_storage_data_476 ^ i_input_data[584 % IN_WIDTH];
                915 / IN_WIDTH: pong_storage_data_476 <= (fillup_transition == 1'b1) ? i_input_data[915 % IN_WIDTH] : pong_storage_data_476 ^ i_input_data[915 % IN_WIDTH];
                980 / IN_WIDTH: pong_storage_data_476 <= (fillup_transition == 1'b1) ? i_input_data[980 % IN_WIDTH] : pong_storage_data_476 ^ i_input_data[980 % IN_WIDTH];
                default: pong_storage_data_476 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_476;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_476 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_476;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_476 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_476;
            end
        end
    end
end

logic ping_storage_data_477;
logic pong_storage_data_477;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_477 <= 1'b0;
        pong_storage_data_477 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                246 / IN_WIDTH: ping_storage_data_477 <= (fillup_transition == 1'b1) ? i_input_data[246 % IN_WIDTH] : ping_storage_data_477 ^ i_input_data[246 % IN_WIDTH];
                585 / IN_WIDTH: ping_storage_data_477 <= (fillup_transition == 1'b1) ? i_input_data[585 % IN_WIDTH] : ping_storage_data_477 ^ i_input_data[585 % IN_WIDTH];
                916 / IN_WIDTH: ping_storage_data_477 <= (fillup_transition == 1'b1) ? i_input_data[916 % IN_WIDTH] : ping_storage_data_477 ^ i_input_data[916 % IN_WIDTH];
                981 / IN_WIDTH: ping_storage_data_477 <= (fillup_transition == 1'b1) ? i_input_data[981 % IN_WIDTH] : ping_storage_data_477 ^ i_input_data[981 % IN_WIDTH];
                default: ping_storage_data_477 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_477;
                endcase
            end else begin
                case (input_count)
                246 / IN_WIDTH: pong_storage_data_477 <= (fillup_transition == 1'b1) ? i_input_data[246 % IN_WIDTH] : pong_storage_data_477 ^ i_input_data[246 % IN_WIDTH];
                585 / IN_WIDTH: pong_storage_data_477 <= (fillup_transition == 1'b1) ? i_input_data[585 % IN_WIDTH] : pong_storage_data_477 ^ i_input_data[585 % IN_WIDTH];
                916 / IN_WIDTH: pong_storage_data_477 <= (fillup_transition == 1'b1) ? i_input_data[916 % IN_WIDTH] : pong_storage_data_477 ^ i_input_data[916 % IN_WIDTH];
                981 / IN_WIDTH: pong_storage_data_477 <= (fillup_transition == 1'b1) ? i_input_data[981 % IN_WIDTH] : pong_storage_data_477 ^ i_input_data[981 % IN_WIDTH];
                default: pong_storage_data_477 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_477;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_477 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_477;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_477 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_477;
            end
        end
    end
end

logic ping_storage_data_478;
logic pong_storage_data_478;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_478 <= 1'b0;
        pong_storage_data_478 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                247 / IN_WIDTH: ping_storage_data_478 <= (fillup_transition == 1'b1) ? i_input_data[247 % IN_WIDTH] : ping_storage_data_478 ^ i_input_data[247 % IN_WIDTH];
                586 / IN_WIDTH: ping_storage_data_478 <= (fillup_transition == 1'b1) ? i_input_data[586 % IN_WIDTH] : ping_storage_data_478 ^ i_input_data[586 % IN_WIDTH];
                917 / IN_WIDTH: ping_storage_data_478 <= (fillup_transition == 1'b1) ? i_input_data[917 % IN_WIDTH] : ping_storage_data_478 ^ i_input_data[917 % IN_WIDTH];
                982 / IN_WIDTH: ping_storage_data_478 <= (fillup_transition == 1'b1) ? i_input_data[982 % IN_WIDTH] : ping_storage_data_478 ^ i_input_data[982 % IN_WIDTH];
                default: ping_storage_data_478 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_478;
                endcase
            end else begin
                case (input_count)
                247 / IN_WIDTH: pong_storage_data_478 <= (fillup_transition == 1'b1) ? i_input_data[247 % IN_WIDTH] : pong_storage_data_478 ^ i_input_data[247 % IN_WIDTH];
                586 / IN_WIDTH: pong_storage_data_478 <= (fillup_transition == 1'b1) ? i_input_data[586 % IN_WIDTH] : pong_storage_data_478 ^ i_input_data[586 % IN_WIDTH];
                917 / IN_WIDTH: pong_storage_data_478 <= (fillup_transition == 1'b1) ? i_input_data[917 % IN_WIDTH] : pong_storage_data_478 ^ i_input_data[917 % IN_WIDTH];
                982 / IN_WIDTH: pong_storage_data_478 <= (fillup_transition == 1'b1) ? i_input_data[982 % IN_WIDTH] : pong_storage_data_478 ^ i_input_data[982 % IN_WIDTH];
                default: pong_storage_data_478 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_478;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_478 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_478;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_478 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_478;
            end
        end
    end
end

logic ping_storage_data_479;
logic pong_storage_data_479;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_479 <= 1'b0;
        pong_storage_data_479 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                248 / IN_WIDTH: ping_storage_data_479 <= (fillup_transition == 1'b1) ? i_input_data[248 % IN_WIDTH] : ping_storage_data_479 ^ i_input_data[248 % IN_WIDTH];
                587 / IN_WIDTH: ping_storage_data_479 <= (fillup_transition == 1'b1) ? i_input_data[587 % IN_WIDTH] : ping_storage_data_479 ^ i_input_data[587 % IN_WIDTH];
                918 / IN_WIDTH: ping_storage_data_479 <= (fillup_transition == 1'b1) ? i_input_data[918 % IN_WIDTH] : ping_storage_data_479 ^ i_input_data[918 % IN_WIDTH];
                983 / IN_WIDTH: ping_storage_data_479 <= (fillup_transition == 1'b1) ? i_input_data[983 % IN_WIDTH] : ping_storage_data_479 ^ i_input_data[983 % IN_WIDTH];
                default: ping_storage_data_479 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_479;
                endcase
            end else begin
                case (input_count)
                248 / IN_WIDTH: pong_storage_data_479 <= (fillup_transition == 1'b1) ? i_input_data[248 % IN_WIDTH] : pong_storage_data_479 ^ i_input_data[248 % IN_WIDTH];
                587 / IN_WIDTH: pong_storage_data_479 <= (fillup_transition == 1'b1) ? i_input_data[587 % IN_WIDTH] : pong_storage_data_479 ^ i_input_data[587 % IN_WIDTH];
                918 / IN_WIDTH: pong_storage_data_479 <= (fillup_transition == 1'b1) ? i_input_data[918 % IN_WIDTH] : pong_storage_data_479 ^ i_input_data[918 % IN_WIDTH];
                983 / IN_WIDTH: pong_storage_data_479 <= (fillup_transition == 1'b1) ? i_input_data[983 % IN_WIDTH] : pong_storage_data_479 ^ i_input_data[983 % IN_WIDTH];
                default: pong_storage_data_479 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_479;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_479 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_479;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_479 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_479;
            end
        end
    end
end

logic ping_storage_data_480;
logic pong_storage_data_480;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_480 <= 1'b0;
        pong_storage_data_480 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                434 / IN_WIDTH: ping_storage_data_480 <= (fillup_transition == 1'b1) ? i_input_data[434 % IN_WIDTH] : ping_storage_data_480 ^ i_input_data[434 % IN_WIDTH];
                536 / IN_WIDTH: ping_storage_data_480 <= (fillup_transition == 1'b1) ? i_input_data[536 % IN_WIDTH] : ping_storage_data_480 ^ i_input_data[536 % IN_WIDTH];
                686 / IN_WIDTH: ping_storage_data_480 <= (fillup_transition == 1'b1) ? i_input_data[686 % IN_WIDTH] : ping_storage_data_480 ^ i_input_data[686 % IN_WIDTH];
                1073 / IN_WIDTH: ping_storage_data_480 <= (fillup_transition == 1'b1) ? i_input_data[1073 % IN_WIDTH] : ping_storage_data_480 ^ i_input_data[1073 % IN_WIDTH];
                default: ping_storage_data_480 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_480;
                endcase
            end else begin
                case (input_count)
                434 / IN_WIDTH: pong_storage_data_480 <= (fillup_transition == 1'b1) ? i_input_data[434 % IN_WIDTH] : pong_storage_data_480 ^ i_input_data[434 % IN_WIDTH];
                536 / IN_WIDTH: pong_storage_data_480 <= (fillup_transition == 1'b1) ? i_input_data[536 % IN_WIDTH] : pong_storage_data_480 ^ i_input_data[536 % IN_WIDTH];
                686 / IN_WIDTH: pong_storage_data_480 <= (fillup_transition == 1'b1) ? i_input_data[686 % IN_WIDTH] : pong_storage_data_480 ^ i_input_data[686 % IN_WIDTH];
                1073 / IN_WIDTH: pong_storage_data_480 <= (fillup_transition == 1'b1) ? i_input_data[1073 % IN_WIDTH] : pong_storage_data_480 ^ i_input_data[1073 % IN_WIDTH];
                default: pong_storage_data_480 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_480;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_480 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_480;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_480 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_480;
            end
        end
    end
end

logic ping_storage_data_481;
logic pong_storage_data_481;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_481 <= 1'b0;
        pong_storage_data_481 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                435 / IN_WIDTH: ping_storage_data_481 <= (fillup_transition == 1'b1) ? i_input_data[435 % IN_WIDTH] : ping_storage_data_481 ^ i_input_data[435 % IN_WIDTH];
                537 / IN_WIDTH: ping_storage_data_481 <= (fillup_transition == 1'b1) ? i_input_data[537 % IN_WIDTH] : ping_storage_data_481 ^ i_input_data[537 % IN_WIDTH];
                687 / IN_WIDTH: ping_storage_data_481 <= (fillup_transition == 1'b1) ? i_input_data[687 % IN_WIDTH] : ping_storage_data_481 ^ i_input_data[687 % IN_WIDTH];
                1074 / IN_WIDTH: ping_storage_data_481 <= (fillup_transition == 1'b1) ? i_input_data[1074 % IN_WIDTH] : ping_storage_data_481 ^ i_input_data[1074 % IN_WIDTH];
                default: ping_storage_data_481 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_481;
                endcase
            end else begin
                case (input_count)
                435 / IN_WIDTH: pong_storage_data_481 <= (fillup_transition == 1'b1) ? i_input_data[435 % IN_WIDTH] : pong_storage_data_481 ^ i_input_data[435 % IN_WIDTH];
                537 / IN_WIDTH: pong_storage_data_481 <= (fillup_transition == 1'b1) ? i_input_data[537 % IN_WIDTH] : pong_storage_data_481 ^ i_input_data[537 % IN_WIDTH];
                687 / IN_WIDTH: pong_storage_data_481 <= (fillup_transition == 1'b1) ? i_input_data[687 % IN_WIDTH] : pong_storage_data_481 ^ i_input_data[687 % IN_WIDTH];
                1074 / IN_WIDTH: pong_storage_data_481 <= (fillup_transition == 1'b1) ? i_input_data[1074 % IN_WIDTH] : pong_storage_data_481 ^ i_input_data[1074 % IN_WIDTH];
                default: pong_storage_data_481 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_481;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_481 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_481;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_481 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_481;
            end
        end
    end
end

logic ping_storage_data_482;
logic pong_storage_data_482;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_482 <= 1'b0;
        pong_storage_data_482 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                436 / IN_WIDTH: ping_storage_data_482 <= (fillup_transition == 1'b1) ? i_input_data[436 % IN_WIDTH] : ping_storage_data_482 ^ i_input_data[436 % IN_WIDTH];
                538 / IN_WIDTH: ping_storage_data_482 <= (fillup_transition == 1'b1) ? i_input_data[538 % IN_WIDTH] : ping_storage_data_482 ^ i_input_data[538 % IN_WIDTH];
                688 / IN_WIDTH: ping_storage_data_482 <= (fillup_transition == 1'b1) ? i_input_data[688 % IN_WIDTH] : ping_storage_data_482 ^ i_input_data[688 % IN_WIDTH];
                1075 / IN_WIDTH: ping_storage_data_482 <= (fillup_transition == 1'b1) ? i_input_data[1075 % IN_WIDTH] : ping_storage_data_482 ^ i_input_data[1075 % IN_WIDTH];
                default: ping_storage_data_482 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_482;
                endcase
            end else begin
                case (input_count)
                436 / IN_WIDTH: pong_storage_data_482 <= (fillup_transition == 1'b1) ? i_input_data[436 % IN_WIDTH] : pong_storage_data_482 ^ i_input_data[436 % IN_WIDTH];
                538 / IN_WIDTH: pong_storage_data_482 <= (fillup_transition == 1'b1) ? i_input_data[538 % IN_WIDTH] : pong_storage_data_482 ^ i_input_data[538 % IN_WIDTH];
                688 / IN_WIDTH: pong_storage_data_482 <= (fillup_transition == 1'b1) ? i_input_data[688 % IN_WIDTH] : pong_storage_data_482 ^ i_input_data[688 % IN_WIDTH];
                1075 / IN_WIDTH: pong_storage_data_482 <= (fillup_transition == 1'b1) ? i_input_data[1075 % IN_WIDTH] : pong_storage_data_482 ^ i_input_data[1075 % IN_WIDTH];
                default: pong_storage_data_482 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_482;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_482 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_482;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_482 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_482;
            end
        end
    end
end

logic ping_storage_data_483;
logic pong_storage_data_483;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_483 <= 1'b0;
        pong_storage_data_483 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                437 / IN_WIDTH: ping_storage_data_483 <= (fillup_transition == 1'b1) ? i_input_data[437 % IN_WIDTH] : ping_storage_data_483 ^ i_input_data[437 % IN_WIDTH];
                539 / IN_WIDTH: ping_storage_data_483 <= (fillup_transition == 1'b1) ? i_input_data[539 % IN_WIDTH] : ping_storage_data_483 ^ i_input_data[539 % IN_WIDTH];
                689 / IN_WIDTH: ping_storage_data_483 <= (fillup_transition == 1'b1) ? i_input_data[689 % IN_WIDTH] : ping_storage_data_483 ^ i_input_data[689 % IN_WIDTH];
                1076 / IN_WIDTH: ping_storage_data_483 <= (fillup_transition == 1'b1) ? i_input_data[1076 % IN_WIDTH] : ping_storage_data_483 ^ i_input_data[1076 % IN_WIDTH];
                default: ping_storage_data_483 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_483;
                endcase
            end else begin
                case (input_count)
                437 / IN_WIDTH: pong_storage_data_483 <= (fillup_transition == 1'b1) ? i_input_data[437 % IN_WIDTH] : pong_storage_data_483 ^ i_input_data[437 % IN_WIDTH];
                539 / IN_WIDTH: pong_storage_data_483 <= (fillup_transition == 1'b1) ? i_input_data[539 % IN_WIDTH] : pong_storage_data_483 ^ i_input_data[539 % IN_WIDTH];
                689 / IN_WIDTH: pong_storage_data_483 <= (fillup_transition == 1'b1) ? i_input_data[689 % IN_WIDTH] : pong_storage_data_483 ^ i_input_data[689 % IN_WIDTH];
                1076 / IN_WIDTH: pong_storage_data_483 <= (fillup_transition == 1'b1) ? i_input_data[1076 % IN_WIDTH] : pong_storage_data_483 ^ i_input_data[1076 % IN_WIDTH];
                default: pong_storage_data_483 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_483;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_483 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_483;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_483 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_483;
            end
        end
    end
end

logic ping_storage_data_484;
logic pong_storage_data_484;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_484 <= 1'b0;
        pong_storage_data_484 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                438 / IN_WIDTH: ping_storage_data_484 <= (fillup_transition == 1'b1) ? i_input_data[438 % IN_WIDTH] : ping_storage_data_484 ^ i_input_data[438 % IN_WIDTH];
                540 / IN_WIDTH: ping_storage_data_484 <= (fillup_transition == 1'b1) ? i_input_data[540 % IN_WIDTH] : ping_storage_data_484 ^ i_input_data[540 % IN_WIDTH];
                690 / IN_WIDTH: ping_storage_data_484 <= (fillup_transition == 1'b1) ? i_input_data[690 % IN_WIDTH] : ping_storage_data_484 ^ i_input_data[690 % IN_WIDTH];
                1077 / IN_WIDTH: ping_storage_data_484 <= (fillup_transition == 1'b1) ? i_input_data[1077 % IN_WIDTH] : ping_storage_data_484 ^ i_input_data[1077 % IN_WIDTH];
                default: ping_storage_data_484 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_484;
                endcase
            end else begin
                case (input_count)
                438 / IN_WIDTH: pong_storage_data_484 <= (fillup_transition == 1'b1) ? i_input_data[438 % IN_WIDTH] : pong_storage_data_484 ^ i_input_data[438 % IN_WIDTH];
                540 / IN_WIDTH: pong_storage_data_484 <= (fillup_transition == 1'b1) ? i_input_data[540 % IN_WIDTH] : pong_storage_data_484 ^ i_input_data[540 % IN_WIDTH];
                690 / IN_WIDTH: pong_storage_data_484 <= (fillup_transition == 1'b1) ? i_input_data[690 % IN_WIDTH] : pong_storage_data_484 ^ i_input_data[690 % IN_WIDTH];
                1077 / IN_WIDTH: pong_storage_data_484 <= (fillup_transition == 1'b1) ? i_input_data[1077 % IN_WIDTH] : pong_storage_data_484 ^ i_input_data[1077 % IN_WIDTH];
                default: pong_storage_data_484 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_484;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_484 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_484;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_484 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_484;
            end
        end
    end
end

logic ping_storage_data_485;
logic pong_storage_data_485;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_485 <= 1'b0;
        pong_storage_data_485 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                439 / IN_WIDTH: ping_storage_data_485 <= (fillup_transition == 1'b1) ? i_input_data[439 % IN_WIDTH] : ping_storage_data_485 ^ i_input_data[439 % IN_WIDTH];
                541 / IN_WIDTH: ping_storage_data_485 <= (fillup_transition == 1'b1) ? i_input_data[541 % IN_WIDTH] : ping_storage_data_485 ^ i_input_data[541 % IN_WIDTH];
                691 / IN_WIDTH: ping_storage_data_485 <= (fillup_transition == 1'b1) ? i_input_data[691 % IN_WIDTH] : ping_storage_data_485 ^ i_input_data[691 % IN_WIDTH];
                1078 / IN_WIDTH: ping_storage_data_485 <= (fillup_transition == 1'b1) ? i_input_data[1078 % IN_WIDTH] : ping_storage_data_485 ^ i_input_data[1078 % IN_WIDTH];
                default: ping_storage_data_485 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_485;
                endcase
            end else begin
                case (input_count)
                439 / IN_WIDTH: pong_storage_data_485 <= (fillup_transition == 1'b1) ? i_input_data[439 % IN_WIDTH] : pong_storage_data_485 ^ i_input_data[439 % IN_WIDTH];
                541 / IN_WIDTH: pong_storage_data_485 <= (fillup_transition == 1'b1) ? i_input_data[541 % IN_WIDTH] : pong_storage_data_485 ^ i_input_data[541 % IN_WIDTH];
                691 / IN_WIDTH: pong_storage_data_485 <= (fillup_transition == 1'b1) ? i_input_data[691 % IN_WIDTH] : pong_storage_data_485 ^ i_input_data[691 % IN_WIDTH];
                1078 / IN_WIDTH: pong_storage_data_485 <= (fillup_transition == 1'b1) ? i_input_data[1078 % IN_WIDTH] : pong_storage_data_485 ^ i_input_data[1078 % IN_WIDTH];
                default: pong_storage_data_485 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_485;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_485 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_485;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_485 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_485;
            end
        end
    end
end

logic ping_storage_data_486;
logic pong_storage_data_486;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_486 <= 1'b0;
        pong_storage_data_486 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                440 / IN_WIDTH: ping_storage_data_486 <= (fillup_transition == 1'b1) ? i_input_data[440 % IN_WIDTH] : ping_storage_data_486 ^ i_input_data[440 % IN_WIDTH];
                542 / IN_WIDTH: ping_storage_data_486 <= (fillup_transition == 1'b1) ? i_input_data[542 % IN_WIDTH] : ping_storage_data_486 ^ i_input_data[542 % IN_WIDTH];
                692 / IN_WIDTH: ping_storage_data_486 <= (fillup_transition == 1'b1) ? i_input_data[692 % IN_WIDTH] : ping_storage_data_486 ^ i_input_data[692 % IN_WIDTH];
                1079 / IN_WIDTH: ping_storage_data_486 <= (fillup_transition == 1'b1) ? i_input_data[1079 % IN_WIDTH] : ping_storage_data_486 ^ i_input_data[1079 % IN_WIDTH];
                default: ping_storage_data_486 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_486;
                endcase
            end else begin
                case (input_count)
                440 / IN_WIDTH: pong_storage_data_486 <= (fillup_transition == 1'b1) ? i_input_data[440 % IN_WIDTH] : pong_storage_data_486 ^ i_input_data[440 % IN_WIDTH];
                542 / IN_WIDTH: pong_storage_data_486 <= (fillup_transition == 1'b1) ? i_input_data[542 % IN_WIDTH] : pong_storage_data_486 ^ i_input_data[542 % IN_WIDTH];
                692 / IN_WIDTH: pong_storage_data_486 <= (fillup_transition == 1'b1) ? i_input_data[692 % IN_WIDTH] : pong_storage_data_486 ^ i_input_data[692 % IN_WIDTH];
                1079 / IN_WIDTH: pong_storage_data_486 <= (fillup_transition == 1'b1) ? i_input_data[1079 % IN_WIDTH] : pong_storage_data_486 ^ i_input_data[1079 % IN_WIDTH];
                default: pong_storage_data_486 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_486;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_486 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_486;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_486 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_486;
            end
        end
    end
end

logic ping_storage_data_487;
logic pong_storage_data_487;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_487 <= 1'b0;
        pong_storage_data_487 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                441 / IN_WIDTH: ping_storage_data_487 <= (fillup_transition == 1'b1) ? i_input_data[441 % IN_WIDTH] : ping_storage_data_487 ^ i_input_data[441 % IN_WIDTH];
                543 / IN_WIDTH: ping_storage_data_487 <= (fillup_transition == 1'b1) ? i_input_data[543 % IN_WIDTH] : ping_storage_data_487 ^ i_input_data[543 % IN_WIDTH];
                693 / IN_WIDTH: ping_storage_data_487 <= (fillup_transition == 1'b1) ? i_input_data[693 % IN_WIDTH] : ping_storage_data_487 ^ i_input_data[693 % IN_WIDTH];
                1080 / IN_WIDTH: ping_storage_data_487 <= (fillup_transition == 1'b1) ? i_input_data[1080 % IN_WIDTH] : ping_storage_data_487 ^ i_input_data[1080 % IN_WIDTH];
                default: ping_storage_data_487 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_487;
                endcase
            end else begin
                case (input_count)
                441 / IN_WIDTH: pong_storage_data_487 <= (fillup_transition == 1'b1) ? i_input_data[441 % IN_WIDTH] : pong_storage_data_487 ^ i_input_data[441 % IN_WIDTH];
                543 / IN_WIDTH: pong_storage_data_487 <= (fillup_transition == 1'b1) ? i_input_data[543 % IN_WIDTH] : pong_storage_data_487 ^ i_input_data[543 % IN_WIDTH];
                693 / IN_WIDTH: pong_storage_data_487 <= (fillup_transition == 1'b1) ? i_input_data[693 % IN_WIDTH] : pong_storage_data_487 ^ i_input_data[693 % IN_WIDTH];
                1080 / IN_WIDTH: pong_storage_data_487 <= (fillup_transition == 1'b1) ? i_input_data[1080 % IN_WIDTH] : pong_storage_data_487 ^ i_input_data[1080 % IN_WIDTH];
                default: pong_storage_data_487 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_487;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_487 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_487;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_487 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_487;
            end
        end
    end
end

logic ping_storage_data_488;
logic pong_storage_data_488;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_488 <= 1'b0;
        pong_storage_data_488 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                442 / IN_WIDTH: ping_storage_data_488 <= (fillup_transition == 1'b1) ? i_input_data[442 % IN_WIDTH] : ping_storage_data_488 ^ i_input_data[442 % IN_WIDTH];
                544 / IN_WIDTH: ping_storage_data_488 <= (fillup_transition == 1'b1) ? i_input_data[544 % IN_WIDTH] : ping_storage_data_488 ^ i_input_data[544 % IN_WIDTH];
                694 / IN_WIDTH: ping_storage_data_488 <= (fillup_transition == 1'b1) ? i_input_data[694 % IN_WIDTH] : ping_storage_data_488 ^ i_input_data[694 % IN_WIDTH];
                1081 / IN_WIDTH: ping_storage_data_488 <= (fillup_transition == 1'b1) ? i_input_data[1081 % IN_WIDTH] : ping_storage_data_488 ^ i_input_data[1081 % IN_WIDTH];
                default: ping_storage_data_488 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_488;
                endcase
            end else begin
                case (input_count)
                442 / IN_WIDTH: pong_storage_data_488 <= (fillup_transition == 1'b1) ? i_input_data[442 % IN_WIDTH] : pong_storage_data_488 ^ i_input_data[442 % IN_WIDTH];
                544 / IN_WIDTH: pong_storage_data_488 <= (fillup_transition == 1'b1) ? i_input_data[544 % IN_WIDTH] : pong_storage_data_488 ^ i_input_data[544 % IN_WIDTH];
                694 / IN_WIDTH: pong_storage_data_488 <= (fillup_transition == 1'b1) ? i_input_data[694 % IN_WIDTH] : pong_storage_data_488 ^ i_input_data[694 % IN_WIDTH];
                1081 / IN_WIDTH: pong_storage_data_488 <= (fillup_transition == 1'b1) ? i_input_data[1081 % IN_WIDTH] : pong_storage_data_488 ^ i_input_data[1081 % IN_WIDTH];
                default: pong_storage_data_488 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_488;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_488 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_488;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_488 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_488;
            end
        end
    end
end

logic ping_storage_data_489;
logic pong_storage_data_489;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_489 <= 1'b0;
        pong_storage_data_489 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                443 / IN_WIDTH: ping_storage_data_489 <= (fillup_transition == 1'b1) ? i_input_data[443 % IN_WIDTH] : ping_storage_data_489 ^ i_input_data[443 % IN_WIDTH];
                545 / IN_WIDTH: ping_storage_data_489 <= (fillup_transition == 1'b1) ? i_input_data[545 % IN_WIDTH] : ping_storage_data_489 ^ i_input_data[545 % IN_WIDTH];
                695 / IN_WIDTH: ping_storage_data_489 <= (fillup_transition == 1'b1) ? i_input_data[695 % IN_WIDTH] : ping_storage_data_489 ^ i_input_data[695 % IN_WIDTH];
                1082 / IN_WIDTH: ping_storage_data_489 <= (fillup_transition == 1'b1) ? i_input_data[1082 % IN_WIDTH] : ping_storage_data_489 ^ i_input_data[1082 % IN_WIDTH];
                default: ping_storage_data_489 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_489;
                endcase
            end else begin
                case (input_count)
                443 / IN_WIDTH: pong_storage_data_489 <= (fillup_transition == 1'b1) ? i_input_data[443 % IN_WIDTH] : pong_storage_data_489 ^ i_input_data[443 % IN_WIDTH];
                545 / IN_WIDTH: pong_storage_data_489 <= (fillup_transition == 1'b1) ? i_input_data[545 % IN_WIDTH] : pong_storage_data_489 ^ i_input_data[545 % IN_WIDTH];
                695 / IN_WIDTH: pong_storage_data_489 <= (fillup_transition == 1'b1) ? i_input_data[695 % IN_WIDTH] : pong_storage_data_489 ^ i_input_data[695 % IN_WIDTH];
                1082 / IN_WIDTH: pong_storage_data_489 <= (fillup_transition == 1'b1) ? i_input_data[1082 % IN_WIDTH] : pong_storage_data_489 ^ i_input_data[1082 % IN_WIDTH];
                default: pong_storage_data_489 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_489;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_489 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_489;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_489 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_489;
            end
        end
    end
end

logic ping_storage_data_490;
logic pong_storage_data_490;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_490 <= 1'b0;
        pong_storage_data_490 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                444 / IN_WIDTH: ping_storage_data_490 <= (fillup_transition == 1'b1) ? i_input_data[444 % IN_WIDTH] : ping_storage_data_490 ^ i_input_data[444 % IN_WIDTH];
                546 / IN_WIDTH: ping_storage_data_490 <= (fillup_transition == 1'b1) ? i_input_data[546 % IN_WIDTH] : ping_storage_data_490 ^ i_input_data[546 % IN_WIDTH];
                696 / IN_WIDTH: ping_storage_data_490 <= (fillup_transition == 1'b1) ? i_input_data[696 % IN_WIDTH] : ping_storage_data_490 ^ i_input_data[696 % IN_WIDTH];
                1083 / IN_WIDTH: ping_storage_data_490 <= (fillup_transition == 1'b1) ? i_input_data[1083 % IN_WIDTH] : ping_storage_data_490 ^ i_input_data[1083 % IN_WIDTH];
                default: ping_storage_data_490 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_490;
                endcase
            end else begin
                case (input_count)
                444 / IN_WIDTH: pong_storage_data_490 <= (fillup_transition == 1'b1) ? i_input_data[444 % IN_WIDTH] : pong_storage_data_490 ^ i_input_data[444 % IN_WIDTH];
                546 / IN_WIDTH: pong_storage_data_490 <= (fillup_transition == 1'b1) ? i_input_data[546 % IN_WIDTH] : pong_storage_data_490 ^ i_input_data[546 % IN_WIDTH];
                696 / IN_WIDTH: pong_storage_data_490 <= (fillup_transition == 1'b1) ? i_input_data[696 % IN_WIDTH] : pong_storage_data_490 ^ i_input_data[696 % IN_WIDTH];
                1083 / IN_WIDTH: pong_storage_data_490 <= (fillup_transition == 1'b1) ? i_input_data[1083 % IN_WIDTH] : pong_storage_data_490 ^ i_input_data[1083 % IN_WIDTH];
                default: pong_storage_data_490 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_490;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_490 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_490;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_490 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_490;
            end
        end
    end
end

logic ping_storage_data_491;
logic pong_storage_data_491;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_491 <= 1'b0;
        pong_storage_data_491 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                445 / IN_WIDTH: ping_storage_data_491 <= (fillup_transition == 1'b1) ? i_input_data[445 % IN_WIDTH] : ping_storage_data_491 ^ i_input_data[445 % IN_WIDTH];
                547 / IN_WIDTH: ping_storage_data_491 <= (fillup_transition == 1'b1) ? i_input_data[547 % IN_WIDTH] : ping_storage_data_491 ^ i_input_data[547 % IN_WIDTH];
                697 / IN_WIDTH: ping_storage_data_491 <= (fillup_transition == 1'b1) ? i_input_data[697 % IN_WIDTH] : ping_storage_data_491 ^ i_input_data[697 % IN_WIDTH];
                1084 / IN_WIDTH: ping_storage_data_491 <= (fillup_transition == 1'b1) ? i_input_data[1084 % IN_WIDTH] : ping_storage_data_491 ^ i_input_data[1084 % IN_WIDTH];
                default: ping_storage_data_491 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_491;
                endcase
            end else begin
                case (input_count)
                445 / IN_WIDTH: pong_storage_data_491 <= (fillup_transition == 1'b1) ? i_input_data[445 % IN_WIDTH] : pong_storage_data_491 ^ i_input_data[445 % IN_WIDTH];
                547 / IN_WIDTH: pong_storage_data_491 <= (fillup_transition == 1'b1) ? i_input_data[547 % IN_WIDTH] : pong_storage_data_491 ^ i_input_data[547 % IN_WIDTH];
                697 / IN_WIDTH: pong_storage_data_491 <= (fillup_transition == 1'b1) ? i_input_data[697 % IN_WIDTH] : pong_storage_data_491 ^ i_input_data[697 % IN_WIDTH];
                1084 / IN_WIDTH: pong_storage_data_491 <= (fillup_transition == 1'b1) ? i_input_data[1084 % IN_WIDTH] : pong_storage_data_491 ^ i_input_data[1084 % IN_WIDTH];
                default: pong_storage_data_491 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_491;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_491 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_491;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_491 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_491;
            end
        end
    end
end

logic ping_storage_data_492;
logic pong_storage_data_492;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_492 <= 1'b0;
        pong_storage_data_492 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                446 / IN_WIDTH: ping_storage_data_492 <= (fillup_transition == 1'b1) ? i_input_data[446 % IN_WIDTH] : ping_storage_data_492 ^ i_input_data[446 % IN_WIDTH];
                548 / IN_WIDTH: ping_storage_data_492 <= (fillup_transition == 1'b1) ? i_input_data[548 % IN_WIDTH] : ping_storage_data_492 ^ i_input_data[548 % IN_WIDTH];
                698 / IN_WIDTH: ping_storage_data_492 <= (fillup_transition == 1'b1) ? i_input_data[698 % IN_WIDTH] : ping_storage_data_492 ^ i_input_data[698 % IN_WIDTH];
                1085 / IN_WIDTH: ping_storage_data_492 <= (fillup_transition == 1'b1) ? i_input_data[1085 % IN_WIDTH] : ping_storage_data_492 ^ i_input_data[1085 % IN_WIDTH];
                default: ping_storage_data_492 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_492;
                endcase
            end else begin
                case (input_count)
                446 / IN_WIDTH: pong_storage_data_492 <= (fillup_transition == 1'b1) ? i_input_data[446 % IN_WIDTH] : pong_storage_data_492 ^ i_input_data[446 % IN_WIDTH];
                548 / IN_WIDTH: pong_storage_data_492 <= (fillup_transition == 1'b1) ? i_input_data[548 % IN_WIDTH] : pong_storage_data_492 ^ i_input_data[548 % IN_WIDTH];
                698 / IN_WIDTH: pong_storage_data_492 <= (fillup_transition == 1'b1) ? i_input_data[698 % IN_WIDTH] : pong_storage_data_492 ^ i_input_data[698 % IN_WIDTH];
                1085 / IN_WIDTH: pong_storage_data_492 <= (fillup_transition == 1'b1) ? i_input_data[1085 % IN_WIDTH] : pong_storage_data_492 ^ i_input_data[1085 % IN_WIDTH];
                default: pong_storage_data_492 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_492;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_492 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_492;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_492 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_492;
            end
        end
    end
end

logic ping_storage_data_493;
logic pong_storage_data_493;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_493 <= 1'b0;
        pong_storage_data_493 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                447 / IN_WIDTH: ping_storage_data_493 <= (fillup_transition == 1'b1) ? i_input_data[447 % IN_WIDTH] : ping_storage_data_493 ^ i_input_data[447 % IN_WIDTH];
                549 / IN_WIDTH: ping_storage_data_493 <= (fillup_transition == 1'b1) ? i_input_data[549 % IN_WIDTH] : ping_storage_data_493 ^ i_input_data[549 % IN_WIDTH];
                699 / IN_WIDTH: ping_storage_data_493 <= (fillup_transition == 1'b1) ? i_input_data[699 % IN_WIDTH] : ping_storage_data_493 ^ i_input_data[699 % IN_WIDTH];
                1086 / IN_WIDTH: ping_storage_data_493 <= (fillup_transition == 1'b1) ? i_input_data[1086 % IN_WIDTH] : ping_storage_data_493 ^ i_input_data[1086 % IN_WIDTH];
                default: ping_storage_data_493 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_493;
                endcase
            end else begin
                case (input_count)
                447 / IN_WIDTH: pong_storage_data_493 <= (fillup_transition == 1'b1) ? i_input_data[447 % IN_WIDTH] : pong_storage_data_493 ^ i_input_data[447 % IN_WIDTH];
                549 / IN_WIDTH: pong_storage_data_493 <= (fillup_transition == 1'b1) ? i_input_data[549 % IN_WIDTH] : pong_storage_data_493 ^ i_input_data[549 % IN_WIDTH];
                699 / IN_WIDTH: pong_storage_data_493 <= (fillup_transition == 1'b1) ? i_input_data[699 % IN_WIDTH] : pong_storage_data_493 ^ i_input_data[699 % IN_WIDTH];
                1086 / IN_WIDTH: pong_storage_data_493 <= (fillup_transition == 1'b1) ? i_input_data[1086 % IN_WIDTH] : pong_storage_data_493 ^ i_input_data[1086 % IN_WIDTH];
                default: pong_storage_data_493 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_493;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_493 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_493;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_493 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_493;
            end
        end
    end
end

logic ping_storage_data_494;
logic pong_storage_data_494;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_494 <= 1'b0;
        pong_storage_data_494 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                448 / IN_WIDTH: ping_storage_data_494 <= (fillup_transition == 1'b1) ? i_input_data[448 % IN_WIDTH] : ping_storage_data_494 ^ i_input_data[448 % IN_WIDTH];
                550 / IN_WIDTH: ping_storage_data_494 <= (fillup_transition == 1'b1) ? i_input_data[550 % IN_WIDTH] : ping_storage_data_494 ^ i_input_data[550 % IN_WIDTH];
                700 / IN_WIDTH: ping_storage_data_494 <= (fillup_transition == 1'b1) ? i_input_data[700 % IN_WIDTH] : ping_storage_data_494 ^ i_input_data[700 % IN_WIDTH];
                1087 / IN_WIDTH: ping_storage_data_494 <= (fillup_transition == 1'b1) ? i_input_data[1087 % IN_WIDTH] : ping_storage_data_494 ^ i_input_data[1087 % IN_WIDTH];
                default: ping_storage_data_494 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_494;
                endcase
            end else begin
                case (input_count)
                448 / IN_WIDTH: pong_storage_data_494 <= (fillup_transition == 1'b1) ? i_input_data[448 % IN_WIDTH] : pong_storage_data_494 ^ i_input_data[448 % IN_WIDTH];
                550 / IN_WIDTH: pong_storage_data_494 <= (fillup_transition == 1'b1) ? i_input_data[550 % IN_WIDTH] : pong_storage_data_494 ^ i_input_data[550 % IN_WIDTH];
                700 / IN_WIDTH: pong_storage_data_494 <= (fillup_transition == 1'b1) ? i_input_data[700 % IN_WIDTH] : pong_storage_data_494 ^ i_input_data[700 % IN_WIDTH];
                1087 / IN_WIDTH: pong_storage_data_494 <= (fillup_transition == 1'b1) ? i_input_data[1087 % IN_WIDTH] : pong_storage_data_494 ^ i_input_data[1087 % IN_WIDTH];
                default: pong_storage_data_494 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_494;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_494 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_494;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_494 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_494;
            end
        end
    end
end

logic ping_storage_data_495;
logic pong_storage_data_495;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_495 <= 1'b0;
        pong_storage_data_495 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                449 / IN_WIDTH: ping_storage_data_495 <= (fillup_transition == 1'b1) ? i_input_data[449 % IN_WIDTH] : ping_storage_data_495 ^ i_input_data[449 % IN_WIDTH];
                551 / IN_WIDTH: ping_storage_data_495 <= (fillup_transition == 1'b1) ? i_input_data[551 % IN_WIDTH] : ping_storage_data_495 ^ i_input_data[551 % IN_WIDTH];
                701 / IN_WIDTH: ping_storage_data_495 <= (fillup_transition == 1'b1) ? i_input_data[701 % IN_WIDTH] : ping_storage_data_495 ^ i_input_data[701 % IN_WIDTH];
                1088 / IN_WIDTH: ping_storage_data_495 <= (fillup_transition == 1'b1) ? i_input_data[1088 % IN_WIDTH] : ping_storage_data_495 ^ i_input_data[1088 % IN_WIDTH];
                default: ping_storage_data_495 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_495;
                endcase
            end else begin
                case (input_count)
                449 / IN_WIDTH: pong_storage_data_495 <= (fillup_transition == 1'b1) ? i_input_data[449 % IN_WIDTH] : pong_storage_data_495 ^ i_input_data[449 % IN_WIDTH];
                551 / IN_WIDTH: pong_storage_data_495 <= (fillup_transition == 1'b1) ? i_input_data[551 % IN_WIDTH] : pong_storage_data_495 ^ i_input_data[551 % IN_WIDTH];
                701 / IN_WIDTH: pong_storage_data_495 <= (fillup_transition == 1'b1) ? i_input_data[701 % IN_WIDTH] : pong_storage_data_495 ^ i_input_data[701 % IN_WIDTH];
                1088 / IN_WIDTH: pong_storage_data_495 <= (fillup_transition == 1'b1) ? i_input_data[1088 % IN_WIDTH] : pong_storage_data_495 ^ i_input_data[1088 % IN_WIDTH];
                default: pong_storage_data_495 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_495;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_495 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_495;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_495 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_495;
            end
        end
    end
end

logic ping_storage_data_496;
logic pong_storage_data_496;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_496 <= 1'b0;
        pong_storage_data_496 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                450 / IN_WIDTH: ping_storage_data_496 <= (fillup_transition == 1'b1) ? i_input_data[450 % IN_WIDTH] : ping_storage_data_496 ^ i_input_data[450 % IN_WIDTH];
                552 / IN_WIDTH: ping_storage_data_496 <= (fillup_transition == 1'b1) ? i_input_data[552 % IN_WIDTH] : ping_storage_data_496 ^ i_input_data[552 % IN_WIDTH];
                702 / IN_WIDTH: ping_storage_data_496 <= (fillup_transition == 1'b1) ? i_input_data[702 % IN_WIDTH] : ping_storage_data_496 ^ i_input_data[702 % IN_WIDTH];
                1089 / IN_WIDTH: ping_storage_data_496 <= (fillup_transition == 1'b1) ? i_input_data[1089 % IN_WIDTH] : ping_storage_data_496 ^ i_input_data[1089 % IN_WIDTH];
                default: ping_storage_data_496 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_496;
                endcase
            end else begin
                case (input_count)
                450 / IN_WIDTH: pong_storage_data_496 <= (fillup_transition == 1'b1) ? i_input_data[450 % IN_WIDTH] : pong_storage_data_496 ^ i_input_data[450 % IN_WIDTH];
                552 / IN_WIDTH: pong_storage_data_496 <= (fillup_transition == 1'b1) ? i_input_data[552 % IN_WIDTH] : pong_storage_data_496 ^ i_input_data[552 % IN_WIDTH];
                702 / IN_WIDTH: pong_storage_data_496 <= (fillup_transition == 1'b1) ? i_input_data[702 % IN_WIDTH] : pong_storage_data_496 ^ i_input_data[702 % IN_WIDTH];
                1089 / IN_WIDTH: pong_storage_data_496 <= (fillup_transition == 1'b1) ? i_input_data[1089 % IN_WIDTH] : pong_storage_data_496 ^ i_input_data[1089 % IN_WIDTH];
                default: pong_storage_data_496 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_496;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_496 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_496;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_496 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_496;
            end
        end
    end
end

logic ping_storage_data_497;
logic pong_storage_data_497;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_497 <= 1'b0;
        pong_storage_data_497 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                451 / IN_WIDTH: ping_storage_data_497 <= (fillup_transition == 1'b1) ? i_input_data[451 % IN_WIDTH] : ping_storage_data_497 ^ i_input_data[451 % IN_WIDTH];
                553 / IN_WIDTH: ping_storage_data_497 <= (fillup_transition == 1'b1) ? i_input_data[553 % IN_WIDTH] : ping_storage_data_497 ^ i_input_data[553 % IN_WIDTH];
                703 / IN_WIDTH: ping_storage_data_497 <= (fillup_transition == 1'b1) ? i_input_data[703 % IN_WIDTH] : ping_storage_data_497 ^ i_input_data[703 % IN_WIDTH];
                1090 / IN_WIDTH: ping_storage_data_497 <= (fillup_transition == 1'b1) ? i_input_data[1090 % IN_WIDTH] : ping_storage_data_497 ^ i_input_data[1090 % IN_WIDTH];
                default: ping_storage_data_497 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_497;
                endcase
            end else begin
                case (input_count)
                451 / IN_WIDTH: pong_storage_data_497 <= (fillup_transition == 1'b1) ? i_input_data[451 % IN_WIDTH] : pong_storage_data_497 ^ i_input_data[451 % IN_WIDTH];
                553 / IN_WIDTH: pong_storage_data_497 <= (fillup_transition == 1'b1) ? i_input_data[553 % IN_WIDTH] : pong_storage_data_497 ^ i_input_data[553 % IN_WIDTH];
                703 / IN_WIDTH: pong_storage_data_497 <= (fillup_transition == 1'b1) ? i_input_data[703 % IN_WIDTH] : pong_storage_data_497 ^ i_input_data[703 % IN_WIDTH];
                1090 / IN_WIDTH: pong_storage_data_497 <= (fillup_transition == 1'b1) ? i_input_data[1090 % IN_WIDTH] : pong_storage_data_497 ^ i_input_data[1090 % IN_WIDTH];
                default: pong_storage_data_497 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_497;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_497 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_497;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_497 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_497;
            end
        end
    end
end

logic ping_storage_data_498;
logic pong_storage_data_498;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_498 <= 1'b0;
        pong_storage_data_498 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                452 / IN_WIDTH: ping_storage_data_498 <= (fillup_transition == 1'b1) ? i_input_data[452 % IN_WIDTH] : ping_storage_data_498 ^ i_input_data[452 % IN_WIDTH];
                554 / IN_WIDTH: ping_storage_data_498 <= (fillup_transition == 1'b1) ? i_input_data[554 % IN_WIDTH] : ping_storage_data_498 ^ i_input_data[554 % IN_WIDTH];
                704 / IN_WIDTH: ping_storage_data_498 <= (fillup_transition == 1'b1) ? i_input_data[704 % IN_WIDTH] : ping_storage_data_498 ^ i_input_data[704 % IN_WIDTH];
                1091 / IN_WIDTH: ping_storage_data_498 <= (fillup_transition == 1'b1) ? i_input_data[1091 % IN_WIDTH] : ping_storage_data_498 ^ i_input_data[1091 % IN_WIDTH];
                default: ping_storage_data_498 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_498;
                endcase
            end else begin
                case (input_count)
                452 / IN_WIDTH: pong_storage_data_498 <= (fillup_transition == 1'b1) ? i_input_data[452 % IN_WIDTH] : pong_storage_data_498 ^ i_input_data[452 % IN_WIDTH];
                554 / IN_WIDTH: pong_storage_data_498 <= (fillup_transition == 1'b1) ? i_input_data[554 % IN_WIDTH] : pong_storage_data_498 ^ i_input_data[554 % IN_WIDTH];
                704 / IN_WIDTH: pong_storage_data_498 <= (fillup_transition == 1'b1) ? i_input_data[704 % IN_WIDTH] : pong_storage_data_498 ^ i_input_data[704 % IN_WIDTH];
                1091 / IN_WIDTH: pong_storage_data_498 <= (fillup_transition == 1'b1) ? i_input_data[1091 % IN_WIDTH] : pong_storage_data_498 ^ i_input_data[1091 % IN_WIDTH];
                default: pong_storage_data_498 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_498;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_498 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_498;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_498 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_498;
            end
        end
    end
end

logic ping_storage_data_499;
logic pong_storage_data_499;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_499 <= 1'b0;
        pong_storage_data_499 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                453 / IN_WIDTH: ping_storage_data_499 <= (fillup_transition == 1'b1) ? i_input_data[453 % IN_WIDTH] : ping_storage_data_499 ^ i_input_data[453 % IN_WIDTH];
                555 / IN_WIDTH: ping_storage_data_499 <= (fillup_transition == 1'b1) ? i_input_data[555 % IN_WIDTH] : ping_storage_data_499 ^ i_input_data[555 % IN_WIDTH];
                705 / IN_WIDTH: ping_storage_data_499 <= (fillup_transition == 1'b1) ? i_input_data[705 % IN_WIDTH] : ping_storage_data_499 ^ i_input_data[705 % IN_WIDTH];
                1092 / IN_WIDTH: ping_storage_data_499 <= (fillup_transition == 1'b1) ? i_input_data[1092 % IN_WIDTH] : ping_storage_data_499 ^ i_input_data[1092 % IN_WIDTH];
                default: ping_storage_data_499 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_499;
                endcase
            end else begin
                case (input_count)
                453 / IN_WIDTH: pong_storage_data_499 <= (fillup_transition == 1'b1) ? i_input_data[453 % IN_WIDTH] : pong_storage_data_499 ^ i_input_data[453 % IN_WIDTH];
                555 / IN_WIDTH: pong_storage_data_499 <= (fillup_transition == 1'b1) ? i_input_data[555 % IN_WIDTH] : pong_storage_data_499 ^ i_input_data[555 % IN_WIDTH];
                705 / IN_WIDTH: pong_storage_data_499 <= (fillup_transition == 1'b1) ? i_input_data[705 % IN_WIDTH] : pong_storage_data_499 ^ i_input_data[705 % IN_WIDTH];
                1092 / IN_WIDTH: pong_storage_data_499 <= (fillup_transition == 1'b1) ? i_input_data[1092 % IN_WIDTH] : pong_storage_data_499 ^ i_input_data[1092 % IN_WIDTH];
                default: pong_storage_data_499 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_499;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_499 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_499;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_499 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_499;
            end
        end
    end
end

logic ping_storage_data_500;
logic pong_storage_data_500;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_500 <= 1'b0;
        pong_storage_data_500 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                454 / IN_WIDTH: ping_storage_data_500 <= (fillup_transition == 1'b1) ? i_input_data[454 % IN_WIDTH] : ping_storage_data_500 ^ i_input_data[454 % IN_WIDTH];
                556 / IN_WIDTH: ping_storage_data_500 <= (fillup_transition == 1'b1) ? i_input_data[556 % IN_WIDTH] : ping_storage_data_500 ^ i_input_data[556 % IN_WIDTH];
                706 / IN_WIDTH: ping_storage_data_500 <= (fillup_transition == 1'b1) ? i_input_data[706 % IN_WIDTH] : ping_storage_data_500 ^ i_input_data[706 % IN_WIDTH];
                1093 / IN_WIDTH: ping_storage_data_500 <= (fillup_transition == 1'b1) ? i_input_data[1093 % IN_WIDTH] : ping_storage_data_500 ^ i_input_data[1093 % IN_WIDTH];
                default: ping_storage_data_500 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_500;
                endcase
            end else begin
                case (input_count)
                454 / IN_WIDTH: pong_storage_data_500 <= (fillup_transition == 1'b1) ? i_input_data[454 % IN_WIDTH] : pong_storage_data_500 ^ i_input_data[454 % IN_WIDTH];
                556 / IN_WIDTH: pong_storage_data_500 <= (fillup_transition == 1'b1) ? i_input_data[556 % IN_WIDTH] : pong_storage_data_500 ^ i_input_data[556 % IN_WIDTH];
                706 / IN_WIDTH: pong_storage_data_500 <= (fillup_transition == 1'b1) ? i_input_data[706 % IN_WIDTH] : pong_storage_data_500 ^ i_input_data[706 % IN_WIDTH];
                1093 / IN_WIDTH: pong_storage_data_500 <= (fillup_transition == 1'b1) ? i_input_data[1093 % IN_WIDTH] : pong_storage_data_500 ^ i_input_data[1093 % IN_WIDTH];
                default: pong_storage_data_500 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_500;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_500 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_500;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_500 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_500;
            end
        end
    end
end

logic ping_storage_data_501;
logic pong_storage_data_501;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_501 <= 1'b0;
        pong_storage_data_501 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                455 / IN_WIDTH: ping_storage_data_501 <= (fillup_transition == 1'b1) ? i_input_data[455 % IN_WIDTH] : ping_storage_data_501 ^ i_input_data[455 % IN_WIDTH];
                557 / IN_WIDTH: ping_storage_data_501 <= (fillup_transition == 1'b1) ? i_input_data[557 % IN_WIDTH] : ping_storage_data_501 ^ i_input_data[557 % IN_WIDTH];
                707 / IN_WIDTH: ping_storage_data_501 <= (fillup_transition == 1'b1) ? i_input_data[707 % IN_WIDTH] : ping_storage_data_501 ^ i_input_data[707 % IN_WIDTH];
                1094 / IN_WIDTH: ping_storage_data_501 <= (fillup_transition == 1'b1) ? i_input_data[1094 % IN_WIDTH] : ping_storage_data_501 ^ i_input_data[1094 % IN_WIDTH];
                default: ping_storage_data_501 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_501;
                endcase
            end else begin
                case (input_count)
                455 / IN_WIDTH: pong_storage_data_501 <= (fillup_transition == 1'b1) ? i_input_data[455 % IN_WIDTH] : pong_storage_data_501 ^ i_input_data[455 % IN_WIDTH];
                557 / IN_WIDTH: pong_storage_data_501 <= (fillup_transition == 1'b1) ? i_input_data[557 % IN_WIDTH] : pong_storage_data_501 ^ i_input_data[557 % IN_WIDTH];
                707 / IN_WIDTH: pong_storage_data_501 <= (fillup_transition == 1'b1) ? i_input_data[707 % IN_WIDTH] : pong_storage_data_501 ^ i_input_data[707 % IN_WIDTH];
                1094 / IN_WIDTH: pong_storage_data_501 <= (fillup_transition == 1'b1) ? i_input_data[1094 % IN_WIDTH] : pong_storage_data_501 ^ i_input_data[1094 % IN_WIDTH];
                default: pong_storage_data_501 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_501;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_501 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_501;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_501 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_501;
            end
        end
    end
end

logic ping_storage_data_502;
logic pong_storage_data_502;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_502 <= 1'b0;
        pong_storage_data_502 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                456 / IN_WIDTH: ping_storage_data_502 <= (fillup_transition == 1'b1) ? i_input_data[456 % IN_WIDTH] : ping_storage_data_502 ^ i_input_data[456 % IN_WIDTH];
                558 / IN_WIDTH: ping_storage_data_502 <= (fillup_transition == 1'b1) ? i_input_data[558 % IN_WIDTH] : ping_storage_data_502 ^ i_input_data[558 % IN_WIDTH];
                708 / IN_WIDTH: ping_storage_data_502 <= (fillup_transition == 1'b1) ? i_input_data[708 % IN_WIDTH] : ping_storage_data_502 ^ i_input_data[708 % IN_WIDTH];
                1095 / IN_WIDTH: ping_storage_data_502 <= (fillup_transition == 1'b1) ? i_input_data[1095 % IN_WIDTH] : ping_storage_data_502 ^ i_input_data[1095 % IN_WIDTH];
                default: ping_storage_data_502 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_502;
                endcase
            end else begin
                case (input_count)
                456 / IN_WIDTH: pong_storage_data_502 <= (fillup_transition == 1'b1) ? i_input_data[456 % IN_WIDTH] : pong_storage_data_502 ^ i_input_data[456 % IN_WIDTH];
                558 / IN_WIDTH: pong_storage_data_502 <= (fillup_transition == 1'b1) ? i_input_data[558 % IN_WIDTH] : pong_storage_data_502 ^ i_input_data[558 % IN_WIDTH];
                708 / IN_WIDTH: pong_storage_data_502 <= (fillup_transition == 1'b1) ? i_input_data[708 % IN_WIDTH] : pong_storage_data_502 ^ i_input_data[708 % IN_WIDTH];
                1095 / IN_WIDTH: pong_storage_data_502 <= (fillup_transition == 1'b1) ? i_input_data[1095 % IN_WIDTH] : pong_storage_data_502 ^ i_input_data[1095 % IN_WIDTH];
                default: pong_storage_data_502 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_502;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_502 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_502;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_502 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_502;
            end
        end
    end
end

logic ping_storage_data_503;
logic pong_storage_data_503;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_503 <= 1'b0;
        pong_storage_data_503 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                457 / IN_WIDTH: ping_storage_data_503 <= (fillup_transition == 1'b1) ? i_input_data[457 % IN_WIDTH] : ping_storage_data_503 ^ i_input_data[457 % IN_WIDTH];
                559 / IN_WIDTH: ping_storage_data_503 <= (fillup_transition == 1'b1) ? i_input_data[559 % IN_WIDTH] : ping_storage_data_503 ^ i_input_data[559 % IN_WIDTH];
                709 / IN_WIDTH: ping_storage_data_503 <= (fillup_transition == 1'b1) ? i_input_data[709 % IN_WIDTH] : ping_storage_data_503 ^ i_input_data[709 % IN_WIDTH];
                1096 / IN_WIDTH: ping_storage_data_503 <= (fillup_transition == 1'b1) ? i_input_data[1096 % IN_WIDTH] : ping_storage_data_503 ^ i_input_data[1096 % IN_WIDTH];
                default: ping_storage_data_503 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_503;
                endcase
            end else begin
                case (input_count)
                457 / IN_WIDTH: pong_storage_data_503 <= (fillup_transition == 1'b1) ? i_input_data[457 % IN_WIDTH] : pong_storage_data_503 ^ i_input_data[457 % IN_WIDTH];
                559 / IN_WIDTH: pong_storage_data_503 <= (fillup_transition == 1'b1) ? i_input_data[559 % IN_WIDTH] : pong_storage_data_503 ^ i_input_data[559 % IN_WIDTH];
                709 / IN_WIDTH: pong_storage_data_503 <= (fillup_transition == 1'b1) ? i_input_data[709 % IN_WIDTH] : pong_storage_data_503 ^ i_input_data[709 % IN_WIDTH];
                1096 / IN_WIDTH: pong_storage_data_503 <= (fillup_transition == 1'b1) ? i_input_data[1096 % IN_WIDTH] : pong_storage_data_503 ^ i_input_data[1096 % IN_WIDTH];
                default: pong_storage_data_503 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_503;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_503 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_503;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_503 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_503;
            end
        end
    end
end

logic ping_storage_data_504;
logic pong_storage_data_504;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_504 <= 1'b0;
        pong_storage_data_504 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                458 / IN_WIDTH: ping_storage_data_504 <= (fillup_transition == 1'b1) ? i_input_data[458 % IN_WIDTH] : ping_storage_data_504 ^ i_input_data[458 % IN_WIDTH];
                560 / IN_WIDTH: ping_storage_data_504 <= (fillup_transition == 1'b1) ? i_input_data[560 % IN_WIDTH] : ping_storage_data_504 ^ i_input_data[560 % IN_WIDTH];
                710 / IN_WIDTH: ping_storage_data_504 <= (fillup_transition == 1'b1) ? i_input_data[710 % IN_WIDTH] : ping_storage_data_504 ^ i_input_data[710 % IN_WIDTH];
                1097 / IN_WIDTH: ping_storage_data_504 <= (fillup_transition == 1'b1) ? i_input_data[1097 % IN_WIDTH] : ping_storage_data_504 ^ i_input_data[1097 % IN_WIDTH];
                default: ping_storage_data_504 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_504;
                endcase
            end else begin
                case (input_count)
                458 / IN_WIDTH: pong_storage_data_504 <= (fillup_transition == 1'b1) ? i_input_data[458 % IN_WIDTH] : pong_storage_data_504 ^ i_input_data[458 % IN_WIDTH];
                560 / IN_WIDTH: pong_storage_data_504 <= (fillup_transition == 1'b1) ? i_input_data[560 % IN_WIDTH] : pong_storage_data_504 ^ i_input_data[560 % IN_WIDTH];
                710 / IN_WIDTH: pong_storage_data_504 <= (fillup_transition == 1'b1) ? i_input_data[710 % IN_WIDTH] : pong_storage_data_504 ^ i_input_data[710 % IN_WIDTH];
                1097 / IN_WIDTH: pong_storage_data_504 <= (fillup_transition == 1'b1) ? i_input_data[1097 % IN_WIDTH] : pong_storage_data_504 ^ i_input_data[1097 % IN_WIDTH];
                default: pong_storage_data_504 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_504;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_504 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_504;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_504 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_504;
            end
        end
    end
end

logic ping_storage_data_505;
logic pong_storage_data_505;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_505 <= 1'b0;
        pong_storage_data_505 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                459 / IN_WIDTH: ping_storage_data_505 <= (fillup_transition == 1'b1) ? i_input_data[459 % IN_WIDTH] : ping_storage_data_505 ^ i_input_data[459 % IN_WIDTH];
                561 / IN_WIDTH: ping_storage_data_505 <= (fillup_transition == 1'b1) ? i_input_data[561 % IN_WIDTH] : ping_storage_data_505 ^ i_input_data[561 % IN_WIDTH];
                711 / IN_WIDTH: ping_storage_data_505 <= (fillup_transition == 1'b1) ? i_input_data[711 % IN_WIDTH] : ping_storage_data_505 ^ i_input_data[711 % IN_WIDTH];
                1098 / IN_WIDTH: ping_storage_data_505 <= (fillup_transition == 1'b1) ? i_input_data[1098 % IN_WIDTH] : ping_storage_data_505 ^ i_input_data[1098 % IN_WIDTH];
                default: ping_storage_data_505 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_505;
                endcase
            end else begin
                case (input_count)
                459 / IN_WIDTH: pong_storage_data_505 <= (fillup_transition == 1'b1) ? i_input_data[459 % IN_WIDTH] : pong_storage_data_505 ^ i_input_data[459 % IN_WIDTH];
                561 / IN_WIDTH: pong_storage_data_505 <= (fillup_transition == 1'b1) ? i_input_data[561 % IN_WIDTH] : pong_storage_data_505 ^ i_input_data[561 % IN_WIDTH];
                711 / IN_WIDTH: pong_storage_data_505 <= (fillup_transition == 1'b1) ? i_input_data[711 % IN_WIDTH] : pong_storage_data_505 ^ i_input_data[711 % IN_WIDTH];
                1098 / IN_WIDTH: pong_storage_data_505 <= (fillup_transition == 1'b1) ? i_input_data[1098 % IN_WIDTH] : pong_storage_data_505 ^ i_input_data[1098 % IN_WIDTH];
                default: pong_storage_data_505 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_505;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_505 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_505;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_505 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_505;
            end
        end
    end
end

logic ping_storage_data_506;
logic pong_storage_data_506;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_506 <= 1'b0;
        pong_storage_data_506 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                460 / IN_WIDTH: ping_storage_data_506 <= (fillup_transition == 1'b1) ? i_input_data[460 % IN_WIDTH] : ping_storage_data_506 ^ i_input_data[460 % IN_WIDTH];
                562 / IN_WIDTH: ping_storage_data_506 <= (fillup_transition == 1'b1) ? i_input_data[562 % IN_WIDTH] : ping_storage_data_506 ^ i_input_data[562 % IN_WIDTH];
                712 / IN_WIDTH: ping_storage_data_506 <= (fillup_transition == 1'b1) ? i_input_data[712 % IN_WIDTH] : ping_storage_data_506 ^ i_input_data[712 % IN_WIDTH];
                1099 / IN_WIDTH: ping_storage_data_506 <= (fillup_transition == 1'b1) ? i_input_data[1099 % IN_WIDTH] : ping_storage_data_506 ^ i_input_data[1099 % IN_WIDTH];
                default: ping_storage_data_506 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_506;
                endcase
            end else begin
                case (input_count)
                460 / IN_WIDTH: pong_storage_data_506 <= (fillup_transition == 1'b1) ? i_input_data[460 % IN_WIDTH] : pong_storage_data_506 ^ i_input_data[460 % IN_WIDTH];
                562 / IN_WIDTH: pong_storage_data_506 <= (fillup_transition == 1'b1) ? i_input_data[562 % IN_WIDTH] : pong_storage_data_506 ^ i_input_data[562 % IN_WIDTH];
                712 / IN_WIDTH: pong_storage_data_506 <= (fillup_transition == 1'b1) ? i_input_data[712 % IN_WIDTH] : pong_storage_data_506 ^ i_input_data[712 % IN_WIDTH];
                1099 / IN_WIDTH: pong_storage_data_506 <= (fillup_transition == 1'b1) ? i_input_data[1099 % IN_WIDTH] : pong_storage_data_506 ^ i_input_data[1099 % IN_WIDTH];
                default: pong_storage_data_506 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_506;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_506 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_506;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_506 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_506;
            end
        end
    end
end

logic ping_storage_data_507;
logic pong_storage_data_507;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_507 <= 1'b0;
        pong_storage_data_507 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                461 / IN_WIDTH: ping_storage_data_507 <= (fillup_transition == 1'b1) ? i_input_data[461 % IN_WIDTH] : ping_storage_data_507 ^ i_input_data[461 % IN_WIDTH];
                563 / IN_WIDTH: ping_storage_data_507 <= (fillup_transition == 1'b1) ? i_input_data[563 % IN_WIDTH] : ping_storage_data_507 ^ i_input_data[563 % IN_WIDTH];
                713 / IN_WIDTH: ping_storage_data_507 <= (fillup_transition == 1'b1) ? i_input_data[713 % IN_WIDTH] : ping_storage_data_507 ^ i_input_data[713 % IN_WIDTH];
                1100 / IN_WIDTH: ping_storage_data_507 <= (fillup_transition == 1'b1) ? i_input_data[1100 % IN_WIDTH] : ping_storage_data_507 ^ i_input_data[1100 % IN_WIDTH];
                default: ping_storage_data_507 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_507;
                endcase
            end else begin
                case (input_count)
                461 / IN_WIDTH: pong_storage_data_507 <= (fillup_transition == 1'b1) ? i_input_data[461 % IN_WIDTH] : pong_storage_data_507 ^ i_input_data[461 % IN_WIDTH];
                563 / IN_WIDTH: pong_storage_data_507 <= (fillup_transition == 1'b1) ? i_input_data[563 % IN_WIDTH] : pong_storage_data_507 ^ i_input_data[563 % IN_WIDTH];
                713 / IN_WIDTH: pong_storage_data_507 <= (fillup_transition == 1'b1) ? i_input_data[713 % IN_WIDTH] : pong_storage_data_507 ^ i_input_data[713 % IN_WIDTH];
                1100 / IN_WIDTH: pong_storage_data_507 <= (fillup_transition == 1'b1) ? i_input_data[1100 % IN_WIDTH] : pong_storage_data_507 ^ i_input_data[1100 % IN_WIDTH];
                default: pong_storage_data_507 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_507;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_507 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_507;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_507 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_507;
            end
        end
    end
end

logic ping_storage_data_508;
logic pong_storage_data_508;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_508 <= 1'b0;
        pong_storage_data_508 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                462 / IN_WIDTH: ping_storage_data_508 <= (fillup_transition == 1'b1) ? i_input_data[462 % IN_WIDTH] : ping_storage_data_508 ^ i_input_data[462 % IN_WIDTH];
                564 / IN_WIDTH: ping_storage_data_508 <= (fillup_transition == 1'b1) ? i_input_data[564 % IN_WIDTH] : ping_storage_data_508 ^ i_input_data[564 % IN_WIDTH];
                714 / IN_WIDTH: ping_storage_data_508 <= (fillup_transition == 1'b1) ? i_input_data[714 % IN_WIDTH] : ping_storage_data_508 ^ i_input_data[714 % IN_WIDTH];
                1101 / IN_WIDTH: ping_storage_data_508 <= (fillup_transition == 1'b1) ? i_input_data[1101 % IN_WIDTH] : ping_storage_data_508 ^ i_input_data[1101 % IN_WIDTH];
                default: ping_storage_data_508 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_508;
                endcase
            end else begin
                case (input_count)
                462 / IN_WIDTH: pong_storage_data_508 <= (fillup_transition == 1'b1) ? i_input_data[462 % IN_WIDTH] : pong_storage_data_508 ^ i_input_data[462 % IN_WIDTH];
                564 / IN_WIDTH: pong_storage_data_508 <= (fillup_transition == 1'b1) ? i_input_data[564 % IN_WIDTH] : pong_storage_data_508 ^ i_input_data[564 % IN_WIDTH];
                714 / IN_WIDTH: pong_storage_data_508 <= (fillup_transition == 1'b1) ? i_input_data[714 % IN_WIDTH] : pong_storage_data_508 ^ i_input_data[714 % IN_WIDTH];
                1101 / IN_WIDTH: pong_storage_data_508 <= (fillup_transition == 1'b1) ? i_input_data[1101 % IN_WIDTH] : pong_storage_data_508 ^ i_input_data[1101 % IN_WIDTH];
                default: pong_storage_data_508 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_508;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_508 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_508;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_508 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_508;
            end
        end
    end
end

logic ping_storage_data_509;
logic pong_storage_data_509;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_509 <= 1'b0;
        pong_storage_data_509 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                463 / IN_WIDTH: ping_storage_data_509 <= (fillup_transition == 1'b1) ? i_input_data[463 % IN_WIDTH] : ping_storage_data_509 ^ i_input_data[463 % IN_WIDTH];
                565 / IN_WIDTH: ping_storage_data_509 <= (fillup_transition == 1'b1) ? i_input_data[565 % IN_WIDTH] : ping_storage_data_509 ^ i_input_data[565 % IN_WIDTH];
                715 / IN_WIDTH: ping_storage_data_509 <= (fillup_transition == 1'b1) ? i_input_data[715 % IN_WIDTH] : ping_storage_data_509 ^ i_input_data[715 % IN_WIDTH];
                1102 / IN_WIDTH: ping_storage_data_509 <= (fillup_transition == 1'b1) ? i_input_data[1102 % IN_WIDTH] : ping_storage_data_509 ^ i_input_data[1102 % IN_WIDTH];
                default: ping_storage_data_509 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_509;
                endcase
            end else begin
                case (input_count)
                463 / IN_WIDTH: pong_storage_data_509 <= (fillup_transition == 1'b1) ? i_input_data[463 % IN_WIDTH] : pong_storage_data_509 ^ i_input_data[463 % IN_WIDTH];
                565 / IN_WIDTH: pong_storage_data_509 <= (fillup_transition == 1'b1) ? i_input_data[565 % IN_WIDTH] : pong_storage_data_509 ^ i_input_data[565 % IN_WIDTH];
                715 / IN_WIDTH: pong_storage_data_509 <= (fillup_transition == 1'b1) ? i_input_data[715 % IN_WIDTH] : pong_storage_data_509 ^ i_input_data[715 % IN_WIDTH];
                1102 / IN_WIDTH: pong_storage_data_509 <= (fillup_transition == 1'b1) ? i_input_data[1102 % IN_WIDTH] : pong_storage_data_509 ^ i_input_data[1102 % IN_WIDTH];
                default: pong_storage_data_509 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_509;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_509 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_509;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_509 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_509;
            end
        end
    end
end

logic ping_storage_data_510;
logic pong_storage_data_510;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_510 <= 1'b0;
        pong_storage_data_510 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                464 / IN_WIDTH: ping_storage_data_510 <= (fillup_transition == 1'b1) ? i_input_data[464 % IN_WIDTH] : ping_storage_data_510 ^ i_input_data[464 % IN_WIDTH];
                566 / IN_WIDTH: ping_storage_data_510 <= (fillup_transition == 1'b1) ? i_input_data[566 % IN_WIDTH] : ping_storage_data_510 ^ i_input_data[566 % IN_WIDTH];
                716 / IN_WIDTH: ping_storage_data_510 <= (fillup_transition == 1'b1) ? i_input_data[716 % IN_WIDTH] : ping_storage_data_510 ^ i_input_data[716 % IN_WIDTH];
                1103 / IN_WIDTH: ping_storage_data_510 <= (fillup_transition == 1'b1) ? i_input_data[1103 % IN_WIDTH] : ping_storage_data_510 ^ i_input_data[1103 % IN_WIDTH];
                default: ping_storage_data_510 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_510;
                endcase
            end else begin
                case (input_count)
                464 / IN_WIDTH: pong_storage_data_510 <= (fillup_transition == 1'b1) ? i_input_data[464 % IN_WIDTH] : pong_storage_data_510 ^ i_input_data[464 % IN_WIDTH];
                566 / IN_WIDTH: pong_storage_data_510 <= (fillup_transition == 1'b1) ? i_input_data[566 % IN_WIDTH] : pong_storage_data_510 ^ i_input_data[566 % IN_WIDTH];
                716 / IN_WIDTH: pong_storage_data_510 <= (fillup_transition == 1'b1) ? i_input_data[716 % IN_WIDTH] : pong_storage_data_510 ^ i_input_data[716 % IN_WIDTH];
                1103 / IN_WIDTH: pong_storage_data_510 <= (fillup_transition == 1'b1) ? i_input_data[1103 % IN_WIDTH] : pong_storage_data_510 ^ i_input_data[1103 % IN_WIDTH];
                default: pong_storage_data_510 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_510;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_510 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_510;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_510 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_510;
            end
        end
    end
end

logic ping_storage_data_511;
logic pong_storage_data_511;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_511 <= 1'b0;
        pong_storage_data_511 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                465 / IN_WIDTH: ping_storage_data_511 <= (fillup_transition == 1'b1) ? i_input_data[465 % IN_WIDTH] : ping_storage_data_511 ^ i_input_data[465 % IN_WIDTH];
                567 / IN_WIDTH: ping_storage_data_511 <= (fillup_transition == 1'b1) ? i_input_data[567 % IN_WIDTH] : ping_storage_data_511 ^ i_input_data[567 % IN_WIDTH];
                717 / IN_WIDTH: ping_storage_data_511 <= (fillup_transition == 1'b1) ? i_input_data[717 % IN_WIDTH] : ping_storage_data_511 ^ i_input_data[717 % IN_WIDTH];
                1104 / IN_WIDTH: ping_storage_data_511 <= (fillup_transition == 1'b1) ? i_input_data[1104 % IN_WIDTH] : ping_storage_data_511 ^ i_input_data[1104 % IN_WIDTH];
                default: ping_storage_data_511 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_511;
                endcase
            end else begin
                case (input_count)
                465 / IN_WIDTH: pong_storage_data_511 <= (fillup_transition == 1'b1) ? i_input_data[465 % IN_WIDTH] : pong_storage_data_511 ^ i_input_data[465 % IN_WIDTH];
                567 / IN_WIDTH: pong_storage_data_511 <= (fillup_transition == 1'b1) ? i_input_data[567 % IN_WIDTH] : pong_storage_data_511 ^ i_input_data[567 % IN_WIDTH];
                717 / IN_WIDTH: pong_storage_data_511 <= (fillup_transition == 1'b1) ? i_input_data[717 % IN_WIDTH] : pong_storage_data_511 ^ i_input_data[717 % IN_WIDTH];
                1104 / IN_WIDTH: pong_storage_data_511 <= (fillup_transition == 1'b1) ? i_input_data[1104 % IN_WIDTH] : pong_storage_data_511 ^ i_input_data[1104 % IN_WIDTH];
                default: pong_storage_data_511 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_511;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_511 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_511;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_511 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_511;
            end
        end
    end
end

logic ping_storage_data_512;
logic pong_storage_data_512;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_512 <= 1'b0;
        pong_storage_data_512 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                466 / IN_WIDTH: ping_storage_data_512 <= (fillup_transition == 1'b1) ? i_input_data[466 % IN_WIDTH] : ping_storage_data_512 ^ i_input_data[466 % IN_WIDTH];
                568 / IN_WIDTH: ping_storage_data_512 <= (fillup_transition == 1'b1) ? i_input_data[568 % IN_WIDTH] : ping_storage_data_512 ^ i_input_data[568 % IN_WIDTH];
                718 / IN_WIDTH: ping_storage_data_512 <= (fillup_transition == 1'b1) ? i_input_data[718 % IN_WIDTH] : ping_storage_data_512 ^ i_input_data[718 % IN_WIDTH];
                1105 / IN_WIDTH: ping_storage_data_512 <= (fillup_transition == 1'b1) ? i_input_data[1105 % IN_WIDTH] : ping_storage_data_512 ^ i_input_data[1105 % IN_WIDTH];
                default: ping_storage_data_512 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_512;
                endcase
            end else begin
                case (input_count)
                466 / IN_WIDTH: pong_storage_data_512 <= (fillup_transition == 1'b1) ? i_input_data[466 % IN_WIDTH] : pong_storage_data_512 ^ i_input_data[466 % IN_WIDTH];
                568 / IN_WIDTH: pong_storage_data_512 <= (fillup_transition == 1'b1) ? i_input_data[568 % IN_WIDTH] : pong_storage_data_512 ^ i_input_data[568 % IN_WIDTH];
                718 / IN_WIDTH: pong_storage_data_512 <= (fillup_transition == 1'b1) ? i_input_data[718 % IN_WIDTH] : pong_storage_data_512 ^ i_input_data[718 % IN_WIDTH];
                1105 / IN_WIDTH: pong_storage_data_512 <= (fillup_transition == 1'b1) ? i_input_data[1105 % IN_WIDTH] : pong_storage_data_512 ^ i_input_data[1105 % IN_WIDTH];
                default: pong_storage_data_512 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_512;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_512 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_512;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_512 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_512;
            end
        end
    end
end

logic ping_storage_data_513;
logic pong_storage_data_513;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_513 <= 1'b0;
        pong_storage_data_513 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                467 / IN_WIDTH: ping_storage_data_513 <= (fillup_transition == 1'b1) ? i_input_data[467 % IN_WIDTH] : ping_storage_data_513 ^ i_input_data[467 % IN_WIDTH];
                569 / IN_WIDTH: ping_storage_data_513 <= (fillup_transition == 1'b1) ? i_input_data[569 % IN_WIDTH] : ping_storage_data_513 ^ i_input_data[569 % IN_WIDTH];
                719 / IN_WIDTH: ping_storage_data_513 <= (fillup_transition == 1'b1) ? i_input_data[719 % IN_WIDTH] : ping_storage_data_513 ^ i_input_data[719 % IN_WIDTH];
                1106 / IN_WIDTH: ping_storage_data_513 <= (fillup_transition == 1'b1) ? i_input_data[1106 % IN_WIDTH] : ping_storage_data_513 ^ i_input_data[1106 % IN_WIDTH];
                default: ping_storage_data_513 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_513;
                endcase
            end else begin
                case (input_count)
                467 / IN_WIDTH: pong_storage_data_513 <= (fillup_transition == 1'b1) ? i_input_data[467 % IN_WIDTH] : pong_storage_data_513 ^ i_input_data[467 % IN_WIDTH];
                569 / IN_WIDTH: pong_storage_data_513 <= (fillup_transition == 1'b1) ? i_input_data[569 % IN_WIDTH] : pong_storage_data_513 ^ i_input_data[569 % IN_WIDTH];
                719 / IN_WIDTH: pong_storage_data_513 <= (fillup_transition == 1'b1) ? i_input_data[719 % IN_WIDTH] : pong_storage_data_513 ^ i_input_data[719 % IN_WIDTH];
                1106 / IN_WIDTH: pong_storage_data_513 <= (fillup_transition == 1'b1) ? i_input_data[1106 % IN_WIDTH] : pong_storage_data_513 ^ i_input_data[1106 % IN_WIDTH];
                default: pong_storage_data_513 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_513;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_513 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_513;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_513 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_513;
            end
        end
    end
end

logic ping_storage_data_514;
logic pong_storage_data_514;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_514 <= 1'b0;
        pong_storage_data_514 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                468 / IN_WIDTH: ping_storage_data_514 <= (fillup_transition == 1'b1) ? i_input_data[468 % IN_WIDTH] : ping_storage_data_514 ^ i_input_data[468 % IN_WIDTH];
                570 / IN_WIDTH: ping_storage_data_514 <= (fillup_transition == 1'b1) ? i_input_data[570 % IN_WIDTH] : ping_storage_data_514 ^ i_input_data[570 % IN_WIDTH];
                720 / IN_WIDTH: ping_storage_data_514 <= (fillup_transition == 1'b1) ? i_input_data[720 % IN_WIDTH] : ping_storage_data_514 ^ i_input_data[720 % IN_WIDTH];
                1107 / IN_WIDTH: ping_storage_data_514 <= (fillup_transition == 1'b1) ? i_input_data[1107 % IN_WIDTH] : ping_storage_data_514 ^ i_input_data[1107 % IN_WIDTH];
                default: ping_storage_data_514 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_514;
                endcase
            end else begin
                case (input_count)
                468 / IN_WIDTH: pong_storage_data_514 <= (fillup_transition == 1'b1) ? i_input_data[468 % IN_WIDTH] : pong_storage_data_514 ^ i_input_data[468 % IN_WIDTH];
                570 / IN_WIDTH: pong_storage_data_514 <= (fillup_transition == 1'b1) ? i_input_data[570 % IN_WIDTH] : pong_storage_data_514 ^ i_input_data[570 % IN_WIDTH];
                720 / IN_WIDTH: pong_storage_data_514 <= (fillup_transition == 1'b1) ? i_input_data[720 % IN_WIDTH] : pong_storage_data_514 ^ i_input_data[720 % IN_WIDTH];
                1107 / IN_WIDTH: pong_storage_data_514 <= (fillup_transition == 1'b1) ? i_input_data[1107 % IN_WIDTH] : pong_storage_data_514 ^ i_input_data[1107 % IN_WIDTH];
                default: pong_storage_data_514 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_514;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_514 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_514;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_514 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_514;
            end
        end
    end
end

logic ping_storage_data_515;
logic pong_storage_data_515;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_515 <= 1'b0;
        pong_storage_data_515 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                469 / IN_WIDTH: ping_storage_data_515 <= (fillup_transition == 1'b1) ? i_input_data[469 % IN_WIDTH] : ping_storage_data_515 ^ i_input_data[469 % IN_WIDTH];
                571 / IN_WIDTH: ping_storage_data_515 <= (fillup_transition == 1'b1) ? i_input_data[571 % IN_WIDTH] : ping_storage_data_515 ^ i_input_data[571 % IN_WIDTH];
                721 / IN_WIDTH: ping_storage_data_515 <= (fillup_transition == 1'b1) ? i_input_data[721 % IN_WIDTH] : ping_storage_data_515 ^ i_input_data[721 % IN_WIDTH];
                1108 / IN_WIDTH: ping_storage_data_515 <= (fillup_transition == 1'b1) ? i_input_data[1108 % IN_WIDTH] : ping_storage_data_515 ^ i_input_data[1108 % IN_WIDTH];
                default: ping_storage_data_515 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_515;
                endcase
            end else begin
                case (input_count)
                469 / IN_WIDTH: pong_storage_data_515 <= (fillup_transition == 1'b1) ? i_input_data[469 % IN_WIDTH] : pong_storage_data_515 ^ i_input_data[469 % IN_WIDTH];
                571 / IN_WIDTH: pong_storage_data_515 <= (fillup_transition == 1'b1) ? i_input_data[571 % IN_WIDTH] : pong_storage_data_515 ^ i_input_data[571 % IN_WIDTH];
                721 / IN_WIDTH: pong_storage_data_515 <= (fillup_transition == 1'b1) ? i_input_data[721 % IN_WIDTH] : pong_storage_data_515 ^ i_input_data[721 % IN_WIDTH];
                1108 / IN_WIDTH: pong_storage_data_515 <= (fillup_transition == 1'b1) ? i_input_data[1108 % IN_WIDTH] : pong_storage_data_515 ^ i_input_data[1108 % IN_WIDTH];
                default: pong_storage_data_515 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_515;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_515 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_515;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_515 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_515;
            end
        end
    end
end

logic ping_storage_data_516;
logic pong_storage_data_516;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_516 <= 1'b0;
        pong_storage_data_516 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                470 / IN_WIDTH: ping_storage_data_516 <= (fillup_transition == 1'b1) ? i_input_data[470 % IN_WIDTH] : ping_storage_data_516 ^ i_input_data[470 % IN_WIDTH];
                572 / IN_WIDTH: ping_storage_data_516 <= (fillup_transition == 1'b1) ? i_input_data[572 % IN_WIDTH] : ping_storage_data_516 ^ i_input_data[572 % IN_WIDTH];
                722 / IN_WIDTH: ping_storage_data_516 <= (fillup_transition == 1'b1) ? i_input_data[722 % IN_WIDTH] : ping_storage_data_516 ^ i_input_data[722 % IN_WIDTH];
                1109 / IN_WIDTH: ping_storage_data_516 <= (fillup_transition == 1'b1) ? i_input_data[1109 % IN_WIDTH] : ping_storage_data_516 ^ i_input_data[1109 % IN_WIDTH];
                default: ping_storage_data_516 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_516;
                endcase
            end else begin
                case (input_count)
                470 / IN_WIDTH: pong_storage_data_516 <= (fillup_transition == 1'b1) ? i_input_data[470 % IN_WIDTH] : pong_storage_data_516 ^ i_input_data[470 % IN_WIDTH];
                572 / IN_WIDTH: pong_storage_data_516 <= (fillup_transition == 1'b1) ? i_input_data[572 % IN_WIDTH] : pong_storage_data_516 ^ i_input_data[572 % IN_WIDTH];
                722 / IN_WIDTH: pong_storage_data_516 <= (fillup_transition == 1'b1) ? i_input_data[722 % IN_WIDTH] : pong_storage_data_516 ^ i_input_data[722 % IN_WIDTH];
                1109 / IN_WIDTH: pong_storage_data_516 <= (fillup_transition == 1'b1) ? i_input_data[1109 % IN_WIDTH] : pong_storage_data_516 ^ i_input_data[1109 % IN_WIDTH];
                default: pong_storage_data_516 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_516;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_516 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_516;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_516 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_516;
            end
        end
    end
end

logic ping_storage_data_517;
logic pong_storage_data_517;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_517 <= 1'b0;
        pong_storage_data_517 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                471 / IN_WIDTH: ping_storage_data_517 <= (fillup_transition == 1'b1) ? i_input_data[471 % IN_WIDTH] : ping_storage_data_517 ^ i_input_data[471 % IN_WIDTH];
                573 / IN_WIDTH: ping_storage_data_517 <= (fillup_transition == 1'b1) ? i_input_data[573 % IN_WIDTH] : ping_storage_data_517 ^ i_input_data[573 % IN_WIDTH];
                723 / IN_WIDTH: ping_storage_data_517 <= (fillup_transition == 1'b1) ? i_input_data[723 % IN_WIDTH] : ping_storage_data_517 ^ i_input_data[723 % IN_WIDTH];
                1110 / IN_WIDTH: ping_storage_data_517 <= (fillup_transition == 1'b1) ? i_input_data[1110 % IN_WIDTH] : ping_storage_data_517 ^ i_input_data[1110 % IN_WIDTH];
                default: ping_storage_data_517 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_517;
                endcase
            end else begin
                case (input_count)
                471 / IN_WIDTH: pong_storage_data_517 <= (fillup_transition == 1'b1) ? i_input_data[471 % IN_WIDTH] : pong_storage_data_517 ^ i_input_data[471 % IN_WIDTH];
                573 / IN_WIDTH: pong_storage_data_517 <= (fillup_transition == 1'b1) ? i_input_data[573 % IN_WIDTH] : pong_storage_data_517 ^ i_input_data[573 % IN_WIDTH];
                723 / IN_WIDTH: pong_storage_data_517 <= (fillup_transition == 1'b1) ? i_input_data[723 % IN_WIDTH] : pong_storage_data_517 ^ i_input_data[723 % IN_WIDTH];
                1110 / IN_WIDTH: pong_storage_data_517 <= (fillup_transition == 1'b1) ? i_input_data[1110 % IN_WIDTH] : pong_storage_data_517 ^ i_input_data[1110 % IN_WIDTH];
                default: pong_storage_data_517 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_517;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_517 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_517;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_517 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_517;
            end
        end
    end
end

logic ping_storage_data_518;
logic pong_storage_data_518;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_518 <= 1'b0;
        pong_storage_data_518 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                472 / IN_WIDTH: ping_storage_data_518 <= (fillup_transition == 1'b1) ? i_input_data[472 % IN_WIDTH] : ping_storage_data_518 ^ i_input_data[472 % IN_WIDTH];
                574 / IN_WIDTH: ping_storage_data_518 <= (fillup_transition == 1'b1) ? i_input_data[574 % IN_WIDTH] : ping_storage_data_518 ^ i_input_data[574 % IN_WIDTH];
                724 / IN_WIDTH: ping_storage_data_518 <= (fillup_transition == 1'b1) ? i_input_data[724 % IN_WIDTH] : ping_storage_data_518 ^ i_input_data[724 % IN_WIDTH];
                1111 / IN_WIDTH: ping_storage_data_518 <= (fillup_transition == 1'b1) ? i_input_data[1111 % IN_WIDTH] : ping_storage_data_518 ^ i_input_data[1111 % IN_WIDTH];
                default: ping_storage_data_518 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_518;
                endcase
            end else begin
                case (input_count)
                472 / IN_WIDTH: pong_storage_data_518 <= (fillup_transition == 1'b1) ? i_input_data[472 % IN_WIDTH] : pong_storage_data_518 ^ i_input_data[472 % IN_WIDTH];
                574 / IN_WIDTH: pong_storage_data_518 <= (fillup_transition == 1'b1) ? i_input_data[574 % IN_WIDTH] : pong_storage_data_518 ^ i_input_data[574 % IN_WIDTH];
                724 / IN_WIDTH: pong_storage_data_518 <= (fillup_transition == 1'b1) ? i_input_data[724 % IN_WIDTH] : pong_storage_data_518 ^ i_input_data[724 % IN_WIDTH];
                1111 / IN_WIDTH: pong_storage_data_518 <= (fillup_transition == 1'b1) ? i_input_data[1111 % IN_WIDTH] : pong_storage_data_518 ^ i_input_data[1111 % IN_WIDTH];
                default: pong_storage_data_518 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_518;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_518 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_518;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_518 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_518;
            end
        end
    end
end

logic ping_storage_data_519;
logic pong_storage_data_519;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_519 <= 1'b0;
        pong_storage_data_519 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                473 / IN_WIDTH: ping_storage_data_519 <= (fillup_transition == 1'b1) ? i_input_data[473 % IN_WIDTH] : ping_storage_data_519 ^ i_input_data[473 % IN_WIDTH];
                575 / IN_WIDTH: ping_storage_data_519 <= (fillup_transition == 1'b1) ? i_input_data[575 % IN_WIDTH] : ping_storage_data_519 ^ i_input_data[575 % IN_WIDTH];
                725 / IN_WIDTH: ping_storage_data_519 <= (fillup_transition == 1'b1) ? i_input_data[725 % IN_WIDTH] : ping_storage_data_519 ^ i_input_data[725 % IN_WIDTH];
                1112 / IN_WIDTH: ping_storage_data_519 <= (fillup_transition == 1'b1) ? i_input_data[1112 % IN_WIDTH] : ping_storage_data_519 ^ i_input_data[1112 % IN_WIDTH];
                default: ping_storage_data_519 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_519;
                endcase
            end else begin
                case (input_count)
                473 / IN_WIDTH: pong_storage_data_519 <= (fillup_transition == 1'b1) ? i_input_data[473 % IN_WIDTH] : pong_storage_data_519 ^ i_input_data[473 % IN_WIDTH];
                575 / IN_WIDTH: pong_storage_data_519 <= (fillup_transition == 1'b1) ? i_input_data[575 % IN_WIDTH] : pong_storage_data_519 ^ i_input_data[575 % IN_WIDTH];
                725 / IN_WIDTH: pong_storage_data_519 <= (fillup_transition == 1'b1) ? i_input_data[725 % IN_WIDTH] : pong_storage_data_519 ^ i_input_data[725 % IN_WIDTH];
                1112 / IN_WIDTH: pong_storage_data_519 <= (fillup_transition == 1'b1) ? i_input_data[1112 % IN_WIDTH] : pong_storage_data_519 ^ i_input_data[1112 % IN_WIDTH];
                default: pong_storage_data_519 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_519;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_519 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_519;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_519 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_519;
            end
        end
    end
end

logic ping_storage_data_520;
logic pong_storage_data_520;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_520 <= 1'b0;
        pong_storage_data_520 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                474 / IN_WIDTH: ping_storage_data_520 <= (fillup_transition == 1'b1) ? i_input_data[474 % IN_WIDTH] : ping_storage_data_520 ^ i_input_data[474 % IN_WIDTH];
                480 / IN_WIDTH: ping_storage_data_520 <= (fillup_transition == 1'b1) ? i_input_data[480 % IN_WIDTH] : ping_storage_data_520 ^ i_input_data[480 % IN_WIDTH];
                726 / IN_WIDTH: ping_storage_data_520 <= (fillup_transition == 1'b1) ? i_input_data[726 % IN_WIDTH] : ping_storage_data_520 ^ i_input_data[726 % IN_WIDTH];
                1113 / IN_WIDTH: ping_storage_data_520 <= (fillup_transition == 1'b1) ? i_input_data[1113 % IN_WIDTH] : ping_storage_data_520 ^ i_input_data[1113 % IN_WIDTH];
                default: ping_storage_data_520 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_520;
                endcase
            end else begin
                case (input_count)
                474 / IN_WIDTH: pong_storage_data_520 <= (fillup_transition == 1'b1) ? i_input_data[474 % IN_WIDTH] : pong_storage_data_520 ^ i_input_data[474 % IN_WIDTH];
                480 / IN_WIDTH: pong_storage_data_520 <= (fillup_transition == 1'b1) ? i_input_data[480 % IN_WIDTH] : pong_storage_data_520 ^ i_input_data[480 % IN_WIDTH];
                726 / IN_WIDTH: pong_storage_data_520 <= (fillup_transition == 1'b1) ? i_input_data[726 % IN_WIDTH] : pong_storage_data_520 ^ i_input_data[726 % IN_WIDTH];
                1113 / IN_WIDTH: pong_storage_data_520 <= (fillup_transition == 1'b1) ? i_input_data[1113 % IN_WIDTH] : pong_storage_data_520 ^ i_input_data[1113 % IN_WIDTH];
                default: pong_storage_data_520 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_520;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_520 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_520;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_520 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_520;
            end
        end
    end
end

logic ping_storage_data_521;
logic pong_storage_data_521;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_521 <= 1'b0;
        pong_storage_data_521 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                475 / IN_WIDTH: ping_storage_data_521 <= (fillup_transition == 1'b1) ? i_input_data[475 % IN_WIDTH] : ping_storage_data_521 ^ i_input_data[475 % IN_WIDTH];
                481 / IN_WIDTH: ping_storage_data_521 <= (fillup_transition == 1'b1) ? i_input_data[481 % IN_WIDTH] : ping_storage_data_521 ^ i_input_data[481 % IN_WIDTH];
                727 / IN_WIDTH: ping_storage_data_521 <= (fillup_transition == 1'b1) ? i_input_data[727 % IN_WIDTH] : ping_storage_data_521 ^ i_input_data[727 % IN_WIDTH];
                1114 / IN_WIDTH: ping_storage_data_521 <= (fillup_transition == 1'b1) ? i_input_data[1114 % IN_WIDTH] : ping_storage_data_521 ^ i_input_data[1114 % IN_WIDTH];
                default: ping_storage_data_521 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_521;
                endcase
            end else begin
                case (input_count)
                475 / IN_WIDTH: pong_storage_data_521 <= (fillup_transition == 1'b1) ? i_input_data[475 % IN_WIDTH] : pong_storage_data_521 ^ i_input_data[475 % IN_WIDTH];
                481 / IN_WIDTH: pong_storage_data_521 <= (fillup_transition == 1'b1) ? i_input_data[481 % IN_WIDTH] : pong_storage_data_521 ^ i_input_data[481 % IN_WIDTH];
                727 / IN_WIDTH: pong_storage_data_521 <= (fillup_transition == 1'b1) ? i_input_data[727 % IN_WIDTH] : pong_storage_data_521 ^ i_input_data[727 % IN_WIDTH];
                1114 / IN_WIDTH: pong_storage_data_521 <= (fillup_transition == 1'b1) ? i_input_data[1114 % IN_WIDTH] : pong_storage_data_521 ^ i_input_data[1114 % IN_WIDTH];
                default: pong_storage_data_521 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_521;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_521 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_521;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_521 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_521;
            end
        end
    end
end

logic ping_storage_data_522;
logic pong_storage_data_522;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_522 <= 1'b0;
        pong_storage_data_522 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                476 / IN_WIDTH: ping_storage_data_522 <= (fillup_transition == 1'b1) ? i_input_data[476 % IN_WIDTH] : ping_storage_data_522 ^ i_input_data[476 % IN_WIDTH];
                482 / IN_WIDTH: ping_storage_data_522 <= (fillup_transition == 1'b1) ? i_input_data[482 % IN_WIDTH] : ping_storage_data_522 ^ i_input_data[482 % IN_WIDTH];
                728 / IN_WIDTH: ping_storage_data_522 <= (fillup_transition == 1'b1) ? i_input_data[728 % IN_WIDTH] : ping_storage_data_522 ^ i_input_data[728 % IN_WIDTH];
                1115 / IN_WIDTH: ping_storage_data_522 <= (fillup_transition == 1'b1) ? i_input_data[1115 % IN_WIDTH] : ping_storage_data_522 ^ i_input_data[1115 % IN_WIDTH];
                default: ping_storage_data_522 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_522;
                endcase
            end else begin
                case (input_count)
                476 / IN_WIDTH: pong_storage_data_522 <= (fillup_transition == 1'b1) ? i_input_data[476 % IN_WIDTH] : pong_storage_data_522 ^ i_input_data[476 % IN_WIDTH];
                482 / IN_WIDTH: pong_storage_data_522 <= (fillup_transition == 1'b1) ? i_input_data[482 % IN_WIDTH] : pong_storage_data_522 ^ i_input_data[482 % IN_WIDTH];
                728 / IN_WIDTH: pong_storage_data_522 <= (fillup_transition == 1'b1) ? i_input_data[728 % IN_WIDTH] : pong_storage_data_522 ^ i_input_data[728 % IN_WIDTH];
                1115 / IN_WIDTH: pong_storage_data_522 <= (fillup_transition == 1'b1) ? i_input_data[1115 % IN_WIDTH] : pong_storage_data_522 ^ i_input_data[1115 % IN_WIDTH];
                default: pong_storage_data_522 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_522;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_522 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_522;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_522 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_522;
            end
        end
    end
end

logic ping_storage_data_523;
logic pong_storage_data_523;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_523 <= 1'b0;
        pong_storage_data_523 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                477 / IN_WIDTH: ping_storage_data_523 <= (fillup_transition == 1'b1) ? i_input_data[477 % IN_WIDTH] : ping_storage_data_523 ^ i_input_data[477 % IN_WIDTH];
                483 / IN_WIDTH: ping_storage_data_523 <= (fillup_transition == 1'b1) ? i_input_data[483 % IN_WIDTH] : ping_storage_data_523 ^ i_input_data[483 % IN_WIDTH];
                729 / IN_WIDTH: ping_storage_data_523 <= (fillup_transition == 1'b1) ? i_input_data[729 % IN_WIDTH] : ping_storage_data_523 ^ i_input_data[729 % IN_WIDTH];
                1116 / IN_WIDTH: ping_storage_data_523 <= (fillup_transition == 1'b1) ? i_input_data[1116 % IN_WIDTH] : ping_storage_data_523 ^ i_input_data[1116 % IN_WIDTH];
                default: ping_storage_data_523 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_523;
                endcase
            end else begin
                case (input_count)
                477 / IN_WIDTH: pong_storage_data_523 <= (fillup_transition == 1'b1) ? i_input_data[477 % IN_WIDTH] : pong_storage_data_523 ^ i_input_data[477 % IN_WIDTH];
                483 / IN_WIDTH: pong_storage_data_523 <= (fillup_transition == 1'b1) ? i_input_data[483 % IN_WIDTH] : pong_storage_data_523 ^ i_input_data[483 % IN_WIDTH];
                729 / IN_WIDTH: pong_storage_data_523 <= (fillup_transition == 1'b1) ? i_input_data[729 % IN_WIDTH] : pong_storage_data_523 ^ i_input_data[729 % IN_WIDTH];
                1116 / IN_WIDTH: pong_storage_data_523 <= (fillup_transition == 1'b1) ? i_input_data[1116 % IN_WIDTH] : pong_storage_data_523 ^ i_input_data[1116 % IN_WIDTH];
                default: pong_storage_data_523 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_523;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_523 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_523;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_523 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_523;
            end
        end
    end
end

logic ping_storage_data_524;
logic pong_storage_data_524;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_524 <= 1'b0;
        pong_storage_data_524 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                478 / IN_WIDTH: ping_storage_data_524 <= (fillup_transition == 1'b1) ? i_input_data[478 % IN_WIDTH] : ping_storage_data_524 ^ i_input_data[478 % IN_WIDTH];
                484 / IN_WIDTH: ping_storage_data_524 <= (fillup_transition == 1'b1) ? i_input_data[484 % IN_WIDTH] : ping_storage_data_524 ^ i_input_data[484 % IN_WIDTH];
                730 / IN_WIDTH: ping_storage_data_524 <= (fillup_transition == 1'b1) ? i_input_data[730 % IN_WIDTH] : ping_storage_data_524 ^ i_input_data[730 % IN_WIDTH];
                1117 / IN_WIDTH: ping_storage_data_524 <= (fillup_transition == 1'b1) ? i_input_data[1117 % IN_WIDTH] : ping_storage_data_524 ^ i_input_data[1117 % IN_WIDTH];
                default: ping_storage_data_524 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_524;
                endcase
            end else begin
                case (input_count)
                478 / IN_WIDTH: pong_storage_data_524 <= (fillup_transition == 1'b1) ? i_input_data[478 % IN_WIDTH] : pong_storage_data_524 ^ i_input_data[478 % IN_WIDTH];
                484 / IN_WIDTH: pong_storage_data_524 <= (fillup_transition == 1'b1) ? i_input_data[484 % IN_WIDTH] : pong_storage_data_524 ^ i_input_data[484 % IN_WIDTH];
                730 / IN_WIDTH: pong_storage_data_524 <= (fillup_transition == 1'b1) ? i_input_data[730 % IN_WIDTH] : pong_storage_data_524 ^ i_input_data[730 % IN_WIDTH];
                1117 / IN_WIDTH: pong_storage_data_524 <= (fillup_transition == 1'b1) ? i_input_data[1117 % IN_WIDTH] : pong_storage_data_524 ^ i_input_data[1117 % IN_WIDTH];
                default: pong_storage_data_524 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_524;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_524 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_524;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_524 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_524;
            end
        end
    end
end

logic ping_storage_data_525;
logic pong_storage_data_525;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_525 <= 1'b0;
        pong_storage_data_525 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                479 / IN_WIDTH: ping_storage_data_525 <= (fillup_transition == 1'b1) ? i_input_data[479 % IN_WIDTH] : ping_storage_data_525 ^ i_input_data[479 % IN_WIDTH];
                485 / IN_WIDTH: ping_storage_data_525 <= (fillup_transition == 1'b1) ? i_input_data[485 % IN_WIDTH] : ping_storage_data_525 ^ i_input_data[485 % IN_WIDTH];
                731 / IN_WIDTH: ping_storage_data_525 <= (fillup_transition == 1'b1) ? i_input_data[731 % IN_WIDTH] : ping_storage_data_525 ^ i_input_data[731 % IN_WIDTH];
                1118 / IN_WIDTH: ping_storage_data_525 <= (fillup_transition == 1'b1) ? i_input_data[1118 % IN_WIDTH] : ping_storage_data_525 ^ i_input_data[1118 % IN_WIDTH];
                default: ping_storage_data_525 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_525;
                endcase
            end else begin
                case (input_count)
                479 / IN_WIDTH: pong_storage_data_525 <= (fillup_transition == 1'b1) ? i_input_data[479 % IN_WIDTH] : pong_storage_data_525 ^ i_input_data[479 % IN_WIDTH];
                485 / IN_WIDTH: pong_storage_data_525 <= (fillup_transition == 1'b1) ? i_input_data[485 % IN_WIDTH] : pong_storage_data_525 ^ i_input_data[485 % IN_WIDTH];
                731 / IN_WIDTH: pong_storage_data_525 <= (fillup_transition == 1'b1) ? i_input_data[731 % IN_WIDTH] : pong_storage_data_525 ^ i_input_data[731 % IN_WIDTH];
                1118 / IN_WIDTH: pong_storage_data_525 <= (fillup_transition == 1'b1) ? i_input_data[1118 % IN_WIDTH] : pong_storage_data_525 ^ i_input_data[1118 % IN_WIDTH];
                default: pong_storage_data_525 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_525;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_525 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_525;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_525 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_525;
            end
        end
    end
end

logic ping_storage_data_526;
logic pong_storage_data_526;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_526 <= 1'b0;
        pong_storage_data_526 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                384 / IN_WIDTH: ping_storage_data_526 <= (fillup_transition == 1'b1) ? i_input_data[384 % IN_WIDTH] : ping_storage_data_526 ^ i_input_data[384 % IN_WIDTH];
                486 / IN_WIDTH: ping_storage_data_526 <= (fillup_transition == 1'b1) ? i_input_data[486 % IN_WIDTH] : ping_storage_data_526 ^ i_input_data[486 % IN_WIDTH];
                732 / IN_WIDTH: ping_storage_data_526 <= (fillup_transition == 1'b1) ? i_input_data[732 % IN_WIDTH] : ping_storage_data_526 ^ i_input_data[732 % IN_WIDTH];
                1119 / IN_WIDTH: ping_storage_data_526 <= (fillup_transition == 1'b1) ? i_input_data[1119 % IN_WIDTH] : ping_storage_data_526 ^ i_input_data[1119 % IN_WIDTH];
                default: ping_storage_data_526 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_526;
                endcase
            end else begin
                case (input_count)
                384 / IN_WIDTH: pong_storage_data_526 <= (fillup_transition == 1'b1) ? i_input_data[384 % IN_WIDTH] : pong_storage_data_526 ^ i_input_data[384 % IN_WIDTH];
                486 / IN_WIDTH: pong_storage_data_526 <= (fillup_transition == 1'b1) ? i_input_data[486 % IN_WIDTH] : pong_storage_data_526 ^ i_input_data[486 % IN_WIDTH];
                732 / IN_WIDTH: pong_storage_data_526 <= (fillup_transition == 1'b1) ? i_input_data[732 % IN_WIDTH] : pong_storage_data_526 ^ i_input_data[732 % IN_WIDTH];
                1119 / IN_WIDTH: pong_storage_data_526 <= (fillup_transition == 1'b1) ? i_input_data[1119 % IN_WIDTH] : pong_storage_data_526 ^ i_input_data[1119 % IN_WIDTH];
                default: pong_storage_data_526 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_526;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_526 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_526;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_526 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_526;
            end
        end
    end
end

logic ping_storage_data_527;
logic pong_storage_data_527;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_527 <= 1'b0;
        pong_storage_data_527 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                385 / IN_WIDTH: ping_storage_data_527 <= (fillup_transition == 1'b1) ? i_input_data[385 % IN_WIDTH] : ping_storage_data_527 ^ i_input_data[385 % IN_WIDTH];
                487 / IN_WIDTH: ping_storage_data_527 <= (fillup_transition == 1'b1) ? i_input_data[487 % IN_WIDTH] : ping_storage_data_527 ^ i_input_data[487 % IN_WIDTH];
                733 / IN_WIDTH: ping_storage_data_527 <= (fillup_transition == 1'b1) ? i_input_data[733 % IN_WIDTH] : ping_storage_data_527 ^ i_input_data[733 % IN_WIDTH];
                1120 / IN_WIDTH: ping_storage_data_527 <= (fillup_transition == 1'b1) ? i_input_data[1120 % IN_WIDTH] : ping_storage_data_527 ^ i_input_data[1120 % IN_WIDTH];
                default: ping_storage_data_527 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_527;
                endcase
            end else begin
                case (input_count)
                385 / IN_WIDTH: pong_storage_data_527 <= (fillup_transition == 1'b1) ? i_input_data[385 % IN_WIDTH] : pong_storage_data_527 ^ i_input_data[385 % IN_WIDTH];
                487 / IN_WIDTH: pong_storage_data_527 <= (fillup_transition == 1'b1) ? i_input_data[487 % IN_WIDTH] : pong_storage_data_527 ^ i_input_data[487 % IN_WIDTH];
                733 / IN_WIDTH: pong_storage_data_527 <= (fillup_transition == 1'b1) ? i_input_data[733 % IN_WIDTH] : pong_storage_data_527 ^ i_input_data[733 % IN_WIDTH];
                1120 / IN_WIDTH: pong_storage_data_527 <= (fillup_transition == 1'b1) ? i_input_data[1120 % IN_WIDTH] : pong_storage_data_527 ^ i_input_data[1120 % IN_WIDTH];
                default: pong_storage_data_527 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_527;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_527 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_527;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_527 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_527;
            end
        end
    end
end

logic ping_storage_data_528;
logic pong_storage_data_528;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_528 <= 1'b0;
        pong_storage_data_528 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                386 / IN_WIDTH: ping_storage_data_528 <= (fillup_transition == 1'b1) ? i_input_data[386 % IN_WIDTH] : ping_storage_data_528 ^ i_input_data[386 % IN_WIDTH];
                488 / IN_WIDTH: ping_storage_data_528 <= (fillup_transition == 1'b1) ? i_input_data[488 % IN_WIDTH] : ping_storage_data_528 ^ i_input_data[488 % IN_WIDTH];
                734 / IN_WIDTH: ping_storage_data_528 <= (fillup_transition == 1'b1) ? i_input_data[734 % IN_WIDTH] : ping_storage_data_528 ^ i_input_data[734 % IN_WIDTH];
                1121 / IN_WIDTH: ping_storage_data_528 <= (fillup_transition == 1'b1) ? i_input_data[1121 % IN_WIDTH] : ping_storage_data_528 ^ i_input_data[1121 % IN_WIDTH];
                default: ping_storage_data_528 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_528;
                endcase
            end else begin
                case (input_count)
                386 / IN_WIDTH: pong_storage_data_528 <= (fillup_transition == 1'b1) ? i_input_data[386 % IN_WIDTH] : pong_storage_data_528 ^ i_input_data[386 % IN_WIDTH];
                488 / IN_WIDTH: pong_storage_data_528 <= (fillup_transition == 1'b1) ? i_input_data[488 % IN_WIDTH] : pong_storage_data_528 ^ i_input_data[488 % IN_WIDTH];
                734 / IN_WIDTH: pong_storage_data_528 <= (fillup_transition == 1'b1) ? i_input_data[734 % IN_WIDTH] : pong_storage_data_528 ^ i_input_data[734 % IN_WIDTH];
                1121 / IN_WIDTH: pong_storage_data_528 <= (fillup_transition == 1'b1) ? i_input_data[1121 % IN_WIDTH] : pong_storage_data_528 ^ i_input_data[1121 % IN_WIDTH];
                default: pong_storage_data_528 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_528;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_528 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_528;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_528 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_528;
            end
        end
    end
end

logic ping_storage_data_529;
logic pong_storage_data_529;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_529 <= 1'b0;
        pong_storage_data_529 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                387 / IN_WIDTH: ping_storage_data_529 <= (fillup_transition == 1'b1) ? i_input_data[387 % IN_WIDTH] : ping_storage_data_529 ^ i_input_data[387 % IN_WIDTH];
                489 / IN_WIDTH: ping_storage_data_529 <= (fillup_transition == 1'b1) ? i_input_data[489 % IN_WIDTH] : ping_storage_data_529 ^ i_input_data[489 % IN_WIDTH];
                735 / IN_WIDTH: ping_storage_data_529 <= (fillup_transition == 1'b1) ? i_input_data[735 % IN_WIDTH] : ping_storage_data_529 ^ i_input_data[735 % IN_WIDTH];
                1122 / IN_WIDTH: ping_storage_data_529 <= (fillup_transition == 1'b1) ? i_input_data[1122 % IN_WIDTH] : ping_storage_data_529 ^ i_input_data[1122 % IN_WIDTH];
                default: ping_storage_data_529 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_529;
                endcase
            end else begin
                case (input_count)
                387 / IN_WIDTH: pong_storage_data_529 <= (fillup_transition == 1'b1) ? i_input_data[387 % IN_WIDTH] : pong_storage_data_529 ^ i_input_data[387 % IN_WIDTH];
                489 / IN_WIDTH: pong_storage_data_529 <= (fillup_transition == 1'b1) ? i_input_data[489 % IN_WIDTH] : pong_storage_data_529 ^ i_input_data[489 % IN_WIDTH];
                735 / IN_WIDTH: pong_storage_data_529 <= (fillup_transition == 1'b1) ? i_input_data[735 % IN_WIDTH] : pong_storage_data_529 ^ i_input_data[735 % IN_WIDTH];
                1122 / IN_WIDTH: pong_storage_data_529 <= (fillup_transition == 1'b1) ? i_input_data[1122 % IN_WIDTH] : pong_storage_data_529 ^ i_input_data[1122 % IN_WIDTH];
                default: pong_storage_data_529 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_529;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_529 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_529;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_529 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_529;
            end
        end
    end
end

logic ping_storage_data_530;
logic pong_storage_data_530;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_530 <= 1'b0;
        pong_storage_data_530 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                388 / IN_WIDTH: ping_storage_data_530 <= (fillup_transition == 1'b1) ? i_input_data[388 % IN_WIDTH] : ping_storage_data_530 ^ i_input_data[388 % IN_WIDTH];
                490 / IN_WIDTH: ping_storage_data_530 <= (fillup_transition == 1'b1) ? i_input_data[490 % IN_WIDTH] : ping_storage_data_530 ^ i_input_data[490 % IN_WIDTH];
                736 / IN_WIDTH: ping_storage_data_530 <= (fillup_transition == 1'b1) ? i_input_data[736 % IN_WIDTH] : ping_storage_data_530 ^ i_input_data[736 % IN_WIDTH];
                1123 / IN_WIDTH: ping_storage_data_530 <= (fillup_transition == 1'b1) ? i_input_data[1123 % IN_WIDTH] : ping_storage_data_530 ^ i_input_data[1123 % IN_WIDTH];
                default: ping_storage_data_530 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_530;
                endcase
            end else begin
                case (input_count)
                388 / IN_WIDTH: pong_storage_data_530 <= (fillup_transition == 1'b1) ? i_input_data[388 % IN_WIDTH] : pong_storage_data_530 ^ i_input_data[388 % IN_WIDTH];
                490 / IN_WIDTH: pong_storage_data_530 <= (fillup_transition == 1'b1) ? i_input_data[490 % IN_WIDTH] : pong_storage_data_530 ^ i_input_data[490 % IN_WIDTH];
                736 / IN_WIDTH: pong_storage_data_530 <= (fillup_transition == 1'b1) ? i_input_data[736 % IN_WIDTH] : pong_storage_data_530 ^ i_input_data[736 % IN_WIDTH];
                1123 / IN_WIDTH: pong_storage_data_530 <= (fillup_transition == 1'b1) ? i_input_data[1123 % IN_WIDTH] : pong_storage_data_530 ^ i_input_data[1123 % IN_WIDTH];
                default: pong_storage_data_530 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_530;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_530 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_530;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_530 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_530;
            end
        end
    end
end

logic ping_storage_data_531;
logic pong_storage_data_531;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_531 <= 1'b0;
        pong_storage_data_531 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                389 / IN_WIDTH: ping_storage_data_531 <= (fillup_transition == 1'b1) ? i_input_data[389 % IN_WIDTH] : ping_storage_data_531 ^ i_input_data[389 % IN_WIDTH];
                491 / IN_WIDTH: ping_storage_data_531 <= (fillup_transition == 1'b1) ? i_input_data[491 % IN_WIDTH] : ping_storage_data_531 ^ i_input_data[491 % IN_WIDTH];
                737 / IN_WIDTH: ping_storage_data_531 <= (fillup_transition == 1'b1) ? i_input_data[737 % IN_WIDTH] : ping_storage_data_531 ^ i_input_data[737 % IN_WIDTH];
                1124 / IN_WIDTH: ping_storage_data_531 <= (fillup_transition == 1'b1) ? i_input_data[1124 % IN_WIDTH] : ping_storage_data_531 ^ i_input_data[1124 % IN_WIDTH];
                default: ping_storage_data_531 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_531;
                endcase
            end else begin
                case (input_count)
                389 / IN_WIDTH: pong_storage_data_531 <= (fillup_transition == 1'b1) ? i_input_data[389 % IN_WIDTH] : pong_storage_data_531 ^ i_input_data[389 % IN_WIDTH];
                491 / IN_WIDTH: pong_storage_data_531 <= (fillup_transition == 1'b1) ? i_input_data[491 % IN_WIDTH] : pong_storage_data_531 ^ i_input_data[491 % IN_WIDTH];
                737 / IN_WIDTH: pong_storage_data_531 <= (fillup_transition == 1'b1) ? i_input_data[737 % IN_WIDTH] : pong_storage_data_531 ^ i_input_data[737 % IN_WIDTH];
                1124 / IN_WIDTH: pong_storage_data_531 <= (fillup_transition == 1'b1) ? i_input_data[1124 % IN_WIDTH] : pong_storage_data_531 ^ i_input_data[1124 % IN_WIDTH];
                default: pong_storage_data_531 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_531;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_531 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_531;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_531 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_531;
            end
        end
    end
end

logic ping_storage_data_532;
logic pong_storage_data_532;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_532 <= 1'b0;
        pong_storage_data_532 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                390 / IN_WIDTH: ping_storage_data_532 <= (fillup_transition == 1'b1) ? i_input_data[390 % IN_WIDTH] : ping_storage_data_532 ^ i_input_data[390 % IN_WIDTH];
                492 / IN_WIDTH: ping_storage_data_532 <= (fillup_transition == 1'b1) ? i_input_data[492 % IN_WIDTH] : ping_storage_data_532 ^ i_input_data[492 % IN_WIDTH];
                738 / IN_WIDTH: ping_storage_data_532 <= (fillup_transition == 1'b1) ? i_input_data[738 % IN_WIDTH] : ping_storage_data_532 ^ i_input_data[738 % IN_WIDTH];
                1125 / IN_WIDTH: ping_storage_data_532 <= (fillup_transition == 1'b1) ? i_input_data[1125 % IN_WIDTH] : ping_storage_data_532 ^ i_input_data[1125 % IN_WIDTH];
                default: ping_storage_data_532 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_532;
                endcase
            end else begin
                case (input_count)
                390 / IN_WIDTH: pong_storage_data_532 <= (fillup_transition == 1'b1) ? i_input_data[390 % IN_WIDTH] : pong_storage_data_532 ^ i_input_data[390 % IN_WIDTH];
                492 / IN_WIDTH: pong_storage_data_532 <= (fillup_transition == 1'b1) ? i_input_data[492 % IN_WIDTH] : pong_storage_data_532 ^ i_input_data[492 % IN_WIDTH];
                738 / IN_WIDTH: pong_storage_data_532 <= (fillup_transition == 1'b1) ? i_input_data[738 % IN_WIDTH] : pong_storage_data_532 ^ i_input_data[738 % IN_WIDTH];
                1125 / IN_WIDTH: pong_storage_data_532 <= (fillup_transition == 1'b1) ? i_input_data[1125 % IN_WIDTH] : pong_storage_data_532 ^ i_input_data[1125 % IN_WIDTH];
                default: pong_storage_data_532 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_532;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_532 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_532;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_532 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_532;
            end
        end
    end
end

logic ping_storage_data_533;
logic pong_storage_data_533;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_533 <= 1'b0;
        pong_storage_data_533 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                391 / IN_WIDTH: ping_storage_data_533 <= (fillup_transition == 1'b1) ? i_input_data[391 % IN_WIDTH] : ping_storage_data_533 ^ i_input_data[391 % IN_WIDTH];
                493 / IN_WIDTH: ping_storage_data_533 <= (fillup_transition == 1'b1) ? i_input_data[493 % IN_WIDTH] : ping_storage_data_533 ^ i_input_data[493 % IN_WIDTH];
                739 / IN_WIDTH: ping_storage_data_533 <= (fillup_transition == 1'b1) ? i_input_data[739 % IN_WIDTH] : ping_storage_data_533 ^ i_input_data[739 % IN_WIDTH];
                1126 / IN_WIDTH: ping_storage_data_533 <= (fillup_transition == 1'b1) ? i_input_data[1126 % IN_WIDTH] : ping_storage_data_533 ^ i_input_data[1126 % IN_WIDTH];
                default: ping_storage_data_533 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_533;
                endcase
            end else begin
                case (input_count)
                391 / IN_WIDTH: pong_storage_data_533 <= (fillup_transition == 1'b1) ? i_input_data[391 % IN_WIDTH] : pong_storage_data_533 ^ i_input_data[391 % IN_WIDTH];
                493 / IN_WIDTH: pong_storage_data_533 <= (fillup_transition == 1'b1) ? i_input_data[493 % IN_WIDTH] : pong_storage_data_533 ^ i_input_data[493 % IN_WIDTH];
                739 / IN_WIDTH: pong_storage_data_533 <= (fillup_transition == 1'b1) ? i_input_data[739 % IN_WIDTH] : pong_storage_data_533 ^ i_input_data[739 % IN_WIDTH];
                1126 / IN_WIDTH: pong_storage_data_533 <= (fillup_transition == 1'b1) ? i_input_data[1126 % IN_WIDTH] : pong_storage_data_533 ^ i_input_data[1126 % IN_WIDTH];
                default: pong_storage_data_533 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_533;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_533 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_533;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_533 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_533;
            end
        end
    end
end

logic ping_storage_data_534;
logic pong_storage_data_534;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_534 <= 1'b0;
        pong_storage_data_534 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                392 / IN_WIDTH: ping_storage_data_534 <= (fillup_transition == 1'b1) ? i_input_data[392 % IN_WIDTH] : ping_storage_data_534 ^ i_input_data[392 % IN_WIDTH];
                494 / IN_WIDTH: ping_storage_data_534 <= (fillup_transition == 1'b1) ? i_input_data[494 % IN_WIDTH] : ping_storage_data_534 ^ i_input_data[494 % IN_WIDTH];
                740 / IN_WIDTH: ping_storage_data_534 <= (fillup_transition == 1'b1) ? i_input_data[740 % IN_WIDTH] : ping_storage_data_534 ^ i_input_data[740 % IN_WIDTH];
                1127 / IN_WIDTH: ping_storage_data_534 <= (fillup_transition == 1'b1) ? i_input_data[1127 % IN_WIDTH] : ping_storage_data_534 ^ i_input_data[1127 % IN_WIDTH];
                default: ping_storage_data_534 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_534;
                endcase
            end else begin
                case (input_count)
                392 / IN_WIDTH: pong_storage_data_534 <= (fillup_transition == 1'b1) ? i_input_data[392 % IN_WIDTH] : pong_storage_data_534 ^ i_input_data[392 % IN_WIDTH];
                494 / IN_WIDTH: pong_storage_data_534 <= (fillup_transition == 1'b1) ? i_input_data[494 % IN_WIDTH] : pong_storage_data_534 ^ i_input_data[494 % IN_WIDTH];
                740 / IN_WIDTH: pong_storage_data_534 <= (fillup_transition == 1'b1) ? i_input_data[740 % IN_WIDTH] : pong_storage_data_534 ^ i_input_data[740 % IN_WIDTH];
                1127 / IN_WIDTH: pong_storage_data_534 <= (fillup_transition == 1'b1) ? i_input_data[1127 % IN_WIDTH] : pong_storage_data_534 ^ i_input_data[1127 % IN_WIDTH];
                default: pong_storage_data_534 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_534;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_534 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_534;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_534 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_534;
            end
        end
    end
end

logic ping_storage_data_535;
logic pong_storage_data_535;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_535 <= 1'b0;
        pong_storage_data_535 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                393 / IN_WIDTH: ping_storage_data_535 <= (fillup_transition == 1'b1) ? i_input_data[393 % IN_WIDTH] : ping_storage_data_535 ^ i_input_data[393 % IN_WIDTH];
                495 / IN_WIDTH: ping_storage_data_535 <= (fillup_transition == 1'b1) ? i_input_data[495 % IN_WIDTH] : ping_storage_data_535 ^ i_input_data[495 % IN_WIDTH];
                741 / IN_WIDTH: ping_storage_data_535 <= (fillup_transition == 1'b1) ? i_input_data[741 % IN_WIDTH] : ping_storage_data_535 ^ i_input_data[741 % IN_WIDTH];
                1128 / IN_WIDTH: ping_storage_data_535 <= (fillup_transition == 1'b1) ? i_input_data[1128 % IN_WIDTH] : ping_storage_data_535 ^ i_input_data[1128 % IN_WIDTH];
                default: ping_storage_data_535 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_535;
                endcase
            end else begin
                case (input_count)
                393 / IN_WIDTH: pong_storage_data_535 <= (fillup_transition == 1'b1) ? i_input_data[393 % IN_WIDTH] : pong_storage_data_535 ^ i_input_data[393 % IN_WIDTH];
                495 / IN_WIDTH: pong_storage_data_535 <= (fillup_transition == 1'b1) ? i_input_data[495 % IN_WIDTH] : pong_storage_data_535 ^ i_input_data[495 % IN_WIDTH];
                741 / IN_WIDTH: pong_storage_data_535 <= (fillup_transition == 1'b1) ? i_input_data[741 % IN_WIDTH] : pong_storage_data_535 ^ i_input_data[741 % IN_WIDTH];
                1128 / IN_WIDTH: pong_storage_data_535 <= (fillup_transition == 1'b1) ? i_input_data[1128 % IN_WIDTH] : pong_storage_data_535 ^ i_input_data[1128 % IN_WIDTH];
                default: pong_storage_data_535 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_535;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_535 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_535;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_535 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_535;
            end
        end
    end
end

logic ping_storage_data_536;
logic pong_storage_data_536;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_536 <= 1'b0;
        pong_storage_data_536 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                394 / IN_WIDTH: ping_storage_data_536 <= (fillup_transition == 1'b1) ? i_input_data[394 % IN_WIDTH] : ping_storage_data_536 ^ i_input_data[394 % IN_WIDTH];
                496 / IN_WIDTH: ping_storage_data_536 <= (fillup_transition == 1'b1) ? i_input_data[496 % IN_WIDTH] : ping_storage_data_536 ^ i_input_data[496 % IN_WIDTH];
                742 / IN_WIDTH: ping_storage_data_536 <= (fillup_transition == 1'b1) ? i_input_data[742 % IN_WIDTH] : ping_storage_data_536 ^ i_input_data[742 % IN_WIDTH];
                1129 / IN_WIDTH: ping_storage_data_536 <= (fillup_transition == 1'b1) ? i_input_data[1129 % IN_WIDTH] : ping_storage_data_536 ^ i_input_data[1129 % IN_WIDTH];
                default: ping_storage_data_536 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_536;
                endcase
            end else begin
                case (input_count)
                394 / IN_WIDTH: pong_storage_data_536 <= (fillup_transition == 1'b1) ? i_input_data[394 % IN_WIDTH] : pong_storage_data_536 ^ i_input_data[394 % IN_WIDTH];
                496 / IN_WIDTH: pong_storage_data_536 <= (fillup_transition == 1'b1) ? i_input_data[496 % IN_WIDTH] : pong_storage_data_536 ^ i_input_data[496 % IN_WIDTH];
                742 / IN_WIDTH: pong_storage_data_536 <= (fillup_transition == 1'b1) ? i_input_data[742 % IN_WIDTH] : pong_storage_data_536 ^ i_input_data[742 % IN_WIDTH];
                1129 / IN_WIDTH: pong_storage_data_536 <= (fillup_transition == 1'b1) ? i_input_data[1129 % IN_WIDTH] : pong_storage_data_536 ^ i_input_data[1129 % IN_WIDTH];
                default: pong_storage_data_536 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_536;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_536 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_536;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_536 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_536;
            end
        end
    end
end

logic ping_storage_data_537;
logic pong_storage_data_537;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_537 <= 1'b0;
        pong_storage_data_537 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                395 / IN_WIDTH: ping_storage_data_537 <= (fillup_transition == 1'b1) ? i_input_data[395 % IN_WIDTH] : ping_storage_data_537 ^ i_input_data[395 % IN_WIDTH];
                497 / IN_WIDTH: ping_storage_data_537 <= (fillup_transition == 1'b1) ? i_input_data[497 % IN_WIDTH] : ping_storage_data_537 ^ i_input_data[497 % IN_WIDTH];
                743 / IN_WIDTH: ping_storage_data_537 <= (fillup_transition == 1'b1) ? i_input_data[743 % IN_WIDTH] : ping_storage_data_537 ^ i_input_data[743 % IN_WIDTH];
                1130 / IN_WIDTH: ping_storage_data_537 <= (fillup_transition == 1'b1) ? i_input_data[1130 % IN_WIDTH] : ping_storage_data_537 ^ i_input_data[1130 % IN_WIDTH];
                default: ping_storage_data_537 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_537;
                endcase
            end else begin
                case (input_count)
                395 / IN_WIDTH: pong_storage_data_537 <= (fillup_transition == 1'b1) ? i_input_data[395 % IN_WIDTH] : pong_storage_data_537 ^ i_input_data[395 % IN_WIDTH];
                497 / IN_WIDTH: pong_storage_data_537 <= (fillup_transition == 1'b1) ? i_input_data[497 % IN_WIDTH] : pong_storage_data_537 ^ i_input_data[497 % IN_WIDTH];
                743 / IN_WIDTH: pong_storage_data_537 <= (fillup_transition == 1'b1) ? i_input_data[743 % IN_WIDTH] : pong_storage_data_537 ^ i_input_data[743 % IN_WIDTH];
                1130 / IN_WIDTH: pong_storage_data_537 <= (fillup_transition == 1'b1) ? i_input_data[1130 % IN_WIDTH] : pong_storage_data_537 ^ i_input_data[1130 % IN_WIDTH];
                default: pong_storage_data_537 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_537;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_537 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_537;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_537 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_537;
            end
        end
    end
end

logic ping_storage_data_538;
logic pong_storage_data_538;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_538 <= 1'b0;
        pong_storage_data_538 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                396 / IN_WIDTH: ping_storage_data_538 <= (fillup_transition == 1'b1) ? i_input_data[396 % IN_WIDTH] : ping_storage_data_538 ^ i_input_data[396 % IN_WIDTH];
                498 / IN_WIDTH: ping_storage_data_538 <= (fillup_transition == 1'b1) ? i_input_data[498 % IN_WIDTH] : ping_storage_data_538 ^ i_input_data[498 % IN_WIDTH];
                744 / IN_WIDTH: ping_storage_data_538 <= (fillup_transition == 1'b1) ? i_input_data[744 % IN_WIDTH] : ping_storage_data_538 ^ i_input_data[744 % IN_WIDTH];
                1131 / IN_WIDTH: ping_storage_data_538 <= (fillup_transition == 1'b1) ? i_input_data[1131 % IN_WIDTH] : ping_storage_data_538 ^ i_input_data[1131 % IN_WIDTH];
                default: ping_storage_data_538 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_538;
                endcase
            end else begin
                case (input_count)
                396 / IN_WIDTH: pong_storage_data_538 <= (fillup_transition == 1'b1) ? i_input_data[396 % IN_WIDTH] : pong_storage_data_538 ^ i_input_data[396 % IN_WIDTH];
                498 / IN_WIDTH: pong_storage_data_538 <= (fillup_transition == 1'b1) ? i_input_data[498 % IN_WIDTH] : pong_storage_data_538 ^ i_input_data[498 % IN_WIDTH];
                744 / IN_WIDTH: pong_storage_data_538 <= (fillup_transition == 1'b1) ? i_input_data[744 % IN_WIDTH] : pong_storage_data_538 ^ i_input_data[744 % IN_WIDTH];
                1131 / IN_WIDTH: pong_storage_data_538 <= (fillup_transition == 1'b1) ? i_input_data[1131 % IN_WIDTH] : pong_storage_data_538 ^ i_input_data[1131 % IN_WIDTH];
                default: pong_storage_data_538 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_538;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_538 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_538;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_538 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_538;
            end
        end
    end
end

logic ping_storage_data_539;
logic pong_storage_data_539;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_539 <= 1'b0;
        pong_storage_data_539 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                397 / IN_WIDTH: ping_storage_data_539 <= (fillup_transition == 1'b1) ? i_input_data[397 % IN_WIDTH] : ping_storage_data_539 ^ i_input_data[397 % IN_WIDTH];
                499 / IN_WIDTH: ping_storage_data_539 <= (fillup_transition == 1'b1) ? i_input_data[499 % IN_WIDTH] : ping_storage_data_539 ^ i_input_data[499 % IN_WIDTH];
                745 / IN_WIDTH: ping_storage_data_539 <= (fillup_transition == 1'b1) ? i_input_data[745 % IN_WIDTH] : ping_storage_data_539 ^ i_input_data[745 % IN_WIDTH];
                1132 / IN_WIDTH: ping_storage_data_539 <= (fillup_transition == 1'b1) ? i_input_data[1132 % IN_WIDTH] : ping_storage_data_539 ^ i_input_data[1132 % IN_WIDTH];
                default: ping_storage_data_539 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_539;
                endcase
            end else begin
                case (input_count)
                397 / IN_WIDTH: pong_storage_data_539 <= (fillup_transition == 1'b1) ? i_input_data[397 % IN_WIDTH] : pong_storage_data_539 ^ i_input_data[397 % IN_WIDTH];
                499 / IN_WIDTH: pong_storage_data_539 <= (fillup_transition == 1'b1) ? i_input_data[499 % IN_WIDTH] : pong_storage_data_539 ^ i_input_data[499 % IN_WIDTH];
                745 / IN_WIDTH: pong_storage_data_539 <= (fillup_transition == 1'b1) ? i_input_data[745 % IN_WIDTH] : pong_storage_data_539 ^ i_input_data[745 % IN_WIDTH];
                1132 / IN_WIDTH: pong_storage_data_539 <= (fillup_transition == 1'b1) ? i_input_data[1132 % IN_WIDTH] : pong_storage_data_539 ^ i_input_data[1132 % IN_WIDTH];
                default: pong_storage_data_539 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_539;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_539 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_539;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_539 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_539;
            end
        end
    end
end

logic ping_storage_data_540;
logic pong_storage_data_540;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_540 <= 1'b0;
        pong_storage_data_540 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                398 / IN_WIDTH: ping_storage_data_540 <= (fillup_transition == 1'b1) ? i_input_data[398 % IN_WIDTH] : ping_storage_data_540 ^ i_input_data[398 % IN_WIDTH];
                500 / IN_WIDTH: ping_storage_data_540 <= (fillup_transition == 1'b1) ? i_input_data[500 % IN_WIDTH] : ping_storage_data_540 ^ i_input_data[500 % IN_WIDTH];
                746 / IN_WIDTH: ping_storage_data_540 <= (fillup_transition == 1'b1) ? i_input_data[746 % IN_WIDTH] : ping_storage_data_540 ^ i_input_data[746 % IN_WIDTH];
                1133 / IN_WIDTH: ping_storage_data_540 <= (fillup_transition == 1'b1) ? i_input_data[1133 % IN_WIDTH] : ping_storage_data_540 ^ i_input_data[1133 % IN_WIDTH];
                default: ping_storage_data_540 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_540;
                endcase
            end else begin
                case (input_count)
                398 / IN_WIDTH: pong_storage_data_540 <= (fillup_transition == 1'b1) ? i_input_data[398 % IN_WIDTH] : pong_storage_data_540 ^ i_input_data[398 % IN_WIDTH];
                500 / IN_WIDTH: pong_storage_data_540 <= (fillup_transition == 1'b1) ? i_input_data[500 % IN_WIDTH] : pong_storage_data_540 ^ i_input_data[500 % IN_WIDTH];
                746 / IN_WIDTH: pong_storage_data_540 <= (fillup_transition == 1'b1) ? i_input_data[746 % IN_WIDTH] : pong_storage_data_540 ^ i_input_data[746 % IN_WIDTH];
                1133 / IN_WIDTH: pong_storage_data_540 <= (fillup_transition == 1'b1) ? i_input_data[1133 % IN_WIDTH] : pong_storage_data_540 ^ i_input_data[1133 % IN_WIDTH];
                default: pong_storage_data_540 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_540;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_540 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_540;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_540 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_540;
            end
        end
    end
end

logic ping_storage_data_541;
logic pong_storage_data_541;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_541 <= 1'b0;
        pong_storage_data_541 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                399 / IN_WIDTH: ping_storage_data_541 <= (fillup_transition == 1'b1) ? i_input_data[399 % IN_WIDTH] : ping_storage_data_541 ^ i_input_data[399 % IN_WIDTH];
                501 / IN_WIDTH: ping_storage_data_541 <= (fillup_transition == 1'b1) ? i_input_data[501 % IN_WIDTH] : ping_storage_data_541 ^ i_input_data[501 % IN_WIDTH];
                747 / IN_WIDTH: ping_storage_data_541 <= (fillup_transition == 1'b1) ? i_input_data[747 % IN_WIDTH] : ping_storage_data_541 ^ i_input_data[747 % IN_WIDTH];
                1134 / IN_WIDTH: ping_storage_data_541 <= (fillup_transition == 1'b1) ? i_input_data[1134 % IN_WIDTH] : ping_storage_data_541 ^ i_input_data[1134 % IN_WIDTH];
                default: ping_storage_data_541 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_541;
                endcase
            end else begin
                case (input_count)
                399 / IN_WIDTH: pong_storage_data_541 <= (fillup_transition == 1'b1) ? i_input_data[399 % IN_WIDTH] : pong_storage_data_541 ^ i_input_data[399 % IN_WIDTH];
                501 / IN_WIDTH: pong_storage_data_541 <= (fillup_transition == 1'b1) ? i_input_data[501 % IN_WIDTH] : pong_storage_data_541 ^ i_input_data[501 % IN_WIDTH];
                747 / IN_WIDTH: pong_storage_data_541 <= (fillup_transition == 1'b1) ? i_input_data[747 % IN_WIDTH] : pong_storage_data_541 ^ i_input_data[747 % IN_WIDTH];
                1134 / IN_WIDTH: pong_storage_data_541 <= (fillup_transition == 1'b1) ? i_input_data[1134 % IN_WIDTH] : pong_storage_data_541 ^ i_input_data[1134 % IN_WIDTH];
                default: pong_storage_data_541 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_541;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_541 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_541;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_541 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_541;
            end
        end
    end
end

logic ping_storage_data_542;
logic pong_storage_data_542;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_542 <= 1'b0;
        pong_storage_data_542 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                400 / IN_WIDTH: ping_storage_data_542 <= (fillup_transition == 1'b1) ? i_input_data[400 % IN_WIDTH] : ping_storage_data_542 ^ i_input_data[400 % IN_WIDTH];
                502 / IN_WIDTH: ping_storage_data_542 <= (fillup_transition == 1'b1) ? i_input_data[502 % IN_WIDTH] : ping_storage_data_542 ^ i_input_data[502 % IN_WIDTH];
                748 / IN_WIDTH: ping_storage_data_542 <= (fillup_transition == 1'b1) ? i_input_data[748 % IN_WIDTH] : ping_storage_data_542 ^ i_input_data[748 % IN_WIDTH];
                1135 / IN_WIDTH: ping_storage_data_542 <= (fillup_transition == 1'b1) ? i_input_data[1135 % IN_WIDTH] : ping_storage_data_542 ^ i_input_data[1135 % IN_WIDTH];
                default: ping_storage_data_542 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_542;
                endcase
            end else begin
                case (input_count)
                400 / IN_WIDTH: pong_storage_data_542 <= (fillup_transition == 1'b1) ? i_input_data[400 % IN_WIDTH] : pong_storage_data_542 ^ i_input_data[400 % IN_WIDTH];
                502 / IN_WIDTH: pong_storage_data_542 <= (fillup_transition == 1'b1) ? i_input_data[502 % IN_WIDTH] : pong_storage_data_542 ^ i_input_data[502 % IN_WIDTH];
                748 / IN_WIDTH: pong_storage_data_542 <= (fillup_transition == 1'b1) ? i_input_data[748 % IN_WIDTH] : pong_storage_data_542 ^ i_input_data[748 % IN_WIDTH];
                1135 / IN_WIDTH: pong_storage_data_542 <= (fillup_transition == 1'b1) ? i_input_data[1135 % IN_WIDTH] : pong_storage_data_542 ^ i_input_data[1135 % IN_WIDTH];
                default: pong_storage_data_542 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_542;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_542 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_542;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_542 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_542;
            end
        end
    end
end

logic ping_storage_data_543;
logic pong_storage_data_543;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_543 <= 1'b0;
        pong_storage_data_543 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                401 / IN_WIDTH: ping_storage_data_543 <= (fillup_transition == 1'b1) ? i_input_data[401 % IN_WIDTH] : ping_storage_data_543 ^ i_input_data[401 % IN_WIDTH];
                503 / IN_WIDTH: ping_storage_data_543 <= (fillup_transition == 1'b1) ? i_input_data[503 % IN_WIDTH] : ping_storage_data_543 ^ i_input_data[503 % IN_WIDTH];
                749 / IN_WIDTH: ping_storage_data_543 <= (fillup_transition == 1'b1) ? i_input_data[749 % IN_WIDTH] : ping_storage_data_543 ^ i_input_data[749 % IN_WIDTH];
                1136 / IN_WIDTH: ping_storage_data_543 <= (fillup_transition == 1'b1) ? i_input_data[1136 % IN_WIDTH] : ping_storage_data_543 ^ i_input_data[1136 % IN_WIDTH];
                default: ping_storage_data_543 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_543;
                endcase
            end else begin
                case (input_count)
                401 / IN_WIDTH: pong_storage_data_543 <= (fillup_transition == 1'b1) ? i_input_data[401 % IN_WIDTH] : pong_storage_data_543 ^ i_input_data[401 % IN_WIDTH];
                503 / IN_WIDTH: pong_storage_data_543 <= (fillup_transition == 1'b1) ? i_input_data[503 % IN_WIDTH] : pong_storage_data_543 ^ i_input_data[503 % IN_WIDTH];
                749 / IN_WIDTH: pong_storage_data_543 <= (fillup_transition == 1'b1) ? i_input_data[749 % IN_WIDTH] : pong_storage_data_543 ^ i_input_data[749 % IN_WIDTH];
                1136 / IN_WIDTH: pong_storage_data_543 <= (fillup_transition == 1'b1) ? i_input_data[1136 % IN_WIDTH] : pong_storage_data_543 ^ i_input_data[1136 % IN_WIDTH];
                default: pong_storage_data_543 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_543;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_543 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_543;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_543 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_543;
            end
        end
    end
end

logic ping_storage_data_544;
logic pong_storage_data_544;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_544 <= 1'b0;
        pong_storage_data_544 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                402 / IN_WIDTH: ping_storage_data_544 <= (fillup_transition == 1'b1) ? i_input_data[402 % IN_WIDTH] : ping_storage_data_544 ^ i_input_data[402 % IN_WIDTH];
                504 / IN_WIDTH: ping_storage_data_544 <= (fillup_transition == 1'b1) ? i_input_data[504 % IN_WIDTH] : ping_storage_data_544 ^ i_input_data[504 % IN_WIDTH];
                750 / IN_WIDTH: ping_storage_data_544 <= (fillup_transition == 1'b1) ? i_input_data[750 % IN_WIDTH] : ping_storage_data_544 ^ i_input_data[750 % IN_WIDTH];
                1137 / IN_WIDTH: ping_storage_data_544 <= (fillup_transition == 1'b1) ? i_input_data[1137 % IN_WIDTH] : ping_storage_data_544 ^ i_input_data[1137 % IN_WIDTH];
                default: ping_storage_data_544 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_544;
                endcase
            end else begin
                case (input_count)
                402 / IN_WIDTH: pong_storage_data_544 <= (fillup_transition == 1'b1) ? i_input_data[402 % IN_WIDTH] : pong_storage_data_544 ^ i_input_data[402 % IN_WIDTH];
                504 / IN_WIDTH: pong_storage_data_544 <= (fillup_transition == 1'b1) ? i_input_data[504 % IN_WIDTH] : pong_storage_data_544 ^ i_input_data[504 % IN_WIDTH];
                750 / IN_WIDTH: pong_storage_data_544 <= (fillup_transition == 1'b1) ? i_input_data[750 % IN_WIDTH] : pong_storage_data_544 ^ i_input_data[750 % IN_WIDTH];
                1137 / IN_WIDTH: pong_storage_data_544 <= (fillup_transition == 1'b1) ? i_input_data[1137 % IN_WIDTH] : pong_storage_data_544 ^ i_input_data[1137 % IN_WIDTH];
                default: pong_storage_data_544 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_544;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_544 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_544;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_544 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_544;
            end
        end
    end
end

logic ping_storage_data_545;
logic pong_storage_data_545;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_545 <= 1'b0;
        pong_storage_data_545 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                403 / IN_WIDTH: ping_storage_data_545 <= (fillup_transition == 1'b1) ? i_input_data[403 % IN_WIDTH] : ping_storage_data_545 ^ i_input_data[403 % IN_WIDTH];
                505 / IN_WIDTH: ping_storage_data_545 <= (fillup_transition == 1'b1) ? i_input_data[505 % IN_WIDTH] : ping_storage_data_545 ^ i_input_data[505 % IN_WIDTH];
                751 / IN_WIDTH: ping_storage_data_545 <= (fillup_transition == 1'b1) ? i_input_data[751 % IN_WIDTH] : ping_storage_data_545 ^ i_input_data[751 % IN_WIDTH];
                1138 / IN_WIDTH: ping_storage_data_545 <= (fillup_transition == 1'b1) ? i_input_data[1138 % IN_WIDTH] : ping_storage_data_545 ^ i_input_data[1138 % IN_WIDTH];
                default: ping_storage_data_545 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_545;
                endcase
            end else begin
                case (input_count)
                403 / IN_WIDTH: pong_storage_data_545 <= (fillup_transition == 1'b1) ? i_input_data[403 % IN_WIDTH] : pong_storage_data_545 ^ i_input_data[403 % IN_WIDTH];
                505 / IN_WIDTH: pong_storage_data_545 <= (fillup_transition == 1'b1) ? i_input_data[505 % IN_WIDTH] : pong_storage_data_545 ^ i_input_data[505 % IN_WIDTH];
                751 / IN_WIDTH: pong_storage_data_545 <= (fillup_transition == 1'b1) ? i_input_data[751 % IN_WIDTH] : pong_storage_data_545 ^ i_input_data[751 % IN_WIDTH];
                1138 / IN_WIDTH: pong_storage_data_545 <= (fillup_transition == 1'b1) ? i_input_data[1138 % IN_WIDTH] : pong_storage_data_545 ^ i_input_data[1138 % IN_WIDTH];
                default: pong_storage_data_545 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_545;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_545 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_545;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_545 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_545;
            end
        end
    end
end

logic ping_storage_data_546;
logic pong_storage_data_546;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_546 <= 1'b0;
        pong_storage_data_546 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                404 / IN_WIDTH: ping_storage_data_546 <= (fillup_transition == 1'b1) ? i_input_data[404 % IN_WIDTH] : ping_storage_data_546 ^ i_input_data[404 % IN_WIDTH];
                506 / IN_WIDTH: ping_storage_data_546 <= (fillup_transition == 1'b1) ? i_input_data[506 % IN_WIDTH] : ping_storage_data_546 ^ i_input_data[506 % IN_WIDTH];
                752 / IN_WIDTH: ping_storage_data_546 <= (fillup_transition == 1'b1) ? i_input_data[752 % IN_WIDTH] : ping_storage_data_546 ^ i_input_data[752 % IN_WIDTH];
                1139 / IN_WIDTH: ping_storage_data_546 <= (fillup_transition == 1'b1) ? i_input_data[1139 % IN_WIDTH] : ping_storage_data_546 ^ i_input_data[1139 % IN_WIDTH];
                default: ping_storage_data_546 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_546;
                endcase
            end else begin
                case (input_count)
                404 / IN_WIDTH: pong_storage_data_546 <= (fillup_transition == 1'b1) ? i_input_data[404 % IN_WIDTH] : pong_storage_data_546 ^ i_input_data[404 % IN_WIDTH];
                506 / IN_WIDTH: pong_storage_data_546 <= (fillup_transition == 1'b1) ? i_input_data[506 % IN_WIDTH] : pong_storage_data_546 ^ i_input_data[506 % IN_WIDTH];
                752 / IN_WIDTH: pong_storage_data_546 <= (fillup_transition == 1'b1) ? i_input_data[752 % IN_WIDTH] : pong_storage_data_546 ^ i_input_data[752 % IN_WIDTH];
                1139 / IN_WIDTH: pong_storage_data_546 <= (fillup_transition == 1'b1) ? i_input_data[1139 % IN_WIDTH] : pong_storage_data_546 ^ i_input_data[1139 % IN_WIDTH];
                default: pong_storage_data_546 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_546;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_546 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_546;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_546 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_546;
            end
        end
    end
end

logic ping_storage_data_547;
logic pong_storage_data_547;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_547 <= 1'b0;
        pong_storage_data_547 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                405 / IN_WIDTH: ping_storage_data_547 <= (fillup_transition == 1'b1) ? i_input_data[405 % IN_WIDTH] : ping_storage_data_547 ^ i_input_data[405 % IN_WIDTH];
                507 / IN_WIDTH: ping_storage_data_547 <= (fillup_transition == 1'b1) ? i_input_data[507 % IN_WIDTH] : ping_storage_data_547 ^ i_input_data[507 % IN_WIDTH];
                753 / IN_WIDTH: ping_storage_data_547 <= (fillup_transition == 1'b1) ? i_input_data[753 % IN_WIDTH] : ping_storage_data_547 ^ i_input_data[753 % IN_WIDTH];
                1140 / IN_WIDTH: ping_storage_data_547 <= (fillup_transition == 1'b1) ? i_input_data[1140 % IN_WIDTH] : ping_storage_data_547 ^ i_input_data[1140 % IN_WIDTH];
                default: ping_storage_data_547 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_547;
                endcase
            end else begin
                case (input_count)
                405 / IN_WIDTH: pong_storage_data_547 <= (fillup_transition == 1'b1) ? i_input_data[405 % IN_WIDTH] : pong_storage_data_547 ^ i_input_data[405 % IN_WIDTH];
                507 / IN_WIDTH: pong_storage_data_547 <= (fillup_transition == 1'b1) ? i_input_data[507 % IN_WIDTH] : pong_storage_data_547 ^ i_input_data[507 % IN_WIDTH];
                753 / IN_WIDTH: pong_storage_data_547 <= (fillup_transition == 1'b1) ? i_input_data[753 % IN_WIDTH] : pong_storage_data_547 ^ i_input_data[753 % IN_WIDTH];
                1140 / IN_WIDTH: pong_storage_data_547 <= (fillup_transition == 1'b1) ? i_input_data[1140 % IN_WIDTH] : pong_storage_data_547 ^ i_input_data[1140 % IN_WIDTH];
                default: pong_storage_data_547 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_547;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_547 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_547;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_547 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_547;
            end
        end
    end
end

logic ping_storage_data_548;
logic pong_storage_data_548;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_548 <= 1'b0;
        pong_storage_data_548 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                406 / IN_WIDTH: ping_storage_data_548 <= (fillup_transition == 1'b1) ? i_input_data[406 % IN_WIDTH] : ping_storage_data_548 ^ i_input_data[406 % IN_WIDTH];
                508 / IN_WIDTH: ping_storage_data_548 <= (fillup_transition == 1'b1) ? i_input_data[508 % IN_WIDTH] : ping_storage_data_548 ^ i_input_data[508 % IN_WIDTH];
                754 / IN_WIDTH: ping_storage_data_548 <= (fillup_transition == 1'b1) ? i_input_data[754 % IN_WIDTH] : ping_storage_data_548 ^ i_input_data[754 % IN_WIDTH];
                1141 / IN_WIDTH: ping_storage_data_548 <= (fillup_transition == 1'b1) ? i_input_data[1141 % IN_WIDTH] : ping_storage_data_548 ^ i_input_data[1141 % IN_WIDTH];
                default: ping_storage_data_548 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_548;
                endcase
            end else begin
                case (input_count)
                406 / IN_WIDTH: pong_storage_data_548 <= (fillup_transition == 1'b1) ? i_input_data[406 % IN_WIDTH] : pong_storage_data_548 ^ i_input_data[406 % IN_WIDTH];
                508 / IN_WIDTH: pong_storage_data_548 <= (fillup_transition == 1'b1) ? i_input_data[508 % IN_WIDTH] : pong_storage_data_548 ^ i_input_data[508 % IN_WIDTH];
                754 / IN_WIDTH: pong_storage_data_548 <= (fillup_transition == 1'b1) ? i_input_data[754 % IN_WIDTH] : pong_storage_data_548 ^ i_input_data[754 % IN_WIDTH];
                1141 / IN_WIDTH: pong_storage_data_548 <= (fillup_transition == 1'b1) ? i_input_data[1141 % IN_WIDTH] : pong_storage_data_548 ^ i_input_data[1141 % IN_WIDTH];
                default: pong_storage_data_548 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_548;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_548 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_548;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_548 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_548;
            end
        end
    end
end

logic ping_storage_data_549;
logic pong_storage_data_549;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_549 <= 1'b0;
        pong_storage_data_549 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                407 / IN_WIDTH: ping_storage_data_549 <= (fillup_transition == 1'b1) ? i_input_data[407 % IN_WIDTH] : ping_storage_data_549 ^ i_input_data[407 % IN_WIDTH];
                509 / IN_WIDTH: ping_storage_data_549 <= (fillup_transition == 1'b1) ? i_input_data[509 % IN_WIDTH] : ping_storage_data_549 ^ i_input_data[509 % IN_WIDTH];
                755 / IN_WIDTH: ping_storage_data_549 <= (fillup_transition == 1'b1) ? i_input_data[755 % IN_WIDTH] : ping_storage_data_549 ^ i_input_data[755 % IN_WIDTH];
                1142 / IN_WIDTH: ping_storage_data_549 <= (fillup_transition == 1'b1) ? i_input_data[1142 % IN_WIDTH] : ping_storage_data_549 ^ i_input_data[1142 % IN_WIDTH];
                default: ping_storage_data_549 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_549;
                endcase
            end else begin
                case (input_count)
                407 / IN_WIDTH: pong_storage_data_549 <= (fillup_transition == 1'b1) ? i_input_data[407 % IN_WIDTH] : pong_storage_data_549 ^ i_input_data[407 % IN_WIDTH];
                509 / IN_WIDTH: pong_storage_data_549 <= (fillup_transition == 1'b1) ? i_input_data[509 % IN_WIDTH] : pong_storage_data_549 ^ i_input_data[509 % IN_WIDTH];
                755 / IN_WIDTH: pong_storage_data_549 <= (fillup_transition == 1'b1) ? i_input_data[755 % IN_WIDTH] : pong_storage_data_549 ^ i_input_data[755 % IN_WIDTH];
                1142 / IN_WIDTH: pong_storage_data_549 <= (fillup_transition == 1'b1) ? i_input_data[1142 % IN_WIDTH] : pong_storage_data_549 ^ i_input_data[1142 % IN_WIDTH];
                default: pong_storage_data_549 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_549;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_549 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_549;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_549 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_549;
            end
        end
    end
end

logic ping_storage_data_550;
logic pong_storage_data_550;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_550 <= 1'b0;
        pong_storage_data_550 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                408 / IN_WIDTH: ping_storage_data_550 <= (fillup_transition == 1'b1) ? i_input_data[408 % IN_WIDTH] : ping_storage_data_550 ^ i_input_data[408 % IN_WIDTH];
                510 / IN_WIDTH: ping_storage_data_550 <= (fillup_transition == 1'b1) ? i_input_data[510 % IN_WIDTH] : ping_storage_data_550 ^ i_input_data[510 % IN_WIDTH];
                756 / IN_WIDTH: ping_storage_data_550 <= (fillup_transition == 1'b1) ? i_input_data[756 % IN_WIDTH] : ping_storage_data_550 ^ i_input_data[756 % IN_WIDTH];
                1143 / IN_WIDTH: ping_storage_data_550 <= (fillup_transition == 1'b1) ? i_input_data[1143 % IN_WIDTH] : ping_storage_data_550 ^ i_input_data[1143 % IN_WIDTH];
                default: ping_storage_data_550 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_550;
                endcase
            end else begin
                case (input_count)
                408 / IN_WIDTH: pong_storage_data_550 <= (fillup_transition == 1'b1) ? i_input_data[408 % IN_WIDTH] : pong_storage_data_550 ^ i_input_data[408 % IN_WIDTH];
                510 / IN_WIDTH: pong_storage_data_550 <= (fillup_transition == 1'b1) ? i_input_data[510 % IN_WIDTH] : pong_storage_data_550 ^ i_input_data[510 % IN_WIDTH];
                756 / IN_WIDTH: pong_storage_data_550 <= (fillup_transition == 1'b1) ? i_input_data[756 % IN_WIDTH] : pong_storage_data_550 ^ i_input_data[756 % IN_WIDTH];
                1143 / IN_WIDTH: pong_storage_data_550 <= (fillup_transition == 1'b1) ? i_input_data[1143 % IN_WIDTH] : pong_storage_data_550 ^ i_input_data[1143 % IN_WIDTH];
                default: pong_storage_data_550 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_550;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_550 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_550;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_550 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_550;
            end
        end
    end
end

logic ping_storage_data_551;
logic pong_storage_data_551;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_551 <= 1'b0;
        pong_storage_data_551 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                409 / IN_WIDTH: ping_storage_data_551 <= (fillup_transition == 1'b1) ? i_input_data[409 % IN_WIDTH] : ping_storage_data_551 ^ i_input_data[409 % IN_WIDTH];
                511 / IN_WIDTH: ping_storage_data_551 <= (fillup_transition == 1'b1) ? i_input_data[511 % IN_WIDTH] : ping_storage_data_551 ^ i_input_data[511 % IN_WIDTH];
                757 / IN_WIDTH: ping_storage_data_551 <= (fillup_transition == 1'b1) ? i_input_data[757 % IN_WIDTH] : ping_storage_data_551 ^ i_input_data[757 % IN_WIDTH];
                1144 / IN_WIDTH: ping_storage_data_551 <= (fillup_transition == 1'b1) ? i_input_data[1144 % IN_WIDTH] : ping_storage_data_551 ^ i_input_data[1144 % IN_WIDTH];
                default: ping_storage_data_551 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_551;
                endcase
            end else begin
                case (input_count)
                409 / IN_WIDTH: pong_storage_data_551 <= (fillup_transition == 1'b1) ? i_input_data[409 % IN_WIDTH] : pong_storage_data_551 ^ i_input_data[409 % IN_WIDTH];
                511 / IN_WIDTH: pong_storage_data_551 <= (fillup_transition == 1'b1) ? i_input_data[511 % IN_WIDTH] : pong_storage_data_551 ^ i_input_data[511 % IN_WIDTH];
                757 / IN_WIDTH: pong_storage_data_551 <= (fillup_transition == 1'b1) ? i_input_data[757 % IN_WIDTH] : pong_storage_data_551 ^ i_input_data[757 % IN_WIDTH];
                1144 / IN_WIDTH: pong_storage_data_551 <= (fillup_transition == 1'b1) ? i_input_data[1144 % IN_WIDTH] : pong_storage_data_551 ^ i_input_data[1144 % IN_WIDTH];
                default: pong_storage_data_551 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_551;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_551 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_551;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_551 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_551;
            end
        end
    end
end

logic ping_storage_data_552;
logic pong_storage_data_552;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_552 <= 1'b0;
        pong_storage_data_552 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                410 / IN_WIDTH: ping_storage_data_552 <= (fillup_transition == 1'b1) ? i_input_data[410 % IN_WIDTH] : ping_storage_data_552 ^ i_input_data[410 % IN_WIDTH];
                512 / IN_WIDTH: ping_storage_data_552 <= (fillup_transition == 1'b1) ? i_input_data[512 % IN_WIDTH] : ping_storage_data_552 ^ i_input_data[512 % IN_WIDTH];
                758 / IN_WIDTH: ping_storage_data_552 <= (fillup_transition == 1'b1) ? i_input_data[758 % IN_WIDTH] : ping_storage_data_552 ^ i_input_data[758 % IN_WIDTH];
                1145 / IN_WIDTH: ping_storage_data_552 <= (fillup_transition == 1'b1) ? i_input_data[1145 % IN_WIDTH] : ping_storage_data_552 ^ i_input_data[1145 % IN_WIDTH];
                default: ping_storage_data_552 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_552;
                endcase
            end else begin
                case (input_count)
                410 / IN_WIDTH: pong_storage_data_552 <= (fillup_transition == 1'b1) ? i_input_data[410 % IN_WIDTH] : pong_storage_data_552 ^ i_input_data[410 % IN_WIDTH];
                512 / IN_WIDTH: pong_storage_data_552 <= (fillup_transition == 1'b1) ? i_input_data[512 % IN_WIDTH] : pong_storage_data_552 ^ i_input_data[512 % IN_WIDTH];
                758 / IN_WIDTH: pong_storage_data_552 <= (fillup_transition == 1'b1) ? i_input_data[758 % IN_WIDTH] : pong_storage_data_552 ^ i_input_data[758 % IN_WIDTH];
                1145 / IN_WIDTH: pong_storage_data_552 <= (fillup_transition == 1'b1) ? i_input_data[1145 % IN_WIDTH] : pong_storage_data_552 ^ i_input_data[1145 % IN_WIDTH];
                default: pong_storage_data_552 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_552;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_552 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_552;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_552 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_552;
            end
        end
    end
end

logic ping_storage_data_553;
logic pong_storage_data_553;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_553 <= 1'b0;
        pong_storage_data_553 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                411 / IN_WIDTH: ping_storage_data_553 <= (fillup_transition == 1'b1) ? i_input_data[411 % IN_WIDTH] : ping_storage_data_553 ^ i_input_data[411 % IN_WIDTH];
                513 / IN_WIDTH: ping_storage_data_553 <= (fillup_transition == 1'b1) ? i_input_data[513 % IN_WIDTH] : ping_storage_data_553 ^ i_input_data[513 % IN_WIDTH];
                759 / IN_WIDTH: ping_storage_data_553 <= (fillup_transition == 1'b1) ? i_input_data[759 % IN_WIDTH] : ping_storage_data_553 ^ i_input_data[759 % IN_WIDTH];
                1146 / IN_WIDTH: ping_storage_data_553 <= (fillup_transition == 1'b1) ? i_input_data[1146 % IN_WIDTH] : ping_storage_data_553 ^ i_input_data[1146 % IN_WIDTH];
                default: ping_storage_data_553 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_553;
                endcase
            end else begin
                case (input_count)
                411 / IN_WIDTH: pong_storage_data_553 <= (fillup_transition == 1'b1) ? i_input_data[411 % IN_WIDTH] : pong_storage_data_553 ^ i_input_data[411 % IN_WIDTH];
                513 / IN_WIDTH: pong_storage_data_553 <= (fillup_transition == 1'b1) ? i_input_data[513 % IN_WIDTH] : pong_storage_data_553 ^ i_input_data[513 % IN_WIDTH];
                759 / IN_WIDTH: pong_storage_data_553 <= (fillup_transition == 1'b1) ? i_input_data[759 % IN_WIDTH] : pong_storage_data_553 ^ i_input_data[759 % IN_WIDTH];
                1146 / IN_WIDTH: pong_storage_data_553 <= (fillup_transition == 1'b1) ? i_input_data[1146 % IN_WIDTH] : pong_storage_data_553 ^ i_input_data[1146 % IN_WIDTH];
                default: pong_storage_data_553 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_553;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_553 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_553;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_553 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_553;
            end
        end
    end
end

logic ping_storage_data_554;
logic pong_storage_data_554;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_554 <= 1'b0;
        pong_storage_data_554 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                412 / IN_WIDTH: ping_storage_data_554 <= (fillup_transition == 1'b1) ? i_input_data[412 % IN_WIDTH] : ping_storage_data_554 ^ i_input_data[412 % IN_WIDTH];
                514 / IN_WIDTH: ping_storage_data_554 <= (fillup_transition == 1'b1) ? i_input_data[514 % IN_WIDTH] : ping_storage_data_554 ^ i_input_data[514 % IN_WIDTH];
                760 / IN_WIDTH: ping_storage_data_554 <= (fillup_transition == 1'b1) ? i_input_data[760 % IN_WIDTH] : ping_storage_data_554 ^ i_input_data[760 % IN_WIDTH];
                1147 / IN_WIDTH: ping_storage_data_554 <= (fillup_transition == 1'b1) ? i_input_data[1147 % IN_WIDTH] : ping_storage_data_554 ^ i_input_data[1147 % IN_WIDTH];
                default: ping_storage_data_554 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_554;
                endcase
            end else begin
                case (input_count)
                412 / IN_WIDTH: pong_storage_data_554 <= (fillup_transition == 1'b1) ? i_input_data[412 % IN_WIDTH] : pong_storage_data_554 ^ i_input_data[412 % IN_WIDTH];
                514 / IN_WIDTH: pong_storage_data_554 <= (fillup_transition == 1'b1) ? i_input_data[514 % IN_WIDTH] : pong_storage_data_554 ^ i_input_data[514 % IN_WIDTH];
                760 / IN_WIDTH: pong_storage_data_554 <= (fillup_transition == 1'b1) ? i_input_data[760 % IN_WIDTH] : pong_storage_data_554 ^ i_input_data[760 % IN_WIDTH];
                1147 / IN_WIDTH: pong_storage_data_554 <= (fillup_transition == 1'b1) ? i_input_data[1147 % IN_WIDTH] : pong_storage_data_554 ^ i_input_data[1147 % IN_WIDTH];
                default: pong_storage_data_554 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_554;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_554 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_554;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_554 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_554;
            end
        end
    end
end

logic ping_storage_data_555;
logic pong_storage_data_555;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_555 <= 1'b0;
        pong_storage_data_555 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                413 / IN_WIDTH: ping_storage_data_555 <= (fillup_transition == 1'b1) ? i_input_data[413 % IN_WIDTH] : ping_storage_data_555 ^ i_input_data[413 % IN_WIDTH];
                515 / IN_WIDTH: ping_storage_data_555 <= (fillup_transition == 1'b1) ? i_input_data[515 % IN_WIDTH] : ping_storage_data_555 ^ i_input_data[515 % IN_WIDTH];
                761 / IN_WIDTH: ping_storage_data_555 <= (fillup_transition == 1'b1) ? i_input_data[761 % IN_WIDTH] : ping_storage_data_555 ^ i_input_data[761 % IN_WIDTH];
                1148 / IN_WIDTH: ping_storage_data_555 <= (fillup_transition == 1'b1) ? i_input_data[1148 % IN_WIDTH] : ping_storage_data_555 ^ i_input_data[1148 % IN_WIDTH];
                default: ping_storage_data_555 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_555;
                endcase
            end else begin
                case (input_count)
                413 / IN_WIDTH: pong_storage_data_555 <= (fillup_transition == 1'b1) ? i_input_data[413 % IN_WIDTH] : pong_storage_data_555 ^ i_input_data[413 % IN_WIDTH];
                515 / IN_WIDTH: pong_storage_data_555 <= (fillup_transition == 1'b1) ? i_input_data[515 % IN_WIDTH] : pong_storage_data_555 ^ i_input_data[515 % IN_WIDTH];
                761 / IN_WIDTH: pong_storage_data_555 <= (fillup_transition == 1'b1) ? i_input_data[761 % IN_WIDTH] : pong_storage_data_555 ^ i_input_data[761 % IN_WIDTH];
                1148 / IN_WIDTH: pong_storage_data_555 <= (fillup_transition == 1'b1) ? i_input_data[1148 % IN_WIDTH] : pong_storage_data_555 ^ i_input_data[1148 % IN_WIDTH];
                default: pong_storage_data_555 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_555;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_555 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_555;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_555 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_555;
            end
        end
    end
end

logic ping_storage_data_556;
logic pong_storage_data_556;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_556 <= 1'b0;
        pong_storage_data_556 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                414 / IN_WIDTH: ping_storage_data_556 <= (fillup_transition == 1'b1) ? i_input_data[414 % IN_WIDTH] : ping_storage_data_556 ^ i_input_data[414 % IN_WIDTH];
                516 / IN_WIDTH: ping_storage_data_556 <= (fillup_transition == 1'b1) ? i_input_data[516 % IN_WIDTH] : ping_storage_data_556 ^ i_input_data[516 % IN_WIDTH];
                762 / IN_WIDTH: ping_storage_data_556 <= (fillup_transition == 1'b1) ? i_input_data[762 % IN_WIDTH] : ping_storage_data_556 ^ i_input_data[762 % IN_WIDTH];
                1149 / IN_WIDTH: ping_storage_data_556 <= (fillup_transition == 1'b1) ? i_input_data[1149 % IN_WIDTH] : ping_storage_data_556 ^ i_input_data[1149 % IN_WIDTH];
                default: ping_storage_data_556 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_556;
                endcase
            end else begin
                case (input_count)
                414 / IN_WIDTH: pong_storage_data_556 <= (fillup_transition == 1'b1) ? i_input_data[414 % IN_WIDTH] : pong_storage_data_556 ^ i_input_data[414 % IN_WIDTH];
                516 / IN_WIDTH: pong_storage_data_556 <= (fillup_transition == 1'b1) ? i_input_data[516 % IN_WIDTH] : pong_storage_data_556 ^ i_input_data[516 % IN_WIDTH];
                762 / IN_WIDTH: pong_storage_data_556 <= (fillup_transition == 1'b1) ? i_input_data[762 % IN_WIDTH] : pong_storage_data_556 ^ i_input_data[762 % IN_WIDTH];
                1149 / IN_WIDTH: pong_storage_data_556 <= (fillup_transition == 1'b1) ? i_input_data[1149 % IN_WIDTH] : pong_storage_data_556 ^ i_input_data[1149 % IN_WIDTH];
                default: pong_storage_data_556 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_556;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_556 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_556;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_556 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_556;
            end
        end
    end
end

logic ping_storage_data_557;
logic pong_storage_data_557;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_557 <= 1'b0;
        pong_storage_data_557 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                415 / IN_WIDTH: ping_storage_data_557 <= (fillup_transition == 1'b1) ? i_input_data[415 % IN_WIDTH] : ping_storage_data_557 ^ i_input_data[415 % IN_WIDTH];
                517 / IN_WIDTH: ping_storage_data_557 <= (fillup_transition == 1'b1) ? i_input_data[517 % IN_WIDTH] : ping_storage_data_557 ^ i_input_data[517 % IN_WIDTH];
                763 / IN_WIDTH: ping_storage_data_557 <= (fillup_transition == 1'b1) ? i_input_data[763 % IN_WIDTH] : ping_storage_data_557 ^ i_input_data[763 % IN_WIDTH];
                1150 / IN_WIDTH: ping_storage_data_557 <= (fillup_transition == 1'b1) ? i_input_data[1150 % IN_WIDTH] : ping_storage_data_557 ^ i_input_data[1150 % IN_WIDTH];
                default: ping_storage_data_557 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_557;
                endcase
            end else begin
                case (input_count)
                415 / IN_WIDTH: pong_storage_data_557 <= (fillup_transition == 1'b1) ? i_input_data[415 % IN_WIDTH] : pong_storage_data_557 ^ i_input_data[415 % IN_WIDTH];
                517 / IN_WIDTH: pong_storage_data_557 <= (fillup_transition == 1'b1) ? i_input_data[517 % IN_WIDTH] : pong_storage_data_557 ^ i_input_data[517 % IN_WIDTH];
                763 / IN_WIDTH: pong_storage_data_557 <= (fillup_transition == 1'b1) ? i_input_data[763 % IN_WIDTH] : pong_storage_data_557 ^ i_input_data[763 % IN_WIDTH];
                1150 / IN_WIDTH: pong_storage_data_557 <= (fillup_transition == 1'b1) ? i_input_data[1150 % IN_WIDTH] : pong_storage_data_557 ^ i_input_data[1150 % IN_WIDTH];
                default: pong_storage_data_557 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_557;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_557 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_557;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_557 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_557;
            end
        end
    end
end

logic ping_storage_data_558;
logic pong_storage_data_558;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_558 <= 1'b0;
        pong_storage_data_558 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                416 / IN_WIDTH: ping_storage_data_558 <= (fillup_transition == 1'b1) ? i_input_data[416 % IN_WIDTH] : ping_storage_data_558 ^ i_input_data[416 % IN_WIDTH];
                518 / IN_WIDTH: ping_storage_data_558 <= (fillup_transition == 1'b1) ? i_input_data[518 % IN_WIDTH] : ping_storage_data_558 ^ i_input_data[518 % IN_WIDTH];
                764 / IN_WIDTH: ping_storage_data_558 <= (fillup_transition == 1'b1) ? i_input_data[764 % IN_WIDTH] : ping_storage_data_558 ^ i_input_data[764 % IN_WIDTH];
                1151 / IN_WIDTH: ping_storage_data_558 <= (fillup_transition == 1'b1) ? i_input_data[1151 % IN_WIDTH] : ping_storage_data_558 ^ i_input_data[1151 % IN_WIDTH];
                default: ping_storage_data_558 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_558;
                endcase
            end else begin
                case (input_count)
                416 / IN_WIDTH: pong_storage_data_558 <= (fillup_transition == 1'b1) ? i_input_data[416 % IN_WIDTH] : pong_storage_data_558 ^ i_input_data[416 % IN_WIDTH];
                518 / IN_WIDTH: pong_storage_data_558 <= (fillup_transition == 1'b1) ? i_input_data[518 % IN_WIDTH] : pong_storage_data_558 ^ i_input_data[518 % IN_WIDTH];
                764 / IN_WIDTH: pong_storage_data_558 <= (fillup_transition == 1'b1) ? i_input_data[764 % IN_WIDTH] : pong_storage_data_558 ^ i_input_data[764 % IN_WIDTH];
                1151 / IN_WIDTH: pong_storage_data_558 <= (fillup_transition == 1'b1) ? i_input_data[1151 % IN_WIDTH] : pong_storage_data_558 ^ i_input_data[1151 % IN_WIDTH];
                default: pong_storage_data_558 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_558;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_558 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_558;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_558 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_558;
            end
        end
    end
end

logic ping_storage_data_559;
logic pong_storage_data_559;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_559 <= 1'b0;
        pong_storage_data_559 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                417 / IN_WIDTH: ping_storage_data_559 <= (fillup_transition == 1'b1) ? i_input_data[417 % IN_WIDTH] : ping_storage_data_559 ^ i_input_data[417 % IN_WIDTH];
                519 / IN_WIDTH: ping_storage_data_559 <= (fillup_transition == 1'b1) ? i_input_data[519 % IN_WIDTH] : ping_storage_data_559 ^ i_input_data[519 % IN_WIDTH];
                765 / IN_WIDTH: ping_storage_data_559 <= (fillup_transition == 1'b1) ? i_input_data[765 % IN_WIDTH] : ping_storage_data_559 ^ i_input_data[765 % IN_WIDTH];
                1056 / IN_WIDTH: ping_storage_data_559 <= (fillup_transition == 1'b1) ? i_input_data[1056 % IN_WIDTH] : ping_storage_data_559 ^ i_input_data[1056 % IN_WIDTH];
                default: ping_storage_data_559 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_559;
                endcase
            end else begin
                case (input_count)
                417 / IN_WIDTH: pong_storage_data_559 <= (fillup_transition == 1'b1) ? i_input_data[417 % IN_WIDTH] : pong_storage_data_559 ^ i_input_data[417 % IN_WIDTH];
                519 / IN_WIDTH: pong_storage_data_559 <= (fillup_transition == 1'b1) ? i_input_data[519 % IN_WIDTH] : pong_storage_data_559 ^ i_input_data[519 % IN_WIDTH];
                765 / IN_WIDTH: pong_storage_data_559 <= (fillup_transition == 1'b1) ? i_input_data[765 % IN_WIDTH] : pong_storage_data_559 ^ i_input_data[765 % IN_WIDTH];
                1056 / IN_WIDTH: pong_storage_data_559 <= (fillup_transition == 1'b1) ? i_input_data[1056 % IN_WIDTH] : pong_storage_data_559 ^ i_input_data[1056 % IN_WIDTH];
                default: pong_storage_data_559 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_559;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_559 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_559;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_559 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_559;
            end
        end
    end
end

logic ping_storage_data_560;
logic pong_storage_data_560;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_560 <= 1'b0;
        pong_storage_data_560 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                418 / IN_WIDTH: ping_storage_data_560 <= (fillup_transition == 1'b1) ? i_input_data[418 % IN_WIDTH] : ping_storage_data_560 ^ i_input_data[418 % IN_WIDTH];
                520 / IN_WIDTH: ping_storage_data_560 <= (fillup_transition == 1'b1) ? i_input_data[520 % IN_WIDTH] : ping_storage_data_560 ^ i_input_data[520 % IN_WIDTH];
                766 / IN_WIDTH: ping_storage_data_560 <= (fillup_transition == 1'b1) ? i_input_data[766 % IN_WIDTH] : ping_storage_data_560 ^ i_input_data[766 % IN_WIDTH];
                1057 / IN_WIDTH: ping_storage_data_560 <= (fillup_transition == 1'b1) ? i_input_data[1057 % IN_WIDTH] : ping_storage_data_560 ^ i_input_data[1057 % IN_WIDTH];
                default: ping_storage_data_560 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_560;
                endcase
            end else begin
                case (input_count)
                418 / IN_WIDTH: pong_storage_data_560 <= (fillup_transition == 1'b1) ? i_input_data[418 % IN_WIDTH] : pong_storage_data_560 ^ i_input_data[418 % IN_WIDTH];
                520 / IN_WIDTH: pong_storage_data_560 <= (fillup_transition == 1'b1) ? i_input_data[520 % IN_WIDTH] : pong_storage_data_560 ^ i_input_data[520 % IN_WIDTH];
                766 / IN_WIDTH: pong_storage_data_560 <= (fillup_transition == 1'b1) ? i_input_data[766 % IN_WIDTH] : pong_storage_data_560 ^ i_input_data[766 % IN_WIDTH];
                1057 / IN_WIDTH: pong_storage_data_560 <= (fillup_transition == 1'b1) ? i_input_data[1057 % IN_WIDTH] : pong_storage_data_560 ^ i_input_data[1057 % IN_WIDTH];
                default: pong_storage_data_560 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_560;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_560 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_560;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_560 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_560;
            end
        end
    end
end

logic ping_storage_data_561;
logic pong_storage_data_561;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_561 <= 1'b0;
        pong_storage_data_561 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                419 / IN_WIDTH: ping_storage_data_561 <= (fillup_transition == 1'b1) ? i_input_data[419 % IN_WIDTH] : ping_storage_data_561 ^ i_input_data[419 % IN_WIDTH];
                521 / IN_WIDTH: ping_storage_data_561 <= (fillup_transition == 1'b1) ? i_input_data[521 % IN_WIDTH] : ping_storage_data_561 ^ i_input_data[521 % IN_WIDTH];
                767 / IN_WIDTH: ping_storage_data_561 <= (fillup_transition == 1'b1) ? i_input_data[767 % IN_WIDTH] : ping_storage_data_561 ^ i_input_data[767 % IN_WIDTH];
                1058 / IN_WIDTH: ping_storage_data_561 <= (fillup_transition == 1'b1) ? i_input_data[1058 % IN_WIDTH] : ping_storage_data_561 ^ i_input_data[1058 % IN_WIDTH];
                default: ping_storage_data_561 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_561;
                endcase
            end else begin
                case (input_count)
                419 / IN_WIDTH: pong_storage_data_561 <= (fillup_transition == 1'b1) ? i_input_data[419 % IN_WIDTH] : pong_storage_data_561 ^ i_input_data[419 % IN_WIDTH];
                521 / IN_WIDTH: pong_storage_data_561 <= (fillup_transition == 1'b1) ? i_input_data[521 % IN_WIDTH] : pong_storage_data_561 ^ i_input_data[521 % IN_WIDTH];
                767 / IN_WIDTH: pong_storage_data_561 <= (fillup_transition == 1'b1) ? i_input_data[767 % IN_WIDTH] : pong_storage_data_561 ^ i_input_data[767 % IN_WIDTH];
                1058 / IN_WIDTH: pong_storage_data_561 <= (fillup_transition == 1'b1) ? i_input_data[1058 % IN_WIDTH] : pong_storage_data_561 ^ i_input_data[1058 % IN_WIDTH];
                default: pong_storage_data_561 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_561;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_561 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_561;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_561 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_561;
            end
        end
    end
end

logic ping_storage_data_562;
logic pong_storage_data_562;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_562 <= 1'b0;
        pong_storage_data_562 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                420 / IN_WIDTH: ping_storage_data_562 <= (fillup_transition == 1'b1) ? i_input_data[420 % IN_WIDTH] : ping_storage_data_562 ^ i_input_data[420 % IN_WIDTH];
                522 / IN_WIDTH: ping_storage_data_562 <= (fillup_transition == 1'b1) ? i_input_data[522 % IN_WIDTH] : ping_storage_data_562 ^ i_input_data[522 % IN_WIDTH];
                672 / IN_WIDTH: ping_storage_data_562 <= (fillup_transition == 1'b1) ? i_input_data[672 % IN_WIDTH] : ping_storage_data_562 ^ i_input_data[672 % IN_WIDTH];
                1059 / IN_WIDTH: ping_storage_data_562 <= (fillup_transition == 1'b1) ? i_input_data[1059 % IN_WIDTH] : ping_storage_data_562 ^ i_input_data[1059 % IN_WIDTH];
                default: ping_storage_data_562 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_562;
                endcase
            end else begin
                case (input_count)
                420 / IN_WIDTH: pong_storage_data_562 <= (fillup_transition == 1'b1) ? i_input_data[420 % IN_WIDTH] : pong_storage_data_562 ^ i_input_data[420 % IN_WIDTH];
                522 / IN_WIDTH: pong_storage_data_562 <= (fillup_transition == 1'b1) ? i_input_data[522 % IN_WIDTH] : pong_storage_data_562 ^ i_input_data[522 % IN_WIDTH];
                672 / IN_WIDTH: pong_storage_data_562 <= (fillup_transition == 1'b1) ? i_input_data[672 % IN_WIDTH] : pong_storage_data_562 ^ i_input_data[672 % IN_WIDTH];
                1059 / IN_WIDTH: pong_storage_data_562 <= (fillup_transition == 1'b1) ? i_input_data[1059 % IN_WIDTH] : pong_storage_data_562 ^ i_input_data[1059 % IN_WIDTH];
                default: pong_storage_data_562 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_562;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_562 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_562;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_562 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_562;
            end
        end
    end
end

logic ping_storage_data_563;
logic pong_storage_data_563;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_563 <= 1'b0;
        pong_storage_data_563 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                421 / IN_WIDTH: ping_storage_data_563 <= (fillup_transition == 1'b1) ? i_input_data[421 % IN_WIDTH] : ping_storage_data_563 ^ i_input_data[421 % IN_WIDTH];
                523 / IN_WIDTH: ping_storage_data_563 <= (fillup_transition == 1'b1) ? i_input_data[523 % IN_WIDTH] : ping_storage_data_563 ^ i_input_data[523 % IN_WIDTH];
                673 / IN_WIDTH: ping_storage_data_563 <= (fillup_transition == 1'b1) ? i_input_data[673 % IN_WIDTH] : ping_storage_data_563 ^ i_input_data[673 % IN_WIDTH];
                1060 / IN_WIDTH: ping_storage_data_563 <= (fillup_transition == 1'b1) ? i_input_data[1060 % IN_WIDTH] : ping_storage_data_563 ^ i_input_data[1060 % IN_WIDTH];
                default: ping_storage_data_563 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_563;
                endcase
            end else begin
                case (input_count)
                421 / IN_WIDTH: pong_storage_data_563 <= (fillup_transition == 1'b1) ? i_input_data[421 % IN_WIDTH] : pong_storage_data_563 ^ i_input_data[421 % IN_WIDTH];
                523 / IN_WIDTH: pong_storage_data_563 <= (fillup_transition == 1'b1) ? i_input_data[523 % IN_WIDTH] : pong_storage_data_563 ^ i_input_data[523 % IN_WIDTH];
                673 / IN_WIDTH: pong_storage_data_563 <= (fillup_transition == 1'b1) ? i_input_data[673 % IN_WIDTH] : pong_storage_data_563 ^ i_input_data[673 % IN_WIDTH];
                1060 / IN_WIDTH: pong_storage_data_563 <= (fillup_transition == 1'b1) ? i_input_data[1060 % IN_WIDTH] : pong_storage_data_563 ^ i_input_data[1060 % IN_WIDTH];
                default: pong_storage_data_563 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_563;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_563 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_563;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_563 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_563;
            end
        end
    end
end

logic ping_storage_data_564;
logic pong_storage_data_564;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_564 <= 1'b0;
        pong_storage_data_564 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                422 / IN_WIDTH: ping_storage_data_564 <= (fillup_transition == 1'b1) ? i_input_data[422 % IN_WIDTH] : ping_storage_data_564 ^ i_input_data[422 % IN_WIDTH];
                524 / IN_WIDTH: ping_storage_data_564 <= (fillup_transition == 1'b1) ? i_input_data[524 % IN_WIDTH] : ping_storage_data_564 ^ i_input_data[524 % IN_WIDTH];
                674 / IN_WIDTH: ping_storage_data_564 <= (fillup_transition == 1'b1) ? i_input_data[674 % IN_WIDTH] : ping_storage_data_564 ^ i_input_data[674 % IN_WIDTH];
                1061 / IN_WIDTH: ping_storage_data_564 <= (fillup_transition == 1'b1) ? i_input_data[1061 % IN_WIDTH] : ping_storage_data_564 ^ i_input_data[1061 % IN_WIDTH];
                default: ping_storage_data_564 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_564;
                endcase
            end else begin
                case (input_count)
                422 / IN_WIDTH: pong_storage_data_564 <= (fillup_transition == 1'b1) ? i_input_data[422 % IN_WIDTH] : pong_storage_data_564 ^ i_input_data[422 % IN_WIDTH];
                524 / IN_WIDTH: pong_storage_data_564 <= (fillup_transition == 1'b1) ? i_input_data[524 % IN_WIDTH] : pong_storage_data_564 ^ i_input_data[524 % IN_WIDTH];
                674 / IN_WIDTH: pong_storage_data_564 <= (fillup_transition == 1'b1) ? i_input_data[674 % IN_WIDTH] : pong_storage_data_564 ^ i_input_data[674 % IN_WIDTH];
                1061 / IN_WIDTH: pong_storage_data_564 <= (fillup_transition == 1'b1) ? i_input_data[1061 % IN_WIDTH] : pong_storage_data_564 ^ i_input_data[1061 % IN_WIDTH];
                default: pong_storage_data_564 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_564;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_564 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_564;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_564 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_564;
            end
        end
    end
end

logic ping_storage_data_565;
logic pong_storage_data_565;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_565 <= 1'b0;
        pong_storage_data_565 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                423 / IN_WIDTH: ping_storage_data_565 <= (fillup_transition == 1'b1) ? i_input_data[423 % IN_WIDTH] : ping_storage_data_565 ^ i_input_data[423 % IN_WIDTH];
                525 / IN_WIDTH: ping_storage_data_565 <= (fillup_transition == 1'b1) ? i_input_data[525 % IN_WIDTH] : ping_storage_data_565 ^ i_input_data[525 % IN_WIDTH];
                675 / IN_WIDTH: ping_storage_data_565 <= (fillup_transition == 1'b1) ? i_input_data[675 % IN_WIDTH] : ping_storage_data_565 ^ i_input_data[675 % IN_WIDTH];
                1062 / IN_WIDTH: ping_storage_data_565 <= (fillup_transition == 1'b1) ? i_input_data[1062 % IN_WIDTH] : ping_storage_data_565 ^ i_input_data[1062 % IN_WIDTH];
                default: ping_storage_data_565 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_565;
                endcase
            end else begin
                case (input_count)
                423 / IN_WIDTH: pong_storage_data_565 <= (fillup_transition == 1'b1) ? i_input_data[423 % IN_WIDTH] : pong_storage_data_565 ^ i_input_data[423 % IN_WIDTH];
                525 / IN_WIDTH: pong_storage_data_565 <= (fillup_transition == 1'b1) ? i_input_data[525 % IN_WIDTH] : pong_storage_data_565 ^ i_input_data[525 % IN_WIDTH];
                675 / IN_WIDTH: pong_storage_data_565 <= (fillup_transition == 1'b1) ? i_input_data[675 % IN_WIDTH] : pong_storage_data_565 ^ i_input_data[675 % IN_WIDTH];
                1062 / IN_WIDTH: pong_storage_data_565 <= (fillup_transition == 1'b1) ? i_input_data[1062 % IN_WIDTH] : pong_storage_data_565 ^ i_input_data[1062 % IN_WIDTH];
                default: pong_storage_data_565 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_565;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_565 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_565;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_565 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_565;
            end
        end
    end
end

logic ping_storage_data_566;
logic pong_storage_data_566;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_566 <= 1'b0;
        pong_storage_data_566 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                424 / IN_WIDTH: ping_storage_data_566 <= (fillup_transition == 1'b1) ? i_input_data[424 % IN_WIDTH] : ping_storage_data_566 ^ i_input_data[424 % IN_WIDTH];
                526 / IN_WIDTH: ping_storage_data_566 <= (fillup_transition == 1'b1) ? i_input_data[526 % IN_WIDTH] : ping_storage_data_566 ^ i_input_data[526 % IN_WIDTH];
                676 / IN_WIDTH: ping_storage_data_566 <= (fillup_transition == 1'b1) ? i_input_data[676 % IN_WIDTH] : ping_storage_data_566 ^ i_input_data[676 % IN_WIDTH];
                1063 / IN_WIDTH: ping_storage_data_566 <= (fillup_transition == 1'b1) ? i_input_data[1063 % IN_WIDTH] : ping_storage_data_566 ^ i_input_data[1063 % IN_WIDTH];
                default: ping_storage_data_566 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_566;
                endcase
            end else begin
                case (input_count)
                424 / IN_WIDTH: pong_storage_data_566 <= (fillup_transition == 1'b1) ? i_input_data[424 % IN_WIDTH] : pong_storage_data_566 ^ i_input_data[424 % IN_WIDTH];
                526 / IN_WIDTH: pong_storage_data_566 <= (fillup_transition == 1'b1) ? i_input_data[526 % IN_WIDTH] : pong_storage_data_566 ^ i_input_data[526 % IN_WIDTH];
                676 / IN_WIDTH: pong_storage_data_566 <= (fillup_transition == 1'b1) ? i_input_data[676 % IN_WIDTH] : pong_storage_data_566 ^ i_input_data[676 % IN_WIDTH];
                1063 / IN_WIDTH: pong_storage_data_566 <= (fillup_transition == 1'b1) ? i_input_data[1063 % IN_WIDTH] : pong_storage_data_566 ^ i_input_data[1063 % IN_WIDTH];
                default: pong_storage_data_566 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_566;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_566 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_566;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_566 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_566;
            end
        end
    end
end

logic ping_storage_data_567;
logic pong_storage_data_567;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_567 <= 1'b0;
        pong_storage_data_567 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                425 / IN_WIDTH: ping_storage_data_567 <= (fillup_transition == 1'b1) ? i_input_data[425 % IN_WIDTH] : ping_storage_data_567 ^ i_input_data[425 % IN_WIDTH];
                527 / IN_WIDTH: ping_storage_data_567 <= (fillup_transition == 1'b1) ? i_input_data[527 % IN_WIDTH] : ping_storage_data_567 ^ i_input_data[527 % IN_WIDTH];
                677 / IN_WIDTH: ping_storage_data_567 <= (fillup_transition == 1'b1) ? i_input_data[677 % IN_WIDTH] : ping_storage_data_567 ^ i_input_data[677 % IN_WIDTH];
                1064 / IN_WIDTH: ping_storage_data_567 <= (fillup_transition == 1'b1) ? i_input_data[1064 % IN_WIDTH] : ping_storage_data_567 ^ i_input_data[1064 % IN_WIDTH];
                default: ping_storage_data_567 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_567;
                endcase
            end else begin
                case (input_count)
                425 / IN_WIDTH: pong_storage_data_567 <= (fillup_transition == 1'b1) ? i_input_data[425 % IN_WIDTH] : pong_storage_data_567 ^ i_input_data[425 % IN_WIDTH];
                527 / IN_WIDTH: pong_storage_data_567 <= (fillup_transition == 1'b1) ? i_input_data[527 % IN_WIDTH] : pong_storage_data_567 ^ i_input_data[527 % IN_WIDTH];
                677 / IN_WIDTH: pong_storage_data_567 <= (fillup_transition == 1'b1) ? i_input_data[677 % IN_WIDTH] : pong_storage_data_567 ^ i_input_data[677 % IN_WIDTH];
                1064 / IN_WIDTH: pong_storage_data_567 <= (fillup_transition == 1'b1) ? i_input_data[1064 % IN_WIDTH] : pong_storage_data_567 ^ i_input_data[1064 % IN_WIDTH];
                default: pong_storage_data_567 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_567;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_567 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_567;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_567 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_567;
            end
        end
    end
end

logic ping_storage_data_568;
logic pong_storage_data_568;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_568 <= 1'b0;
        pong_storage_data_568 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                426 / IN_WIDTH: ping_storage_data_568 <= (fillup_transition == 1'b1) ? i_input_data[426 % IN_WIDTH] : ping_storage_data_568 ^ i_input_data[426 % IN_WIDTH];
                528 / IN_WIDTH: ping_storage_data_568 <= (fillup_transition == 1'b1) ? i_input_data[528 % IN_WIDTH] : ping_storage_data_568 ^ i_input_data[528 % IN_WIDTH];
                678 / IN_WIDTH: ping_storage_data_568 <= (fillup_transition == 1'b1) ? i_input_data[678 % IN_WIDTH] : ping_storage_data_568 ^ i_input_data[678 % IN_WIDTH];
                1065 / IN_WIDTH: ping_storage_data_568 <= (fillup_transition == 1'b1) ? i_input_data[1065 % IN_WIDTH] : ping_storage_data_568 ^ i_input_data[1065 % IN_WIDTH];
                default: ping_storage_data_568 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_568;
                endcase
            end else begin
                case (input_count)
                426 / IN_WIDTH: pong_storage_data_568 <= (fillup_transition == 1'b1) ? i_input_data[426 % IN_WIDTH] : pong_storage_data_568 ^ i_input_data[426 % IN_WIDTH];
                528 / IN_WIDTH: pong_storage_data_568 <= (fillup_transition == 1'b1) ? i_input_data[528 % IN_WIDTH] : pong_storage_data_568 ^ i_input_data[528 % IN_WIDTH];
                678 / IN_WIDTH: pong_storage_data_568 <= (fillup_transition == 1'b1) ? i_input_data[678 % IN_WIDTH] : pong_storage_data_568 ^ i_input_data[678 % IN_WIDTH];
                1065 / IN_WIDTH: pong_storage_data_568 <= (fillup_transition == 1'b1) ? i_input_data[1065 % IN_WIDTH] : pong_storage_data_568 ^ i_input_data[1065 % IN_WIDTH];
                default: pong_storage_data_568 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_568;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_568 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_568;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_568 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_568;
            end
        end
    end
end

logic ping_storage_data_569;
logic pong_storage_data_569;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_569 <= 1'b0;
        pong_storage_data_569 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                427 / IN_WIDTH: ping_storage_data_569 <= (fillup_transition == 1'b1) ? i_input_data[427 % IN_WIDTH] : ping_storage_data_569 ^ i_input_data[427 % IN_WIDTH];
                529 / IN_WIDTH: ping_storage_data_569 <= (fillup_transition == 1'b1) ? i_input_data[529 % IN_WIDTH] : ping_storage_data_569 ^ i_input_data[529 % IN_WIDTH];
                679 / IN_WIDTH: ping_storage_data_569 <= (fillup_transition == 1'b1) ? i_input_data[679 % IN_WIDTH] : ping_storage_data_569 ^ i_input_data[679 % IN_WIDTH];
                1066 / IN_WIDTH: ping_storage_data_569 <= (fillup_transition == 1'b1) ? i_input_data[1066 % IN_WIDTH] : ping_storage_data_569 ^ i_input_data[1066 % IN_WIDTH];
                default: ping_storage_data_569 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_569;
                endcase
            end else begin
                case (input_count)
                427 / IN_WIDTH: pong_storage_data_569 <= (fillup_transition == 1'b1) ? i_input_data[427 % IN_WIDTH] : pong_storage_data_569 ^ i_input_data[427 % IN_WIDTH];
                529 / IN_WIDTH: pong_storage_data_569 <= (fillup_transition == 1'b1) ? i_input_data[529 % IN_WIDTH] : pong_storage_data_569 ^ i_input_data[529 % IN_WIDTH];
                679 / IN_WIDTH: pong_storage_data_569 <= (fillup_transition == 1'b1) ? i_input_data[679 % IN_WIDTH] : pong_storage_data_569 ^ i_input_data[679 % IN_WIDTH];
                1066 / IN_WIDTH: pong_storage_data_569 <= (fillup_transition == 1'b1) ? i_input_data[1066 % IN_WIDTH] : pong_storage_data_569 ^ i_input_data[1066 % IN_WIDTH];
                default: pong_storage_data_569 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_569;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_569 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_569;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_569 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_569;
            end
        end
    end
end

logic ping_storage_data_570;
logic pong_storage_data_570;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_570 <= 1'b0;
        pong_storage_data_570 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                428 / IN_WIDTH: ping_storage_data_570 <= (fillup_transition == 1'b1) ? i_input_data[428 % IN_WIDTH] : ping_storage_data_570 ^ i_input_data[428 % IN_WIDTH];
                530 / IN_WIDTH: ping_storage_data_570 <= (fillup_transition == 1'b1) ? i_input_data[530 % IN_WIDTH] : ping_storage_data_570 ^ i_input_data[530 % IN_WIDTH];
                680 / IN_WIDTH: ping_storage_data_570 <= (fillup_transition == 1'b1) ? i_input_data[680 % IN_WIDTH] : ping_storage_data_570 ^ i_input_data[680 % IN_WIDTH];
                1067 / IN_WIDTH: ping_storage_data_570 <= (fillup_transition == 1'b1) ? i_input_data[1067 % IN_WIDTH] : ping_storage_data_570 ^ i_input_data[1067 % IN_WIDTH];
                default: ping_storage_data_570 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_570;
                endcase
            end else begin
                case (input_count)
                428 / IN_WIDTH: pong_storage_data_570 <= (fillup_transition == 1'b1) ? i_input_data[428 % IN_WIDTH] : pong_storage_data_570 ^ i_input_data[428 % IN_WIDTH];
                530 / IN_WIDTH: pong_storage_data_570 <= (fillup_transition == 1'b1) ? i_input_data[530 % IN_WIDTH] : pong_storage_data_570 ^ i_input_data[530 % IN_WIDTH];
                680 / IN_WIDTH: pong_storage_data_570 <= (fillup_transition == 1'b1) ? i_input_data[680 % IN_WIDTH] : pong_storage_data_570 ^ i_input_data[680 % IN_WIDTH];
                1067 / IN_WIDTH: pong_storage_data_570 <= (fillup_transition == 1'b1) ? i_input_data[1067 % IN_WIDTH] : pong_storage_data_570 ^ i_input_data[1067 % IN_WIDTH];
                default: pong_storage_data_570 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_570;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_570 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_570;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_570 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_570;
            end
        end
    end
end

logic ping_storage_data_571;
logic pong_storage_data_571;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_571 <= 1'b0;
        pong_storage_data_571 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                429 / IN_WIDTH: ping_storage_data_571 <= (fillup_transition == 1'b1) ? i_input_data[429 % IN_WIDTH] : ping_storage_data_571 ^ i_input_data[429 % IN_WIDTH];
                531 / IN_WIDTH: ping_storage_data_571 <= (fillup_transition == 1'b1) ? i_input_data[531 % IN_WIDTH] : ping_storage_data_571 ^ i_input_data[531 % IN_WIDTH];
                681 / IN_WIDTH: ping_storage_data_571 <= (fillup_transition == 1'b1) ? i_input_data[681 % IN_WIDTH] : ping_storage_data_571 ^ i_input_data[681 % IN_WIDTH];
                1068 / IN_WIDTH: ping_storage_data_571 <= (fillup_transition == 1'b1) ? i_input_data[1068 % IN_WIDTH] : ping_storage_data_571 ^ i_input_data[1068 % IN_WIDTH];
                default: ping_storage_data_571 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_571;
                endcase
            end else begin
                case (input_count)
                429 / IN_WIDTH: pong_storage_data_571 <= (fillup_transition == 1'b1) ? i_input_data[429 % IN_WIDTH] : pong_storage_data_571 ^ i_input_data[429 % IN_WIDTH];
                531 / IN_WIDTH: pong_storage_data_571 <= (fillup_transition == 1'b1) ? i_input_data[531 % IN_WIDTH] : pong_storage_data_571 ^ i_input_data[531 % IN_WIDTH];
                681 / IN_WIDTH: pong_storage_data_571 <= (fillup_transition == 1'b1) ? i_input_data[681 % IN_WIDTH] : pong_storage_data_571 ^ i_input_data[681 % IN_WIDTH];
                1068 / IN_WIDTH: pong_storage_data_571 <= (fillup_transition == 1'b1) ? i_input_data[1068 % IN_WIDTH] : pong_storage_data_571 ^ i_input_data[1068 % IN_WIDTH];
                default: pong_storage_data_571 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_571;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_571 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_571;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_571 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_571;
            end
        end
    end
end

logic ping_storage_data_572;
logic pong_storage_data_572;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_572 <= 1'b0;
        pong_storage_data_572 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                430 / IN_WIDTH: ping_storage_data_572 <= (fillup_transition == 1'b1) ? i_input_data[430 % IN_WIDTH] : ping_storage_data_572 ^ i_input_data[430 % IN_WIDTH];
                532 / IN_WIDTH: ping_storage_data_572 <= (fillup_transition == 1'b1) ? i_input_data[532 % IN_WIDTH] : ping_storage_data_572 ^ i_input_data[532 % IN_WIDTH];
                682 / IN_WIDTH: ping_storage_data_572 <= (fillup_transition == 1'b1) ? i_input_data[682 % IN_WIDTH] : ping_storage_data_572 ^ i_input_data[682 % IN_WIDTH];
                1069 / IN_WIDTH: ping_storage_data_572 <= (fillup_transition == 1'b1) ? i_input_data[1069 % IN_WIDTH] : ping_storage_data_572 ^ i_input_data[1069 % IN_WIDTH];
                default: ping_storage_data_572 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_572;
                endcase
            end else begin
                case (input_count)
                430 / IN_WIDTH: pong_storage_data_572 <= (fillup_transition == 1'b1) ? i_input_data[430 % IN_WIDTH] : pong_storage_data_572 ^ i_input_data[430 % IN_WIDTH];
                532 / IN_WIDTH: pong_storage_data_572 <= (fillup_transition == 1'b1) ? i_input_data[532 % IN_WIDTH] : pong_storage_data_572 ^ i_input_data[532 % IN_WIDTH];
                682 / IN_WIDTH: pong_storage_data_572 <= (fillup_transition == 1'b1) ? i_input_data[682 % IN_WIDTH] : pong_storage_data_572 ^ i_input_data[682 % IN_WIDTH];
                1069 / IN_WIDTH: pong_storage_data_572 <= (fillup_transition == 1'b1) ? i_input_data[1069 % IN_WIDTH] : pong_storage_data_572 ^ i_input_data[1069 % IN_WIDTH];
                default: pong_storage_data_572 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_572;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_572 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_572;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_572 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_572;
            end
        end
    end
end

logic ping_storage_data_573;
logic pong_storage_data_573;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_573 <= 1'b0;
        pong_storage_data_573 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                431 / IN_WIDTH: ping_storage_data_573 <= (fillup_transition == 1'b1) ? i_input_data[431 % IN_WIDTH] : ping_storage_data_573 ^ i_input_data[431 % IN_WIDTH];
                533 / IN_WIDTH: ping_storage_data_573 <= (fillup_transition == 1'b1) ? i_input_data[533 % IN_WIDTH] : ping_storage_data_573 ^ i_input_data[533 % IN_WIDTH];
                683 / IN_WIDTH: ping_storage_data_573 <= (fillup_transition == 1'b1) ? i_input_data[683 % IN_WIDTH] : ping_storage_data_573 ^ i_input_data[683 % IN_WIDTH];
                1070 / IN_WIDTH: ping_storage_data_573 <= (fillup_transition == 1'b1) ? i_input_data[1070 % IN_WIDTH] : ping_storage_data_573 ^ i_input_data[1070 % IN_WIDTH];
                default: ping_storage_data_573 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_573;
                endcase
            end else begin
                case (input_count)
                431 / IN_WIDTH: pong_storage_data_573 <= (fillup_transition == 1'b1) ? i_input_data[431 % IN_WIDTH] : pong_storage_data_573 ^ i_input_data[431 % IN_WIDTH];
                533 / IN_WIDTH: pong_storage_data_573 <= (fillup_transition == 1'b1) ? i_input_data[533 % IN_WIDTH] : pong_storage_data_573 ^ i_input_data[533 % IN_WIDTH];
                683 / IN_WIDTH: pong_storage_data_573 <= (fillup_transition == 1'b1) ? i_input_data[683 % IN_WIDTH] : pong_storage_data_573 ^ i_input_data[683 % IN_WIDTH];
                1070 / IN_WIDTH: pong_storage_data_573 <= (fillup_transition == 1'b1) ? i_input_data[1070 % IN_WIDTH] : pong_storage_data_573 ^ i_input_data[1070 % IN_WIDTH];
                default: pong_storage_data_573 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_573;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_573 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_573;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_573 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_573;
            end
        end
    end
end

logic ping_storage_data_574;
logic pong_storage_data_574;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_574 <= 1'b0;
        pong_storage_data_574 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                432 / IN_WIDTH: ping_storage_data_574 <= (fillup_transition == 1'b1) ? i_input_data[432 % IN_WIDTH] : ping_storage_data_574 ^ i_input_data[432 % IN_WIDTH];
                534 / IN_WIDTH: ping_storage_data_574 <= (fillup_transition == 1'b1) ? i_input_data[534 % IN_WIDTH] : ping_storage_data_574 ^ i_input_data[534 % IN_WIDTH];
                684 / IN_WIDTH: ping_storage_data_574 <= (fillup_transition == 1'b1) ? i_input_data[684 % IN_WIDTH] : ping_storage_data_574 ^ i_input_data[684 % IN_WIDTH];
                1071 / IN_WIDTH: ping_storage_data_574 <= (fillup_transition == 1'b1) ? i_input_data[1071 % IN_WIDTH] : ping_storage_data_574 ^ i_input_data[1071 % IN_WIDTH];
                default: ping_storage_data_574 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_574;
                endcase
            end else begin
                case (input_count)
                432 / IN_WIDTH: pong_storage_data_574 <= (fillup_transition == 1'b1) ? i_input_data[432 % IN_WIDTH] : pong_storage_data_574 ^ i_input_data[432 % IN_WIDTH];
                534 / IN_WIDTH: pong_storage_data_574 <= (fillup_transition == 1'b1) ? i_input_data[534 % IN_WIDTH] : pong_storage_data_574 ^ i_input_data[534 % IN_WIDTH];
                684 / IN_WIDTH: pong_storage_data_574 <= (fillup_transition == 1'b1) ? i_input_data[684 % IN_WIDTH] : pong_storage_data_574 ^ i_input_data[684 % IN_WIDTH];
                1071 / IN_WIDTH: pong_storage_data_574 <= (fillup_transition == 1'b1) ? i_input_data[1071 % IN_WIDTH] : pong_storage_data_574 ^ i_input_data[1071 % IN_WIDTH];
                default: pong_storage_data_574 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_574;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_574 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_574;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_574 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_574;
            end
        end
    end
end

logic ping_storage_data_575;
logic pong_storage_data_575;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_575 <= 1'b0;
        pong_storage_data_575 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                433 / IN_WIDTH: ping_storage_data_575 <= (fillup_transition == 1'b1) ? i_input_data[433 % IN_WIDTH] : ping_storage_data_575 ^ i_input_data[433 % IN_WIDTH];
                535 / IN_WIDTH: ping_storage_data_575 <= (fillup_transition == 1'b1) ? i_input_data[535 % IN_WIDTH] : ping_storage_data_575 ^ i_input_data[535 % IN_WIDTH];
                685 / IN_WIDTH: ping_storage_data_575 <= (fillup_transition == 1'b1) ? i_input_data[685 % IN_WIDTH] : ping_storage_data_575 ^ i_input_data[685 % IN_WIDTH];
                1072 / IN_WIDTH: ping_storage_data_575 <= (fillup_transition == 1'b1) ? i_input_data[1072 % IN_WIDTH] : ping_storage_data_575 ^ i_input_data[1072 % IN_WIDTH];
                default: ping_storage_data_575 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_575;
                endcase
            end else begin
                case (input_count)
                433 / IN_WIDTH: pong_storage_data_575 <= (fillup_transition == 1'b1) ? i_input_data[433 % IN_WIDTH] : pong_storage_data_575 ^ i_input_data[433 % IN_WIDTH];
                535 / IN_WIDTH: pong_storage_data_575 <= (fillup_transition == 1'b1) ? i_input_data[535 % IN_WIDTH] : pong_storage_data_575 ^ i_input_data[535 % IN_WIDTH];
                685 / IN_WIDTH: pong_storage_data_575 <= (fillup_transition == 1'b1) ? i_input_data[685 % IN_WIDTH] : pong_storage_data_575 ^ i_input_data[685 % IN_WIDTH];
                1072 / IN_WIDTH: pong_storage_data_575 <= (fillup_transition == 1'b1) ? i_input_data[1072 % IN_WIDTH] : pong_storage_data_575 ^ i_input_data[1072 % IN_WIDTH];
                default: pong_storage_data_575 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_575;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_575 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_575;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_575 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_575;
            end
        end
    end
end

logic ping_storage_data_576;
logic pong_storage_data_576;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_576 <= 1'b0;
        pong_storage_data_576 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                193 / IN_WIDTH: ping_storage_data_576 <= (fillup_transition == 1'b1) ? i_input_data[193 % IN_WIDTH] : ping_storage_data_576 ^ i_input_data[193 % IN_WIDTH];
                331 / IN_WIDTH: ping_storage_data_576 <= (fillup_transition == 1'b1) ? i_input_data[331 % IN_WIDTH] : ping_storage_data_576 ^ i_input_data[331 % IN_WIDTH];
                946 / IN_WIDTH: ping_storage_data_576 <= (fillup_transition == 1'b1) ? i_input_data[946 % IN_WIDTH] : ping_storage_data_576 ^ i_input_data[946 % IN_WIDTH];
                1038 / IN_WIDTH: ping_storage_data_576 <= (fillup_transition == 1'b1) ? i_input_data[1038 % IN_WIDTH] : ping_storage_data_576 ^ i_input_data[1038 % IN_WIDTH];
                default: ping_storage_data_576 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_576;
                endcase
            end else begin
                case (input_count)
                193 / IN_WIDTH: pong_storage_data_576 <= (fillup_transition == 1'b1) ? i_input_data[193 % IN_WIDTH] : pong_storage_data_576 ^ i_input_data[193 % IN_WIDTH];
                331 / IN_WIDTH: pong_storage_data_576 <= (fillup_transition == 1'b1) ? i_input_data[331 % IN_WIDTH] : pong_storage_data_576 ^ i_input_data[331 % IN_WIDTH];
                946 / IN_WIDTH: pong_storage_data_576 <= (fillup_transition == 1'b1) ? i_input_data[946 % IN_WIDTH] : pong_storage_data_576 ^ i_input_data[946 % IN_WIDTH];
                1038 / IN_WIDTH: pong_storage_data_576 <= (fillup_transition == 1'b1) ? i_input_data[1038 % IN_WIDTH] : pong_storage_data_576 ^ i_input_data[1038 % IN_WIDTH];
                default: pong_storage_data_576 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_576;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_576 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_576;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_576 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_576;
            end
        end
    end
end

logic ping_storage_data_577;
logic pong_storage_data_577;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_577 <= 1'b0;
        pong_storage_data_577 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                194 / IN_WIDTH: ping_storage_data_577 <= (fillup_transition == 1'b1) ? i_input_data[194 % IN_WIDTH] : ping_storage_data_577 ^ i_input_data[194 % IN_WIDTH];
                332 / IN_WIDTH: ping_storage_data_577 <= (fillup_transition == 1'b1) ? i_input_data[332 % IN_WIDTH] : ping_storage_data_577 ^ i_input_data[332 % IN_WIDTH];
                947 / IN_WIDTH: ping_storage_data_577 <= (fillup_transition == 1'b1) ? i_input_data[947 % IN_WIDTH] : ping_storage_data_577 ^ i_input_data[947 % IN_WIDTH];
                1039 / IN_WIDTH: ping_storage_data_577 <= (fillup_transition == 1'b1) ? i_input_data[1039 % IN_WIDTH] : ping_storage_data_577 ^ i_input_data[1039 % IN_WIDTH];
                default: ping_storage_data_577 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_577;
                endcase
            end else begin
                case (input_count)
                194 / IN_WIDTH: pong_storage_data_577 <= (fillup_transition == 1'b1) ? i_input_data[194 % IN_WIDTH] : pong_storage_data_577 ^ i_input_data[194 % IN_WIDTH];
                332 / IN_WIDTH: pong_storage_data_577 <= (fillup_transition == 1'b1) ? i_input_data[332 % IN_WIDTH] : pong_storage_data_577 ^ i_input_data[332 % IN_WIDTH];
                947 / IN_WIDTH: pong_storage_data_577 <= (fillup_transition == 1'b1) ? i_input_data[947 % IN_WIDTH] : pong_storage_data_577 ^ i_input_data[947 % IN_WIDTH];
                1039 / IN_WIDTH: pong_storage_data_577 <= (fillup_transition == 1'b1) ? i_input_data[1039 % IN_WIDTH] : pong_storage_data_577 ^ i_input_data[1039 % IN_WIDTH];
                default: pong_storage_data_577 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_577;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_577 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_577;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_577 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_577;
            end
        end
    end
end

logic ping_storage_data_578;
logic pong_storage_data_578;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_578 <= 1'b0;
        pong_storage_data_578 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                195 / IN_WIDTH: ping_storage_data_578 <= (fillup_transition == 1'b1) ? i_input_data[195 % IN_WIDTH] : ping_storage_data_578 ^ i_input_data[195 % IN_WIDTH];
                333 / IN_WIDTH: ping_storage_data_578 <= (fillup_transition == 1'b1) ? i_input_data[333 % IN_WIDTH] : ping_storage_data_578 ^ i_input_data[333 % IN_WIDTH];
                948 / IN_WIDTH: ping_storage_data_578 <= (fillup_transition == 1'b1) ? i_input_data[948 % IN_WIDTH] : ping_storage_data_578 ^ i_input_data[948 % IN_WIDTH];
                1040 / IN_WIDTH: ping_storage_data_578 <= (fillup_transition == 1'b1) ? i_input_data[1040 % IN_WIDTH] : ping_storage_data_578 ^ i_input_data[1040 % IN_WIDTH];
                default: ping_storage_data_578 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_578;
                endcase
            end else begin
                case (input_count)
                195 / IN_WIDTH: pong_storage_data_578 <= (fillup_transition == 1'b1) ? i_input_data[195 % IN_WIDTH] : pong_storage_data_578 ^ i_input_data[195 % IN_WIDTH];
                333 / IN_WIDTH: pong_storage_data_578 <= (fillup_transition == 1'b1) ? i_input_data[333 % IN_WIDTH] : pong_storage_data_578 ^ i_input_data[333 % IN_WIDTH];
                948 / IN_WIDTH: pong_storage_data_578 <= (fillup_transition == 1'b1) ? i_input_data[948 % IN_WIDTH] : pong_storage_data_578 ^ i_input_data[948 % IN_WIDTH];
                1040 / IN_WIDTH: pong_storage_data_578 <= (fillup_transition == 1'b1) ? i_input_data[1040 % IN_WIDTH] : pong_storage_data_578 ^ i_input_data[1040 % IN_WIDTH];
                default: pong_storage_data_578 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_578;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_578 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_578;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_578 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_578;
            end
        end
    end
end

logic ping_storage_data_579;
logic pong_storage_data_579;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_579 <= 1'b0;
        pong_storage_data_579 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                196 / IN_WIDTH: ping_storage_data_579 <= (fillup_transition == 1'b1) ? i_input_data[196 % IN_WIDTH] : ping_storage_data_579 ^ i_input_data[196 % IN_WIDTH];
                334 / IN_WIDTH: ping_storage_data_579 <= (fillup_transition == 1'b1) ? i_input_data[334 % IN_WIDTH] : ping_storage_data_579 ^ i_input_data[334 % IN_WIDTH];
                949 / IN_WIDTH: ping_storage_data_579 <= (fillup_transition == 1'b1) ? i_input_data[949 % IN_WIDTH] : ping_storage_data_579 ^ i_input_data[949 % IN_WIDTH];
                1041 / IN_WIDTH: ping_storage_data_579 <= (fillup_transition == 1'b1) ? i_input_data[1041 % IN_WIDTH] : ping_storage_data_579 ^ i_input_data[1041 % IN_WIDTH];
                default: ping_storage_data_579 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_579;
                endcase
            end else begin
                case (input_count)
                196 / IN_WIDTH: pong_storage_data_579 <= (fillup_transition == 1'b1) ? i_input_data[196 % IN_WIDTH] : pong_storage_data_579 ^ i_input_data[196 % IN_WIDTH];
                334 / IN_WIDTH: pong_storage_data_579 <= (fillup_transition == 1'b1) ? i_input_data[334 % IN_WIDTH] : pong_storage_data_579 ^ i_input_data[334 % IN_WIDTH];
                949 / IN_WIDTH: pong_storage_data_579 <= (fillup_transition == 1'b1) ? i_input_data[949 % IN_WIDTH] : pong_storage_data_579 ^ i_input_data[949 % IN_WIDTH];
                1041 / IN_WIDTH: pong_storage_data_579 <= (fillup_transition == 1'b1) ? i_input_data[1041 % IN_WIDTH] : pong_storage_data_579 ^ i_input_data[1041 % IN_WIDTH];
                default: pong_storage_data_579 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_579;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_579 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_579;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_579 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_579;
            end
        end
    end
end

logic ping_storage_data_580;
logic pong_storage_data_580;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_580 <= 1'b0;
        pong_storage_data_580 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                197 / IN_WIDTH: ping_storage_data_580 <= (fillup_transition == 1'b1) ? i_input_data[197 % IN_WIDTH] : ping_storage_data_580 ^ i_input_data[197 % IN_WIDTH];
                335 / IN_WIDTH: ping_storage_data_580 <= (fillup_transition == 1'b1) ? i_input_data[335 % IN_WIDTH] : ping_storage_data_580 ^ i_input_data[335 % IN_WIDTH];
                950 / IN_WIDTH: ping_storage_data_580 <= (fillup_transition == 1'b1) ? i_input_data[950 % IN_WIDTH] : ping_storage_data_580 ^ i_input_data[950 % IN_WIDTH];
                1042 / IN_WIDTH: ping_storage_data_580 <= (fillup_transition == 1'b1) ? i_input_data[1042 % IN_WIDTH] : ping_storage_data_580 ^ i_input_data[1042 % IN_WIDTH];
                default: ping_storage_data_580 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_580;
                endcase
            end else begin
                case (input_count)
                197 / IN_WIDTH: pong_storage_data_580 <= (fillup_transition == 1'b1) ? i_input_data[197 % IN_WIDTH] : pong_storage_data_580 ^ i_input_data[197 % IN_WIDTH];
                335 / IN_WIDTH: pong_storage_data_580 <= (fillup_transition == 1'b1) ? i_input_data[335 % IN_WIDTH] : pong_storage_data_580 ^ i_input_data[335 % IN_WIDTH];
                950 / IN_WIDTH: pong_storage_data_580 <= (fillup_transition == 1'b1) ? i_input_data[950 % IN_WIDTH] : pong_storage_data_580 ^ i_input_data[950 % IN_WIDTH];
                1042 / IN_WIDTH: pong_storage_data_580 <= (fillup_transition == 1'b1) ? i_input_data[1042 % IN_WIDTH] : pong_storage_data_580 ^ i_input_data[1042 % IN_WIDTH];
                default: pong_storage_data_580 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_580;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_580 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_580;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_580 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_580;
            end
        end
    end
end

logic ping_storage_data_581;
logic pong_storage_data_581;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_581 <= 1'b0;
        pong_storage_data_581 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                198 / IN_WIDTH: ping_storage_data_581 <= (fillup_transition == 1'b1) ? i_input_data[198 % IN_WIDTH] : ping_storage_data_581 ^ i_input_data[198 % IN_WIDTH];
                336 / IN_WIDTH: ping_storage_data_581 <= (fillup_transition == 1'b1) ? i_input_data[336 % IN_WIDTH] : ping_storage_data_581 ^ i_input_data[336 % IN_WIDTH];
                951 / IN_WIDTH: ping_storage_data_581 <= (fillup_transition == 1'b1) ? i_input_data[951 % IN_WIDTH] : ping_storage_data_581 ^ i_input_data[951 % IN_WIDTH];
                1043 / IN_WIDTH: ping_storage_data_581 <= (fillup_transition == 1'b1) ? i_input_data[1043 % IN_WIDTH] : ping_storage_data_581 ^ i_input_data[1043 % IN_WIDTH];
                default: ping_storage_data_581 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_581;
                endcase
            end else begin
                case (input_count)
                198 / IN_WIDTH: pong_storage_data_581 <= (fillup_transition == 1'b1) ? i_input_data[198 % IN_WIDTH] : pong_storage_data_581 ^ i_input_data[198 % IN_WIDTH];
                336 / IN_WIDTH: pong_storage_data_581 <= (fillup_transition == 1'b1) ? i_input_data[336 % IN_WIDTH] : pong_storage_data_581 ^ i_input_data[336 % IN_WIDTH];
                951 / IN_WIDTH: pong_storage_data_581 <= (fillup_transition == 1'b1) ? i_input_data[951 % IN_WIDTH] : pong_storage_data_581 ^ i_input_data[951 % IN_WIDTH];
                1043 / IN_WIDTH: pong_storage_data_581 <= (fillup_transition == 1'b1) ? i_input_data[1043 % IN_WIDTH] : pong_storage_data_581 ^ i_input_data[1043 % IN_WIDTH];
                default: pong_storage_data_581 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_581;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_581 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_581;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_581 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_581;
            end
        end
    end
end

logic ping_storage_data_582;
logic pong_storage_data_582;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_582 <= 1'b0;
        pong_storage_data_582 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                199 / IN_WIDTH: ping_storage_data_582 <= (fillup_transition == 1'b1) ? i_input_data[199 % IN_WIDTH] : ping_storage_data_582 ^ i_input_data[199 % IN_WIDTH];
                337 / IN_WIDTH: ping_storage_data_582 <= (fillup_transition == 1'b1) ? i_input_data[337 % IN_WIDTH] : ping_storage_data_582 ^ i_input_data[337 % IN_WIDTH];
                952 / IN_WIDTH: ping_storage_data_582 <= (fillup_transition == 1'b1) ? i_input_data[952 % IN_WIDTH] : ping_storage_data_582 ^ i_input_data[952 % IN_WIDTH];
                1044 / IN_WIDTH: ping_storage_data_582 <= (fillup_transition == 1'b1) ? i_input_data[1044 % IN_WIDTH] : ping_storage_data_582 ^ i_input_data[1044 % IN_WIDTH];
                default: ping_storage_data_582 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_582;
                endcase
            end else begin
                case (input_count)
                199 / IN_WIDTH: pong_storage_data_582 <= (fillup_transition == 1'b1) ? i_input_data[199 % IN_WIDTH] : pong_storage_data_582 ^ i_input_data[199 % IN_WIDTH];
                337 / IN_WIDTH: pong_storage_data_582 <= (fillup_transition == 1'b1) ? i_input_data[337 % IN_WIDTH] : pong_storage_data_582 ^ i_input_data[337 % IN_WIDTH];
                952 / IN_WIDTH: pong_storage_data_582 <= (fillup_transition == 1'b1) ? i_input_data[952 % IN_WIDTH] : pong_storage_data_582 ^ i_input_data[952 % IN_WIDTH];
                1044 / IN_WIDTH: pong_storage_data_582 <= (fillup_transition == 1'b1) ? i_input_data[1044 % IN_WIDTH] : pong_storage_data_582 ^ i_input_data[1044 % IN_WIDTH];
                default: pong_storage_data_582 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_582;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_582 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_582;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_582 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_582;
            end
        end
    end
end

logic ping_storage_data_583;
logic pong_storage_data_583;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_583 <= 1'b0;
        pong_storage_data_583 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                200 / IN_WIDTH: ping_storage_data_583 <= (fillup_transition == 1'b1) ? i_input_data[200 % IN_WIDTH] : ping_storage_data_583 ^ i_input_data[200 % IN_WIDTH];
                338 / IN_WIDTH: ping_storage_data_583 <= (fillup_transition == 1'b1) ? i_input_data[338 % IN_WIDTH] : ping_storage_data_583 ^ i_input_data[338 % IN_WIDTH];
                953 / IN_WIDTH: ping_storage_data_583 <= (fillup_transition == 1'b1) ? i_input_data[953 % IN_WIDTH] : ping_storage_data_583 ^ i_input_data[953 % IN_WIDTH];
                1045 / IN_WIDTH: ping_storage_data_583 <= (fillup_transition == 1'b1) ? i_input_data[1045 % IN_WIDTH] : ping_storage_data_583 ^ i_input_data[1045 % IN_WIDTH];
                default: ping_storage_data_583 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_583;
                endcase
            end else begin
                case (input_count)
                200 / IN_WIDTH: pong_storage_data_583 <= (fillup_transition == 1'b1) ? i_input_data[200 % IN_WIDTH] : pong_storage_data_583 ^ i_input_data[200 % IN_WIDTH];
                338 / IN_WIDTH: pong_storage_data_583 <= (fillup_transition == 1'b1) ? i_input_data[338 % IN_WIDTH] : pong_storage_data_583 ^ i_input_data[338 % IN_WIDTH];
                953 / IN_WIDTH: pong_storage_data_583 <= (fillup_transition == 1'b1) ? i_input_data[953 % IN_WIDTH] : pong_storage_data_583 ^ i_input_data[953 % IN_WIDTH];
                1045 / IN_WIDTH: pong_storage_data_583 <= (fillup_transition == 1'b1) ? i_input_data[1045 % IN_WIDTH] : pong_storage_data_583 ^ i_input_data[1045 % IN_WIDTH];
                default: pong_storage_data_583 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_583;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_583 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_583;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_583 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_583;
            end
        end
    end
end

logic ping_storage_data_584;
logic pong_storage_data_584;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_584 <= 1'b0;
        pong_storage_data_584 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                201 / IN_WIDTH: ping_storage_data_584 <= (fillup_transition == 1'b1) ? i_input_data[201 % IN_WIDTH] : ping_storage_data_584 ^ i_input_data[201 % IN_WIDTH];
                339 / IN_WIDTH: ping_storage_data_584 <= (fillup_transition == 1'b1) ? i_input_data[339 % IN_WIDTH] : ping_storage_data_584 ^ i_input_data[339 % IN_WIDTH];
                954 / IN_WIDTH: ping_storage_data_584 <= (fillup_transition == 1'b1) ? i_input_data[954 % IN_WIDTH] : ping_storage_data_584 ^ i_input_data[954 % IN_WIDTH];
                1046 / IN_WIDTH: ping_storage_data_584 <= (fillup_transition == 1'b1) ? i_input_data[1046 % IN_WIDTH] : ping_storage_data_584 ^ i_input_data[1046 % IN_WIDTH];
                default: ping_storage_data_584 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_584;
                endcase
            end else begin
                case (input_count)
                201 / IN_WIDTH: pong_storage_data_584 <= (fillup_transition == 1'b1) ? i_input_data[201 % IN_WIDTH] : pong_storage_data_584 ^ i_input_data[201 % IN_WIDTH];
                339 / IN_WIDTH: pong_storage_data_584 <= (fillup_transition == 1'b1) ? i_input_data[339 % IN_WIDTH] : pong_storage_data_584 ^ i_input_data[339 % IN_WIDTH];
                954 / IN_WIDTH: pong_storage_data_584 <= (fillup_transition == 1'b1) ? i_input_data[954 % IN_WIDTH] : pong_storage_data_584 ^ i_input_data[954 % IN_WIDTH];
                1046 / IN_WIDTH: pong_storage_data_584 <= (fillup_transition == 1'b1) ? i_input_data[1046 % IN_WIDTH] : pong_storage_data_584 ^ i_input_data[1046 % IN_WIDTH];
                default: pong_storage_data_584 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_584;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_584 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_584;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_584 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_584;
            end
        end
    end
end

logic ping_storage_data_585;
logic pong_storage_data_585;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_585 <= 1'b0;
        pong_storage_data_585 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                202 / IN_WIDTH: ping_storage_data_585 <= (fillup_transition == 1'b1) ? i_input_data[202 % IN_WIDTH] : ping_storage_data_585 ^ i_input_data[202 % IN_WIDTH];
                340 / IN_WIDTH: ping_storage_data_585 <= (fillup_transition == 1'b1) ? i_input_data[340 % IN_WIDTH] : ping_storage_data_585 ^ i_input_data[340 % IN_WIDTH];
                955 / IN_WIDTH: ping_storage_data_585 <= (fillup_transition == 1'b1) ? i_input_data[955 % IN_WIDTH] : ping_storage_data_585 ^ i_input_data[955 % IN_WIDTH];
                1047 / IN_WIDTH: ping_storage_data_585 <= (fillup_transition == 1'b1) ? i_input_data[1047 % IN_WIDTH] : ping_storage_data_585 ^ i_input_data[1047 % IN_WIDTH];
                default: ping_storage_data_585 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_585;
                endcase
            end else begin
                case (input_count)
                202 / IN_WIDTH: pong_storage_data_585 <= (fillup_transition == 1'b1) ? i_input_data[202 % IN_WIDTH] : pong_storage_data_585 ^ i_input_data[202 % IN_WIDTH];
                340 / IN_WIDTH: pong_storage_data_585 <= (fillup_transition == 1'b1) ? i_input_data[340 % IN_WIDTH] : pong_storage_data_585 ^ i_input_data[340 % IN_WIDTH];
                955 / IN_WIDTH: pong_storage_data_585 <= (fillup_transition == 1'b1) ? i_input_data[955 % IN_WIDTH] : pong_storage_data_585 ^ i_input_data[955 % IN_WIDTH];
                1047 / IN_WIDTH: pong_storage_data_585 <= (fillup_transition == 1'b1) ? i_input_data[1047 % IN_WIDTH] : pong_storage_data_585 ^ i_input_data[1047 % IN_WIDTH];
                default: pong_storage_data_585 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_585;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_585 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_585;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_585 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_585;
            end
        end
    end
end

logic ping_storage_data_586;
logic pong_storage_data_586;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_586 <= 1'b0;
        pong_storage_data_586 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                203 / IN_WIDTH: ping_storage_data_586 <= (fillup_transition == 1'b1) ? i_input_data[203 % IN_WIDTH] : ping_storage_data_586 ^ i_input_data[203 % IN_WIDTH];
                341 / IN_WIDTH: ping_storage_data_586 <= (fillup_transition == 1'b1) ? i_input_data[341 % IN_WIDTH] : ping_storage_data_586 ^ i_input_data[341 % IN_WIDTH];
                956 / IN_WIDTH: ping_storage_data_586 <= (fillup_transition == 1'b1) ? i_input_data[956 % IN_WIDTH] : ping_storage_data_586 ^ i_input_data[956 % IN_WIDTH];
                1048 / IN_WIDTH: ping_storage_data_586 <= (fillup_transition == 1'b1) ? i_input_data[1048 % IN_WIDTH] : ping_storage_data_586 ^ i_input_data[1048 % IN_WIDTH];
                default: ping_storage_data_586 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_586;
                endcase
            end else begin
                case (input_count)
                203 / IN_WIDTH: pong_storage_data_586 <= (fillup_transition == 1'b1) ? i_input_data[203 % IN_WIDTH] : pong_storage_data_586 ^ i_input_data[203 % IN_WIDTH];
                341 / IN_WIDTH: pong_storage_data_586 <= (fillup_transition == 1'b1) ? i_input_data[341 % IN_WIDTH] : pong_storage_data_586 ^ i_input_data[341 % IN_WIDTH];
                956 / IN_WIDTH: pong_storage_data_586 <= (fillup_transition == 1'b1) ? i_input_data[956 % IN_WIDTH] : pong_storage_data_586 ^ i_input_data[956 % IN_WIDTH];
                1048 / IN_WIDTH: pong_storage_data_586 <= (fillup_transition == 1'b1) ? i_input_data[1048 % IN_WIDTH] : pong_storage_data_586 ^ i_input_data[1048 % IN_WIDTH];
                default: pong_storage_data_586 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_586;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_586 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_586;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_586 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_586;
            end
        end
    end
end

logic ping_storage_data_587;
logic pong_storage_data_587;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_587 <= 1'b0;
        pong_storage_data_587 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                204 / IN_WIDTH: ping_storage_data_587 <= (fillup_transition == 1'b1) ? i_input_data[204 % IN_WIDTH] : ping_storage_data_587 ^ i_input_data[204 % IN_WIDTH];
                342 / IN_WIDTH: ping_storage_data_587 <= (fillup_transition == 1'b1) ? i_input_data[342 % IN_WIDTH] : ping_storage_data_587 ^ i_input_data[342 % IN_WIDTH];
                957 / IN_WIDTH: ping_storage_data_587 <= (fillup_transition == 1'b1) ? i_input_data[957 % IN_WIDTH] : ping_storage_data_587 ^ i_input_data[957 % IN_WIDTH];
                1049 / IN_WIDTH: ping_storage_data_587 <= (fillup_transition == 1'b1) ? i_input_data[1049 % IN_WIDTH] : ping_storage_data_587 ^ i_input_data[1049 % IN_WIDTH];
                default: ping_storage_data_587 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_587;
                endcase
            end else begin
                case (input_count)
                204 / IN_WIDTH: pong_storage_data_587 <= (fillup_transition == 1'b1) ? i_input_data[204 % IN_WIDTH] : pong_storage_data_587 ^ i_input_data[204 % IN_WIDTH];
                342 / IN_WIDTH: pong_storage_data_587 <= (fillup_transition == 1'b1) ? i_input_data[342 % IN_WIDTH] : pong_storage_data_587 ^ i_input_data[342 % IN_WIDTH];
                957 / IN_WIDTH: pong_storage_data_587 <= (fillup_transition == 1'b1) ? i_input_data[957 % IN_WIDTH] : pong_storage_data_587 ^ i_input_data[957 % IN_WIDTH];
                1049 / IN_WIDTH: pong_storage_data_587 <= (fillup_transition == 1'b1) ? i_input_data[1049 % IN_WIDTH] : pong_storage_data_587 ^ i_input_data[1049 % IN_WIDTH];
                default: pong_storage_data_587 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_587;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_587 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_587;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_587 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_587;
            end
        end
    end
end

logic ping_storage_data_588;
logic pong_storage_data_588;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_588 <= 1'b0;
        pong_storage_data_588 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                205 / IN_WIDTH: ping_storage_data_588 <= (fillup_transition == 1'b1) ? i_input_data[205 % IN_WIDTH] : ping_storage_data_588 ^ i_input_data[205 % IN_WIDTH];
                343 / IN_WIDTH: ping_storage_data_588 <= (fillup_transition == 1'b1) ? i_input_data[343 % IN_WIDTH] : ping_storage_data_588 ^ i_input_data[343 % IN_WIDTH];
                958 / IN_WIDTH: ping_storage_data_588 <= (fillup_transition == 1'b1) ? i_input_data[958 % IN_WIDTH] : ping_storage_data_588 ^ i_input_data[958 % IN_WIDTH];
                1050 / IN_WIDTH: ping_storage_data_588 <= (fillup_transition == 1'b1) ? i_input_data[1050 % IN_WIDTH] : ping_storage_data_588 ^ i_input_data[1050 % IN_WIDTH];
                default: ping_storage_data_588 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_588;
                endcase
            end else begin
                case (input_count)
                205 / IN_WIDTH: pong_storage_data_588 <= (fillup_transition == 1'b1) ? i_input_data[205 % IN_WIDTH] : pong_storage_data_588 ^ i_input_data[205 % IN_WIDTH];
                343 / IN_WIDTH: pong_storage_data_588 <= (fillup_transition == 1'b1) ? i_input_data[343 % IN_WIDTH] : pong_storage_data_588 ^ i_input_data[343 % IN_WIDTH];
                958 / IN_WIDTH: pong_storage_data_588 <= (fillup_transition == 1'b1) ? i_input_data[958 % IN_WIDTH] : pong_storage_data_588 ^ i_input_data[958 % IN_WIDTH];
                1050 / IN_WIDTH: pong_storage_data_588 <= (fillup_transition == 1'b1) ? i_input_data[1050 % IN_WIDTH] : pong_storage_data_588 ^ i_input_data[1050 % IN_WIDTH];
                default: pong_storage_data_588 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_588;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_588 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_588;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_588 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_588;
            end
        end
    end
end

logic ping_storage_data_589;
logic pong_storage_data_589;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_589 <= 1'b0;
        pong_storage_data_589 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                206 / IN_WIDTH: ping_storage_data_589 <= (fillup_transition == 1'b1) ? i_input_data[206 % IN_WIDTH] : ping_storage_data_589 ^ i_input_data[206 % IN_WIDTH];
                344 / IN_WIDTH: ping_storage_data_589 <= (fillup_transition == 1'b1) ? i_input_data[344 % IN_WIDTH] : ping_storage_data_589 ^ i_input_data[344 % IN_WIDTH];
                959 / IN_WIDTH: ping_storage_data_589 <= (fillup_transition == 1'b1) ? i_input_data[959 % IN_WIDTH] : ping_storage_data_589 ^ i_input_data[959 % IN_WIDTH];
                1051 / IN_WIDTH: ping_storage_data_589 <= (fillup_transition == 1'b1) ? i_input_data[1051 % IN_WIDTH] : ping_storage_data_589 ^ i_input_data[1051 % IN_WIDTH];
                default: ping_storage_data_589 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_589;
                endcase
            end else begin
                case (input_count)
                206 / IN_WIDTH: pong_storage_data_589 <= (fillup_transition == 1'b1) ? i_input_data[206 % IN_WIDTH] : pong_storage_data_589 ^ i_input_data[206 % IN_WIDTH];
                344 / IN_WIDTH: pong_storage_data_589 <= (fillup_transition == 1'b1) ? i_input_data[344 % IN_WIDTH] : pong_storage_data_589 ^ i_input_data[344 % IN_WIDTH];
                959 / IN_WIDTH: pong_storage_data_589 <= (fillup_transition == 1'b1) ? i_input_data[959 % IN_WIDTH] : pong_storage_data_589 ^ i_input_data[959 % IN_WIDTH];
                1051 / IN_WIDTH: pong_storage_data_589 <= (fillup_transition == 1'b1) ? i_input_data[1051 % IN_WIDTH] : pong_storage_data_589 ^ i_input_data[1051 % IN_WIDTH];
                default: pong_storage_data_589 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_589;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_589 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_589;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_589 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_589;
            end
        end
    end
end

logic ping_storage_data_590;
logic pong_storage_data_590;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_590 <= 1'b0;
        pong_storage_data_590 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                207 / IN_WIDTH: ping_storage_data_590 <= (fillup_transition == 1'b1) ? i_input_data[207 % IN_WIDTH] : ping_storage_data_590 ^ i_input_data[207 % IN_WIDTH];
                345 / IN_WIDTH: ping_storage_data_590 <= (fillup_transition == 1'b1) ? i_input_data[345 % IN_WIDTH] : ping_storage_data_590 ^ i_input_data[345 % IN_WIDTH];
                864 / IN_WIDTH: ping_storage_data_590 <= (fillup_transition == 1'b1) ? i_input_data[864 % IN_WIDTH] : ping_storage_data_590 ^ i_input_data[864 % IN_WIDTH];
                1052 / IN_WIDTH: ping_storage_data_590 <= (fillup_transition == 1'b1) ? i_input_data[1052 % IN_WIDTH] : ping_storage_data_590 ^ i_input_data[1052 % IN_WIDTH];
                default: ping_storage_data_590 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_590;
                endcase
            end else begin
                case (input_count)
                207 / IN_WIDTH: pong_storage_data_590 <= (fillup_transition == 1'b1) ? i_input_data[207 % IN_WIDTH] : pong_storage_data_590 ^ i_input_data[207 % IN_WIDTH];
                345 / IN_WIDTH: pong_storage_data_590 <= (fillup_transition == 1'b1) ? i_input_data[345 % IN_WIDTH] : pong_storage_data_590 ^ i_input_data[345 % IN_WIDTH];
                864 / IN_WIDTH: pong_storage_data_590 <= (fillup_transition == 1'b1) ? i_input_data[864 % IN_WIDTH] : pong_storage_data_590 ^ i_input_data[864 % IN_WIDTH];
                1052 / IN_WIDTH: pong_storage_data_590 <= (fillup_transition == 1'b1) ? i_input_data[1052 % IN_WIDTH] : pong_storage_data_590 ^ i_input_data[1052 % IN_WIDTH];
                default: pong_storage_data_590 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_590;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_590 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_590;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_590 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_590;
            end
        end
    end
end

logic ping_storage_data_591;
logic pong_storage_data_591;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_591 <= 1'b0;
        pong_storage_data_591 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                208 / IN_WIDTH: ping_storage_data_591 <= (fillup_transition == 1'b1) ? i_input_data[208 % IN_WIDTH] : ping_storage_data_591 ^ i_input_data[208 % IN_WIDTH];
                346 / IN_WIDTH: ping_storage_data_591 <= (fillup_transition == 1'b1) ? i_input_data[346 % IN_WIDTH] : ping_storage_data_591 ^ i_input_data[346 % IN_WIDTH];
                865 / IN_WIDTH: ping_storage_data_591 <= (fillup_transition == 1'b1) ? i_input_data[865 % IN_WIDTH] : ping_storage_data_591 ^ i_input_data[865 % IN_WIDTH];
                1053 / IN_WIDTH: ping_storage_data_591 <= (fillup_transition == 1'b1) ? i_input_data[1053 % IN_WIDTH] : ping_storage_data_591 ^ i_input_data[1053 % IN_WIDTH];
                default: ping_storage_data_591 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_591;
                endcase
            end else begin
                case (input_count)
                208 / IN_WIDTH: pong_storage_data_591 <= (fillup_transition == 1'b1) ? i_input_data[208 % IN_WIDTH] : pong_storage_data_591 ^ i_input_data[208 % IN_WIDTH];
                346 / IN_WIDTH: pong_storage_data_591 <= (fillup_transition == 1'b1) ? i_input_data[346 % IN_WIDTH] : pong_storage_data_591 ^ i_input_data[346 % IN_WIDTH];
                865 / IN_WIDTH: pong_storage_data_591 <= (fillup_transition == 1'b1) ? i_input_data[865 % IN_WIDTH] : pong_storage_data_591 ^ i_input_data[865 % IN_WIDTH];
                1053 / IN_WIDTH: pong_storage_data_591 <= (fillup_transition == 1'b1) ? i_input_data[1053 % IN_WIDTH] : pong_storage_data_591 ^ i_input_data[1053 % IN_WIDTH];
                default: pong_storage_data_591 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_591;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_591 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_591;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_591 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_591;
            end
        end
    end
end

logic ping_storage_data_592;
logic pong_storage_data_592;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_592 <= 1'b0;
        pong_storage_data_592 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                209 / IN_WIDTH: ping_storage_data_592 <= (fillup_transition == 1'b1) ? i_input_data[209 % IN_WIDTH] : ping_storage_data_592 ^ i_input_data[209 % IN_WIDTH];
                347 / IN_WIDTH: ping_storage_data_592 <= (fillup_transition == 1'b1) ? i_input_data[347 % IN_WIDTH] : ping_storage_data_592 ^ i_input_data[347 % IN_WIDTH];
                866 / IN_WIDTH: ping_storage_data_592 <= (fillup_transition == 1'b1) ? i_input_data[866 % IN_WIDTH] : ping_storage_data_592 ^ i_input_data[866 % IN_WIDTH];
                1054 / IN_WIDTH: ping_storage_data_592 <= (fillup_transition == 1'b1) ? i_input_data[1054 % IN_WIDTH] : ping_storage_data_592 ^ i_input_data[1054 % IN_WIDTH];
                default: ping_storage_data_592 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_592;
                endcase
            end else begin
                case (input_count)
                209 / IN_WIDTH: pong_storage_data_592 <= (fillup_transition == 1'b1) ? i_input_data[209 % IN_WIDTH] : pong_storage_data_592 ^ i_input_data[209 % IN_WIDTH];
                347 / IN_WIDTH: pong_storage_data_592 <= (fillup_transition == 1'b1) ? i_input_data[347 % IN_WIDTH] : pong_storage_data_592 ^ i_input_data[347 % IN_WIDTH];
                866 / IN_WIDTH: pong_storage_data_592 <= (fillup_transition == 1'b1) ? i_input_data[866 % IN_WIDTH] : pong_storage_data_592 ^ i_input_data[866 % IN_WIDTH];
                1054 / IN_WIDTH: pong_storage_data_592 <= (fillup_transition == 1'b1) ? i_input_data[1054 % IN_WIDTH] : pong_storage_data_592 ^ i_input_data[1054 % IN_WIDTH];
                default: pong_storage_data_592 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_592;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_592 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_592;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_592 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_592;
            end
        end
    end
end

logic ping_storage_data_593;
logic pong_storage_data_593;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_593 <= 1'b0;
        pong_storage_data_593 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                210 / IN_WIDTH: ping_storage_data_593 <= (fillup_transition == 1'b1) ? i_input_data[210 % IN_WIDTH] : ping_storage_data_593 ^ i_input_data[210 % IN_WIDTH];
                348 / IN_WIDTH: ping_storage_data_593 <= (fillup_transition == 1'b1) ? i_input_data[348 % IN_WIDTH] : ping_storage_data_593 ^ i_input_data[348 % IN_WIDTH];
                867 / IN_WIDTH: ping_storage_data_593 <= (fillup_transition == 1'b1) ? i_input_data[867 % IN_WIDTH] : ping_storage_data_593 ^ i_input_data[867 % IN_WIDTH];
                1055 / IN_WIDTH: ping_storage_data_593 <= (fillup_transition == 1'b1) ? i_input_data[1055 % IN_WIDTH] : ping_storage_data_593 ^ i_input_data[1055 % IN_WIDTH];
                default: ping_storage_data_593 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_593;
                endcase
            end else begin
                case (input_count)
                210 / IN_WIDTH: pong_storage_data_593 <= (fillup_transition == 1'b1) ? i_input_data[210 % IN_WIDTH] : pong_storage_data_593 ^ i_input_data[210 % IN_WIDTH];
                348 / IN_WIDTH: pong_storage_data_593 <= (fillup_transition == 1'b1) ? i_input_data[348 % IN_WIDTH] : pong_storage_data_593 ^ i_input_data[348 % IN_WIDTH];
                867 / IN_WIDTH: pong_storage_data_593 <= (fillup_transition == 1'b1) ? i_input_data[867 % IN_WIDTH] : pong_storage_data_593 ^ i_input_data[867 % IN_WIDTH];
                1055 / IN_WIDTH: pong_storage_data_593 <= (fillup_transition == 1'b1) ? i_input_data[1055 % IN_WIDTH] : pong_storage_data_593 ^ i_input_data[1055 % IN_WIDTH];
                default: pong_storage_data_593 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_593;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_593 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_593;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_593 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_593;
            end
        end
    end
end

logic ping_storage_data_594;
logic pong_storage_data_594;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_594 <= 1'b0;
        pong_storage_data_594 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                211 / IN_WIDTH: ping_storage_data_594 <= (fillup_transition == 1'b1) ? i_input_data[211 % IN_WIDTH] : ping_storage_data_594 ^ i_input_data[211 % IN_WIDTH];
                349 / IN_WIDTH: ping_storage_data_594 <= (fillup_transition == 1'b1) ? i_input_data[349 % IN_WIDTH] : ping_storage_data_594 ^ i_input_data[349 % IN_WIDTH];
                868 / IN_WIDTH: ping_storage_data_594 <= (fillup_transition == 1'b1) ? i_input_data[868 % IN_WIDTH] : ping_storage_data_594 ^ i_input_data[868 % IN_WIDTH];
                960 / IN_WIDTH: ping_storage_data_594 <= (fillup_transition == 1'b1) ? i_input_data[960 % IN_WIDTH] : ping_storage_data_594 ^ i_input_data[960 % IN_WIDTH];
                default: ping_storage_data_594 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_594;
                endcase
            end else begin
                case (input_count)
                211 / IN_WIDTH: pong_storage_data_594 <= (fillup_transition == 1'b1) ? i_input_data[211 % IN_WIDTH] : pong_storage_data_594 ^ i_input_data[211 % IN_WIDTH];
                349 / IN_WIDTH: pong_storage_data_594 <= (fillup_transition == 1'b1) ? i_input_data[349 % IN_WIDTH] : pong_storage_data_594 ^ i_input_data[349 % IN_WIDTH];
                868 / IN_WIDTH: pong_storage_data_594 <= (fillup_transition == 1'b1) ? i_input_data[868 % IN_WIDTH] : pong_storage_data_594 ^ i_input_data[868 % IN_WIDTH];
                960 / IN_WIDTH: pong_storage_data_594 <= (fillup_transition == 1'b1) ? i_input_data[960 % IN_WIDTH] : pong_storage_data_594 ^ i_input_data[960 % IN_WIDTH];
                default: pong_storage_data_594 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_594;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_594 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_594;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_594 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_594;
            end
        end
    end
end

logic ping_storage_data_595;
logic pong_storage_data_595;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_595 <= 1'b0;
        pong_storage_data_595 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                212 / IN_WIDTH: ping_storage_data_595 <= (fillup_transition == 1'b1) ? i_input_data[212 % IN_WIDTH] : ping_storage_data_595 ^ i_input_data[212 % IN_WIDTH];
                350 / IN_WIDTH: ping_storage_data_595 <= (fillup_transition == 1'b1) ? i_input_data[350 % IN_WIDTH] : ping_storage_data_595 ^ i_input_data[350 % IN_WIDTH];
                869 / IN_WIDTH: ping_storage_data_595 <= (fillup_transition == 1'b1) ? i_input_data[869 % IN_WIDTH] : ping_storage_data_595 ^ i_input_data[869 % IN_WIDTH];
                961 / IN_WIDTH: ping_storage_data_595 <= (fillup_transition == 1'b1) ? i_input_data[961 % IN_WIDTH] : ping_storage_data_595 ^ i_input_data[961 % IN_WIDTH];
                default: ping_storage_data_595 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_595;
                endcase
            end else begin
                case (input_count)
                212 / IN_WIDTH: pong_storage_data_595 <= (fillup_transition == 1'b1) ? i_input_data[212 % IN_WIDTH] : pong_storage_data_595 ^ i_input_data[212 % IN_WIDTH];
                350 / IN_WIDTH: pong_storage_data_595 <= (fillup_transition == 1'b1) ? i_input_data[350 % IN_WIDTH] : pong_storage_data_595 ^ i_input_data[350 % IN_WIDTH];
                869 / IN_WIDTH: pong_storage_data_595 <= (fillup_transition == 1'b1) ? i_input_data[869 % IN_WIDTH] : pong_storage_data_595 ^ i_input_data[869 % IN_WIDTH];
                961 / IN_WIDTH: pong_storage_data_595 <= (fillup_transition == 1'b1) ? i_input_data[961 % IN_WIDTH] : pong_storage_data_595 ^ i_input_data[961 % IN_WIDTH];
                default: pong_storage_data_595 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_595;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_595 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_595;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_595 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_595;
            end
        end
    end
end

logic ping_storage_data_596;
logic pong_storage_data_596;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_596 <= 1'b0;
        pong_storage_data_596 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                213 / IN_WIDTH: ping_storage_data_596 <= (fillup_transition == 1'b1) ? i_input_data[213 % IN_WIDTH] : ping_storage_data_596 ^ i_input_data[213 % IN_WIDTH];
                351 / IN_WIDTH: ping_storage_data_596 <= (fillup_transition == 1'b1) ? i_input_data[351 % IN_WIDTH] : ping_storage_data_596 ^ i_input_data[351 % IN_WIDTH];
                870 / IN_WIDTH: ping_storage_data_596 <= (fillup_transition == 1'b1) ? i_input_data[870 % IN_WIDTH] : ping_storage_data_596 ^ i_input_data[870 % IN_WIDTH];
                962 / IN_WIDTH: ping_storage_data_596 <= (fillup_transition == 1'b1) ? i_input_data[962 % IN_WIDTH] : ping_storage_data_596 ^ i_input_data[962 % IN_WIDTH];
                default: ping_storage_data_596 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_596;
                endcase
            end else begin
                case (input_count)
                213 / IN_WIDTH: pong_storage_data_596 <= (fillup_transition == 1'b1) ? i_input_data[213 % IN_WIDTH] : pong_storage_data_596 ^ i_input_data[213 % IN_WIDTH];
                351 / IN_WIDTH: pong_storage_data_596 <= (fillup_transition == 1'b1) ? i_input_data[351 % IN_WIDTH] : pong_storage_data_596 ^ i_input_data[351 % IN_WIDTH];
                870 / IN_WIDTH: pong_storage_data_596 <= (fillup_transition == 1'b1) ? i_input_data[870 % IN_WIDTH] : pong_storage_data_596 ^ i_input_data[870 % IN_WIDTH];
                962 / IN_WIDTH: pong_storage_data_596 <= (fillup_transition == 1'b1) ? i_input_data[962 % IN_WIDTH] : pong_storage_data_596 ^ i_input_data[962 % IN_WIDTH];
                default: pong_storage_data_596 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_596;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_596 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_596;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_596 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_596;
            end
        end
    end
end

logic ping_storage_data_597;
logic pong_storage_data_597;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_597 <= 1'b0;
        pong_storage_data_597 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                214 / IN_WIDTH: ping_storage_data_597 <= (fillup_transition == 1'b1) ? i_input_data[214 % IN_WIDTH] : ping_storage_data_597 ^ i_input_data[214 % IN_WIDTH];
                352 / IN_WIDTH: ping_storage_data_597 <= (fillup_transition == 1'b1) ? i_input_data[352 % IN_WIDTH] : ping_storage_data_597 ^ i_input_data[352 % IN_WIDTH];
                871 / IN_WIDTH: ping_storage_data_597 <= (fillup_transition == 1'b1) ? i_input_data[871 % IN_WIDTH] : ping_storage_data_597 ^ i_input_data[871 % IN_WIDTH];
                963 / IN_WIDTH: ping_storage_data_597 <= (fillup_transition == 1'b1) ? i_input_data[963 % IN_WIDTH] : ping_storage_data_597 ^ i_input_data[963 % IN_WIDTH];
                default: ping_storage_data_597 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_597;
                endcase
            end else begin
                case (input_count)
                214 / IN_WIDTH: pong_storage_data_597 <= (fillup_transition == 1'b1) ? i_input_data[214 % IN_WIDTH] : pong_storage_data_597 ^ i_input_data[214 % IN_WIDTH];
                352 / IN_WIDTH: pong_storage_data_597 <= (fillup_transition == 1'b1) ? i_input_data[352 % IN_WIDTH] : pong_storage_data_597 ^ i_input_data[352 % IN_WIDTH];
                871 / IN_WIDTH: pong_storage_data_597 <= (fillup_transition == 1'b1) ? i_input_data[871 % IN_WIDTH] : pong_storage_data_597 ^ i_input_data[871 % IN_WIDTH];
                963 / IN_WIDTH: pong_storage_data_597 <= (fillup_transition == 1'b1) ? i_input_data[963 % IN_WIDTH] : pong_storage_data_597 ^ i_input_data[963 % IN_WIDTH];
                default: pong_storage_data_597 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_597;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_597 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_597;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_597 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_597;
            end
        end
    end
end

logic ping_storage_data_598;
logic pong_storage_data_598;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_598 <= 1'b0;
        pong_storage_data_598 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                215 / IN_WIDTH: ping_storage_data_598 <= (fillup_transition == 1'b1) ? i_input_data[215 % IN_WIDTH] : ping_storage_data_598 ^ i_input_data[215 % IN_WIDTH];
                353 / IN_WIDTH: ping_storage_data_598 <= (fillup_transition == 1'b1) ? i_input_data[353 % IN_WIDTH] : ping_storage_data_598 ^ i_input_data[353 % IN_WIDTH];
                872 / IN_WIDTH: ping_storage_data_598 <= (fillup_transition == 1'b1) ? i_input_data[872 % IN_WIDTH] : ping_storage_data_598 ^ i_input_data[872 % IN_WIDTH];
                964 / IN_WIDTH: ping_storage_data_598 <= (fillup_transition == 1'b1) ? i_input_data[964 % IN_WIDTH] : ping_storage_data_598 ^ i_input_data[964 % IN_WIDTH];
                default: ping_storage_data_598 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_598;
                endcase
            end else begin
                case (input_count)
                215 / IN_WIDTH: pong_storage_data_598 <= (fillup_transition == 1'b1) ? i_input_data[215 % IN_WIDTH] : pong_storage_data_598 ^ i_input_data[215 % IN_WIDTH];
                353 / IN_WIDTH: pong_storage_data_598 <= (fillup_transition == 1'b1) ? i_input_data[353 % IN_WIDTH] : pong_storage_data_598 ^ i_input_data[353 % IN_WIDTH];
                872 / IN_WIDTH: pong_storage_data_598 <= (fillup_transition == 1'b1) ? i_input_data[872 % IN_WIDTH] : pong_storage_data_598 ^ i_input_data[872 % IN_WIDTH];
                964 / IN_WIDTH: pong_storage_data_598 <= (fillup_transition == 1'b1) ? i_input_data[964 % IN_WIDTH] : pong_storage_data_598 ^ i_input_data[964 % IN_WIDTH];
                default: pong_storage_data_598 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_598;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_598 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_598;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_598 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_598;
            end
        end
    end
end

logic ping_storage_data_599;
logic pong_storage_data_599;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_599 <= 1'b0;
        pong_storage_data_599 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                216 / IN_WIDTH: ping_storage_data_599 <= (fillup_transition == 1'b1) ? i_input_data[216 % IN_WIDTH] : ping_storage_data_599 ^ i_input_data[216 % IN_WIDTH];
                354 / IN_WIDTH: ping_storage_data_599 <= (fillup_transition == 1'b1) ? i_input_data[354 % IN_WIDTH] : ping_storage_data_599 ^ i_input_data[354 % IN_WIDTH];
                873 / IN_WIDTH: ping_storage_data_599 <= (fillup_transition == 1'b1) ? i_input_data[873 % IN_WIDTH] : ping_storage_data_599 ^ i_input_data[873 % IN_WIDTH];
                965 / IN_WIDTH: ping_storage_data_599 <= (fillup_transition == 1'b1) ? i_input_data[965 % IN_WIDTH] : ping_storage_data_599 ^ i_input_data[965 % IN_WIDTH];
                default: ping_storage_data_599 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_599;
                endcase
            end else begin
                case (input_count)
                216 / IN_WIDTH: pong_storage_data_599 <= (fillup_transition == 1'b1) ? i_input_data[216 % IN_WIDTH] : pong_storage_data_599 ^ i_input_data[216 % IN_WIDTH];
                354 / IN_WIDTH: pong_storage_data_599 <= (fillup_transition == 1'b1) ? i_input_data[354 % IN_WIDTH] : pong_storage_data_599 ^ i_input_data[354 % IN_WIDTH];
                873 / IN_WIDTH: pong_storage_data_599 <= (fillup_transition == 1'b1) ? i_input_data[873 % IN_WIDTH] : pong_storage_data_599 ^ i_input_data[873 % IN_WIDTH];
                965 / IN_WIDTH: pong_storage_data_599 <= (fillup_transition == 1'b1) ? i_input_data[965 % IN_WIDTH] : pong_storage_data_599 ^ i_input_data[965 % IN_WIDTH];
                default: pong_storage_data_599 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_599;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_599 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_599;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_599 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_599;
            end
        end
    end
end

logic ping_storage_data_600;
logic pong_storage_data_600;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_600 <= 1'b0;
        pong_storage_data_600 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                217 / IN_WIDTH: ping_storage_data_600 <= (fillup_transition == 1'b1) ? i_input_data[217 % IN_WIDTH] : ping_storage_data_600 ^ i_input_data[217 % IN_WIDTH];
                355 / IN_WIDTH: ping_storage_data_600 <= (fillup_transition == 1'b1) ? i_input_data[355 % IN_WIDTH] : ping_storage_data_600 ^ i_input_data[355 % IN_WIDTH];
                874 / IN_WIDTH: ping_storage_data_600 <= (fillup_transition == 1'b1) ? i_input_data[874 % IN_WIDTH] : ping_storage_data_600 ^ i_input_data[874 % IN_WIDTH];
                966 / IN_WIDTH: ping_storage_data_600 <= (fillup_transition == 1'b1) ? i_input_data[966 % IN_WIDTH] : ping_storage_data_600 ^ i_input_data[966 % IN_WIDTH];
                default: ping_storage_data_600 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_600;
                endcase
            end else begin
                case (input_count)
                217 / IN_WIDTH: pong_storage_data_600 <= (fillup_transition == 1'b1) ? i_input_data[217 % IN_WIDTH] : pong_storage_data_600 ^ i_input_data[217 % IN_WIDTH];
                355 / IN_WIDTH: pong_storage_data_600 <= (fillup_transition == 1'b1) ? i_input_data[355 % IN_WIDTH] : pong_storage_data_600 ^ i_input_data[355 % IN_WIDTH];
                874 / IN_WIDTH: pong_storage_data_600 <= (fillup_transition == 1'b1) ? i_input_data[874 % IN_WIDTH] : pong_storage_data_600 ^ i_input_data[874 % IN_WIDTH];
                966 / IN_WIDTH: pong_storage_data_600 <= (fillup_transition == 1'b1) ? i_input_data[966 % IN_WIDTH] : pong_storage_data_600 ^ i_input_data[966 % IN_WIDTH];
                default: pong_storage_data_600 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_600;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_600 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_600;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_600 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_600;
            end
        end
    end
end

logic ping_storage_data_601;
logic pong_storage_data_601;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_601 <= 1'b0;
        pong_storage_data_601 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                218 / IN_WIDTH: ping_storage_data_601 <= (fillup_transition == 1'b1) ? i_input_data[218 % IN_WIDTH] : ping_storage_data_601 ^ i_input_data[218 % IN_WIDTH];
                356 / IN_WIDTH: ping_storage_data_601 <= (fillup_transition == 1'b1) ? i_input_data[356 % IN_WIDTH] : ping_storage_data_601 ^ i_input_data[356 % IN_WIDTH];
                875 / IN_WIDTH: ping_storage_data_601 <= (fillup_transition == 1'b1) ? i_input_data[875 % IN_WIDTH] : ping_storage_data_601 ^ i_input_data[875 % IN_WIDTH];
                967 / IN_WIDTH: ping_storage_data_601 <= (fillup_transition == 1'b1) ? i_input_data[967 % IN_WIDTH] : ping_storage_data_601 ^ i_input_data[967 % IN_WIDTH];
                default: ping_storage_data_601 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_601;
                endcase
            end else begin
                case (input_count)
                218 / IN_WIDTH: pong_storage_data_601 <= (fillup_transition == 1'b1) ? i_input_data[218 % IN_WIDTH] : pong_storage_data_601 ^ i_input_data[218 % IN_WIDTH];
                356 / IN_WIDTH: pong_storage_data_601 <= (fillup_transition == 1'b1) ? i_input_data[356 % IN_WIDTH] : pong_storage_data_601 ^ i_input_data[356 % IN_WIDTH];
                875 / IN_WIDTH: pong_storage_data_601 <= (fillup_transition == 1'b1) ? i_input_data[875 % IN_WIDTH] : pong_storage_data_601 ^ i_input_data[875 % IN_WIDTH];
                967 / IN_WIDTH: pong_storage_data_601 <= (fillup_transition == 1'b1) ? i_input_data[967 % IN_WIDTH] : pong_storage_data_601 ^ i_input_data[967 % IN_WIDTH];
                default: pong_storage_data_601 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_601;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_601 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_601;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_601 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_601;
            end
        end
    end
end

logic ping_storage_data_602;
logic pong_storage_data_602;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_602 <= 1'b0;
        pong_storage_data_602 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                219 / IN_WIDTH: ping_storage_data_602 <= (fillup_transition == 1'b1) ? i_input_data[219 % IN_WIDTH] : ping_storage_data_602 ^ i_input_data[219 % IN_WIDTH];
                357 / IN_WIDTH: ping_storage_data_602 <= (fillup_transition == 1'b1) ? i_input_data[357 % IN_WIDTH] : ping_storage_data_602 ^ i_input_data[357 % IN_WIDTH];
                876 / IN_WIDTH: ping_storage_data_602 <= (fillup_transition == 1'b1) ? i_input_data[876 % IN_WIDTH] : ping_storage_data_602 ^ i_input_data[876 % IN_WIDTH];
                968 / IN_WIDTH: ping_storage_data_602 <= (fillup_transition == 1'b1) ? i_input_data[968 % IN_WIDTH] : ping_storage_data_602 ^ i_input_data[968 % IN_WIDTH];
                default: ping_storage_data_602 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_602;
                endcase
            end else begin
                case (input_count)
                219 / IN_WIDTH: pong_storage_data_602 <= (fillup_transition == 1'b1) ? i_input_data[219 % IN_WIDTH] : pong_storage_data_602 ^ i_input_data[219 % IN_WIDTH];
                357 / IN_WIDTH: pong_storage_data_602 <= (fillup_transition == 1'b1) ? i_input_data[357 % IN_WIDTH] : pong_storage_data_602 ^ i_input_data[357 % IN_WIDTH];
                876 / IN_WIDTH: pong_storage_data_602 <= (fillup_transition == 1'b1) ? i_input_data[876 % IN_WIDTH] : pong_storage_data_602 ^ i_input_data[876 % IN_WIDTH];
                968 / IN_WIDTH: pong_storage_data_602 <= (fillup_transition == 1'b1) ? i_input_data[968 % IN_WIDTH] : pong_storage_data_602 ^ i_input_data[968 % IN_WIDTH];
                default: pong_storage_data_602 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_602;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_602 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_602;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_602 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_602;
            end
        end
    end
end

logic ping_storage_data_603;
logic pong_storage_data_603;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_603 <= 1'b0;
        pong_storage_data_603 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                220 / IN_WIDTH: ping_storage_data_603 <= (fillup_transition == 1'b1) ? i_input_data[220 % IN_WIDTH] : ping_storage_data_603 ^ i_input_data[220 % IN_WIDTH];
                358 / IN_WIDTH: ping_storage_data_603 <= (fillup_transition == 1'b1) ? i_input_data[358 % IN_WIDTH] : ping_storage_data_603 ^ i_input_data[358 % IN_WIDTH];
                877 / IN_WIDTH: ping_storage_data_603 <= (fillup_transition == 1'b1) ? i_input_data[877 % IN_WIDTH] : ping_storage_data_603 ^ i_input_data[877 % IN_WIDTH];
                969 / IN_WIDTH: ping_storage_data_603 <= (fillup_transition == 1'b1) ? i_input_data[969 % IN_WIDTH] : ping_storage_data_603 ^ i_input_data[969 % IN_WIDTH];
                default: ping_storage_data_603 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_603;
                endcase
            end else begin
                case (input_count)
                220 / IN_WIDTH: pong_storage_data_603 <= (fillup_transition == 1'b1) ? i_input_data[220 % IN_WIDTH] : pong_storage_data_603 ^ i_input_data[220 % IN_WIDTH];
                358 / IN_WIDTH: pong_storage_data_603 <= (fillup_transition == 1'b1) ? i_input_data[358 % IN_WIDTH] : pong_storage_data_603 ^ i_input_data[358 % IN_WIDTH];
                877 / IN_WIDTH: pong_storage_data_603 <= (fillup_transition == 1'b1) ? i_input_data[877 % IN_WIDTH] : pong_storage_data_603 ^ i_input_data[877 % IN_WIDTH];
                969 / IN_WIDTH: pong_storage_data_603 <= (fillup_transition == 1'b1) ? i_input_data[969 % IN_WIDTH] : pong_storage_data_603 ^ i_input_data[969 % IN_WIDTH];
                default: pong_storage_data_603 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_603;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_603 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_603;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_603 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_603;
            end
        end
    end
end

logic ping_storage_data_604;
logic pong_storage_data_604;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_604 <= 1'b0;
        pong_storage_data_604 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                221 / IN_WIDTH: ping_storage_data_604 <= (fillup_transition == 1'b1) ? i_input_data[221 % IN_WIDTH] : ping_storage_data_604 ^ i_input_data[221 % IN_WIDTH];
                359 / IN_WIDTH: ping_storage_data_604 <= (fillup_transition == 1'b1) ? i_input_data[359 % IN_WIDTH] : ping_storage_data_604 ^ i_input_data[359 % IN_WIDTH];
                878 / IN_WIDTH: ping_storage_data_604 <= (fillup_transition == 1'b1) ? i_input_data[878 % IN_WIDTH] : ping_storage_data_604 ^ i_input_data[878 % IN_WIDTH];
                970 / IN_WIDTH: ping_storage_data_604 <= (fillup_transition == 1'b1) ? i_input_data[970 % IN_WIDTH] : ping_storage_data_604 ^ i_input_data[970 % IN_WIDTH];
                default: ping_storage_data_604 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_604;
                endcase
            end else begin
                case (input_count)
                221 / IN_WIDTH: pong_storage_data_604 <= (fillup_transition == 1'b1) ? i_input_data[221 % IN_WIDTH] : pong_storage_data_604 ^ i_input_data[221 % IN_WIDTH];
                359 / IN_WIDTH: pong_storage_data_604 <= (fillup_transition == 1'b1) ? i_input_data[359 % IN_WIDTH] : pong_storage_data_604 ^ i_input_data[359 % IN_WIDTH];
                878 / IN_WIDTH: pong_storage_data_604 <= (fillup_transition == 1'b1) ? i_input_data[878 % IN_WIDTH] : pong_storage_data_604 ^ i_input_data[878 % IN_WIDTH];
                970 / IN_WIDTH: pong_storage_data_604 <= (fillup_transition == 1'b1) ? i_input_data[970 % IN_WIDTH] : pong_storage_data_604 ^ i_input_data[970 % IN_WIDTH];
                default: pong_storage_data_604 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_604;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_604 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_604;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_604 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_604;
            end
        end
    end
end

logic ping_storage_data_605;
logic pong_storage_data_605;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_605 <= 1'b0;
        pong_storage_data_605 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                222 / IN_WIDTH: ping_storage_data_605 <= (fillup_transition == 1'b1) ? i_input_data[222 % IN_WIDTH] : ping_storage_data_605 ^ i_input_data[222 % IN_WIDTH];
                360 / IN_WIDTH: ping_storage_data_605 <= (fillup_transition == 1'b1) ? i_input_data[360 % IN_WIDTH] : ping_storage_data_605 ^ i_input_data[360 % IN_WIDTH];
                879 / IN_WIDTH: ping_storage_data_605 <= (fillup_transition == 1'b1) ? i_input_data[879 % IN_WIDTH] : ping_storage_data_605 ^ i_input_data[879 % IN_WIDTH];
                971 / IN_WIDTH: ping_storage_data_605 <= (fillup_transition == 1'b1) ? i_input_data[971 % IN_WIDTH] : ping_storage_data_605 ^ i_input_data[971 % IN_WIDTH];
                default: ping_storage_data_605 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_605;
                endcase
            end else begin
                case (input_count)
                222 / IN_WIDTH: pong_storage_data_605 <= (fillup_transition == 1'b1) ? i_input_data[222 % IN_WIDTH] : pong_storage_data_605 ^ i_input_data[222 % IN_WIDTH];
                360 / IN_WIDTH: pong_storage_data_605 <= (fillup_transition == 1'b1) ? i_input_data[360 % IN_WIDTH] : pong_storage_data_605 ^ i_input_data[360 % IN_WIDTH];
                879 / IN_WIDTH: pong_storage_data_605 <= (fillup_transition == 1'b1) ? i_input_data[879 % IN_WIDTH] : pong_storage_data_605 ^ i_input_data[879 % IN_WIDTH];
                971 / IN_WIDTH: pong_storage_data_605 <= (fillup_transition == 1'b1) ? i_input_data[971 % IN_WIDTH] : pong_storage_data_605 ^ i_input_data[971 % IN_WIDTH];
                default: pong_storage_data_605 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_605;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_605 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_605;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_605 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_605;
            end
        end
    end
end

logic ping_storage_data_606;
logic pong_storage_data_606;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_606 <= 1'b0;
        pong_storage_data_606 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                223 / IN_WIDTH: ping_storage_data_606 <= (fillup_transition == 1'b1) ? i_input_data[223 % IN_WIDTH] : ping_storage_data_606 ^ i_input_data[223 % IN_WIDTH];
                361 / IN_WIDTH: ping_storage_data_606 <= (fillup_transition == 1'b1) ? i_input_data[361 % IN_WIDTH] : ping_storage_data_606 ^ i_input_data[361 % IN_WIDTH];
                880 / IN_WIDTH: ping_storage_data_606 <= (fillup_transition == 1'b1) ? i_input_data[880 % IN_WIDTH] : ping_storage_data_606 ^ i_input_data[880 % IN_WIDTH];
                972 / IN_WIDTH: ping_storage_data_606 <= (fillup_transition == 1'b1) ? i_input_data[972 % IN_WIDTH] : ping_storage_data_606 ^ i_input_data[972 % IN_WIDTH];
                default: ping_storage_data_606 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_606;
                endcase
            end else begin
                case (input_count)
                223 / IN_WIDTH: pong_storage_data_606 <= (fillup_transition == 1'b1) ? i_input_data[223 % IN_WIDTH] : pong_storage_data_606 ^ i_input_data[223 % IN_WIDTH];
                361 / IN_WIDTH: pong_storage_data_606 <= (fillup_transition == 1'b1) ? i_input_data[361 % IN_WIDTH] : pong_storage_data_606 ^ i_input_data[361 % IN_WIDTH];
                880 / IN_WIDTH: pong_storage_data_606 <= (fillup_transition == 1'b1) ? i_input_data[880 % IN_WIDTH] : pong_storage_data_606 ^ i_input_data[880 % IN_WIDTH];
                972 / IN_WIDTH: pong_storage_data_606 <= (fillup_transition == 1'b1) ? i_input_data[972 % IN_WIDTH] : pong_storage_data_606 ^ i_input_data[972 % IN_WIDTH];
                default: pong_storage_data_606 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_606;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_606 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_606;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_606 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_606;
            end
        end
    end
end

logic ping_storage_data_607;
logic pong_storage_data_607;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_607 <= 1'b0;
        pong_storage_data_607 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                224 / IN_WIDTH: ping_storage_data_607 <= (fillup_transition == 1'b1) ? i_input_data[224 % IN_WIDTH] : ping_storage_data_607 ^ i_input_data[224 % IN_WIDTH];
                362 / IN_WIDTH: ping_storage_data_607 <= (fillup_transition == 1'b1) ? i_input_data[362 % IN_WIDTH] : ping_storage_data_607 ^ i_input_data[362 % IN_WIDTH];
                881 / IN_WIDTH: ping_storage_data_607 <= (fillup_transition == 1'b1) ? i_input_data[881 % IN_WIDTH] : ping_storage_data_607 ^ i_input_data[881 % IN_WIDTH];
                973 / IN_WIDTH: ping_storage_data_607 <= (fillup_transition == 1'b1) ? i_input_data[973 % IN_WIDTH] : ping_storage_data_607 ^ i_input_data[973 % IN_WIDTH];
                default: ping_storage_data_607 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_607;
                endcase
            end else begin
                case (input_count)
                224 / IN_WIDTH: pong_storage_data_607 <= (fillup_transition == 1'b1) ? i_input_data[224 % IN_WIDTH] : pong_storage_data_607 ^ i_input_data[224 % IN_WIDTH];
                362 / IN_WIDTH: pong_storage_data_607 <= (fillup_transition == 1'b1) ? i_input_data[362 % IN_WIDTH] : pong_storage_data_607 ^ i_input_data[362 % IN_WIDTH];
                881 / IN_WIDTH: pong_storage_data_607 <= (fillup_transition == 1'b1) ? i_input_data[881 % IN_WIDTH] : pong_storage_data_607 ^ i_input_data[881 % IN_WIDTH];
                973 / IN_WIDTH: pong_storage_data_607 <= (fillup_transition == 1'b1) ? i_input_data[973 % IN_WIDTH] : pong_storage_data_607 ^ i_input_data[973 % IN_WIDTH];
                default: pong_storage_data_607 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_607;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_607 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_607;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_607 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_607;
            end
        end
    end
end

logic ping_storage_data_608;
logic pong_storage_data_608;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_608 <= 1'b0;
        pong_storage_data_608 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                225 / IN_WIDTH: ping_storage_data_608 <= (fillup_transition == 1'b1) ? i_input_data[225 % IN_WIDTH] : ping_storage_data_608 ^ i_input_data[225 % IN_WIDTH];
                363 / IN_WIDTH: ping_storage_data_608 <= (fillup_transition == 1'b1) ? i_input_data[363 % IN_WIDTH] : ping_storage_data_608 ^ i_input_data[363 % IN_WIDTH];
                882 / IN_WIDTH: ping_storage_data_608 <= (fillup_transition == 1'b1) ? i_input_data[882 % IN_WIDTH] : ping_storage_data_608 ^ i_input_data[882 % IN_WIDTH];
                974 / IN_WIDTH: ping_storage_data_608 <= (fillup_transition == 1'b1) ? i_input_data[974 % IN_WIDTH] : ping_storage_data_608 ^ i_input_data[974 % IN_WIDTH];
                default: ping_storage_data_608 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_608;
                endcase
            end else begin
                case (input_count)
                225 / IN_WIDTH: pong_storage_data_608 <= (fillup_transition == 1'b1) ? i_input_data[225 % IN_WIDTH] : pong_storage_data_608 ^ i_input_data[225 % IN_WIDTH];
                363 / IN_WIDTH: pong_storage_data_608 <= (fillup_transition == 1'b1) ? i_input_data[363 % IN_WIDTH] : pong_storage_data_608 ^ i_input_data[363 % IN_WIDTH];
                882 / IN_WIDTH: pong_storage_data_608 <= (fillup_transition == 1'b1) ? i_input_data[882 % IN_WIDTH] : pong_storage_data_608 ^ i_input_data[882 % IN_WIDTH];
                974 / IN_WIDTH: pong_storage_data_608 <= (fillup_transition == 1'b1) ? i_input_data[974 % IN_WIDTH] : pong_storage_data_608 ^ i_input_data[974 % IN_WIDTH];
                default: pong_storage_data_608 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_608;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_608 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_608;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_608 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_608;
            end
        end
    end
end

logic ping_storage_data_609;
logic pong_storage_data_609;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_609 <= 1'b0;
        pong_storage_data_609 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                226 / IN_WIDTH: ping_storage_data_609 <= (fillup_transition == 1'b1) ? i_input_data[226 % IN_WIDTH] : ping_storage_data_609 ^ i_input_data[226 % IN_WIDTH];
                364 / IN_WIDTH: ping_storage_data_609 <= (fillup_transition == 1'b1) ? i_input_data[364 % IN_WIDTH] : ping_storage_data_609 ^ i_input_data[364 % IN_WIDTH];
                883 / IN_WIDTH: ping_storage_data_609 <= (fillup_transition == 1'b1) ? i_input_data[883 % IN_WIDTH] : ping_storage_data_609 ^ i_input_data[883 % IN_WIDTH];
                975 / IN_WIDTH: ping_storage_data_609 <= (fillup_transition == 1'b1) ? i_input_data[975 % IN_WIDTH] : ping_storage_data_609 ^ i_input_data[975 % IN_WIDTH];
                default: ping_storage_data_609 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_609;
                endcase
            end else begin
                case (input_count)
                226 / IN_WIDTH: pong_storage_data_609 <= (fillup_transition == 1'b1) ? i_input_data[226 % IN_WIDTH] : pong_storage_data_609 ^ i_input_data[226 % IN_WIDTH];
                364 / IN_WIDTH: pong_storage_data_609 <= (fillup_transition == 1'b1) ? i_input_data[364 % IN_WIDTH] : pong_storage_data_609 ^ i_input_data[364 % IN_WIDTH];
                883 / IN_WIDTH: pong_storage_data_609 <= (fillup_transition == 1'b1) ? i_input_data[883 % IN_WIDTH] : pong_storage_data_609 ^ i_input_data[883 % IN_WIDTH];
                975 / IN_WIDTH: pong_storage_data_609 <= (fillup_transition == 1'b1) ? i_input_data[975 % IN_WIDTH] : pong_storage_data_609 ^ i_input_data[975 % IN_WIDTH];
                default: pong_storage_data_609 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_609;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_609 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_609;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_609 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_609;
            end
        end
    end
end

logic ping_storage_data_610;
logic pong_storage_data_610;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_610 <= 1'b0;
        pong_storage_data_610 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                227 / IN_WIDTH: ping_storage_data_610 <= (fillup_transition == 1'b1) ? i_input_data[227 % IN_WIDTH] : ping_storage_data_610 ^ i_input_data[227 % IN_WIDTH];
                365 / IN_WIDTH: ping_storage_data_610 <= (fillup_transition == 1'b1) ? i_input_data[365 % IN_WIDTH] : ping_storage_data_610 ^ i_input_data[365 % IN_WIDTH];
                884 / IN_WIDTH: ping_storage_data_610 <= (fillup_transition == 1'b1) ? i_input_data[884 % IN_WIDTH] : ping_storage_data_610 ^ i_input_data[884 % IN_WIDTH];
                976 / IN_WIDTH: ping_storage_data_610 <= (fillup_transition == 1'b1) ? i_input_data[976 % IN_WIDTH] : ping_storage_data_610 ^ i_input_data[976 % IN_WIDTH];
                default: ping_storage_data_610 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_610;
                endcase
            end else begin
                case (input_count)
                227 / IN_WIDTH: pong_storage_data_610 <= (fillup_transition == 1'b1) ? i_input_data[227 % IN_WIDTH] : pong_storage_data_610 ^ i_input_data[227 % IN_WIDTH];
                365 / IN_WIDTH: pong_storage_data_610 <= (fillup_transition == 1'b1) ? i_input_data[365 % IN_WIDTH] : pong_storage_data_610 ^ i_input_data[365 % IN_WIDTH];
                884 / IN_WIDTH: pong_storage_data_610 <= (fillup_transition == 1'b1) ? i_input_data[884 % IN_WIDTH] : pong_storage_data_610 ^ i_input_data[884 % IN_WIDTH];
                976 / IN_WIDTH: pong_storage_data_610 <= (fillup_transition == 1'b1) ? i_input_data[976 % IN_WIDTH] : pong_storage_data_610 ^ i_input_data[976 % IN_WIDTH];
                default: pong_storage_data_610 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_610;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_610 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_610;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_610 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_610;
            end
        end
    end
end

logic ping_storage_data_611;
logic pong_storage_data_611;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_611 <= 1'b0;
        pong_storage_data_611 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                228 / IN_WIDTH: ping_storage_data_611 <= (fillup_transition == 1'b1) ? i_input_data[228 % IN_WIDTH] : ping_storage_data_611 ^ i_input_data[228 % IN_WIDTH];
                366 / IN_WIDTH: ping_storage_data_611 <= (fillup_transition == 1'b1) ? i_input_data[366 % IN_WIDTH] : ping_storage_data_611 ^ i_input_data[366 % IN_WIDTH];
                885 / IN_WIDTH: ping_storage_data_611 <= (fillup_transition == 1'b1) ? i_input_data[885 % IN_WIDTH] : ping_storage_data_611 ^ i_input_data[885 % IN_WIDTH];
                977 / IN_WIDTH: ping_storage_data_611 <= (fillup_transition == 1'b1) ? i_input_data[977 % IN_WIDTH] : ping_storage_data_611 ^ i_input_data[977 % IN_WIDTH];
                default: ping_storage_data_611 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_611;
                endcase
            end else begin
                case (input_count)
                228 / IN_WIDTH: pong_storage_data_611 <= (fillup_transition == 1'b1) ? i_input_data[228 % IN_WIDTH] : pong_storage_data_611 ^ i_input_data[228 % IN_WIDTH];
                366 / IN_WIDTH: pong_storage_data_611 <= (fillup_transition == 1'b1) ? i_input_data[366 % IN_WIDTH] : pong_storage_data_611 ^ i_input_data[366 % IN_WIDTH];
                885 / IN_WIDTH: pong_storage_data_611 <= (fillup_transition == 1'b1) ? i_input_data[885 % IN_WIDTH] : pong_storage_data_611 ^ i_input_data[885 % IN_WIDTH];
                977 / IN_WIDTH: pong_storage_data_611 <= (fillup_transition == 1'b1) ? i_input_data[977 % IN_WIDTH] : pong_storage_data_611 ^ i_input_data[977 % IN_WIDTH];
                default: pong_storage_data_611 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_611;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_611 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_611;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_611 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_611;
            end
        end
    end
end

logic ping_storage_data_612;
logic pong_storage_data_612;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_612 <= 1'b0;
        pong_storage_data_612 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                229 / IN_WIDTH: ping_storage_data_612 <= (fillup_transition == 1'b1) ? i_input_data[229 % IN_WIDTH] : ping_storage_data_612 ^ i_input_data[229 % IN_WIDTH];
                367 / IN_WIDTH: ping_storage_data_612 <= (fillup_transition == 1'b1) ? i_input_data[367 % IN_WIDTH] : ping_storage_data_612 ^ i_input_data[367 % IN_WIDTH];
                886 / IN_WIDTH: ping_storage_data_612 <= (fillup_transition == 1'b1) ? i_input_data[886 % IN_WIDTH] : ping_storage_data_612 ^ i_input_data[886 % IN_WIDTH];
                978 / IN_WIDTH: ping_storage_data_612 <= (fillup_transition == 1'b1) ? i_input_data[978 % IN_WIDTH] : ping_storage_data_612 ^ i_input_data[978 % IN_WIDTH];
                default: ping_storage_data_612 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_612;
                endcase
            end else begin
                case (input_count)
                229 / IN_WIDTH: pong_storage_data_612 <= (fillup_transition == 1'b1) ? i_input_data[229 % IN_WIDTH] : pong_storage_data_612 ^ i_input_data[229 % IN_WIDTH];
                367 / IN_WIDTH: pong_storage_data_612 <= (fillup_transition == 1'b1) ? i_input_data[367 % IN_WIDTH] : pong_storage_data_612 ^ i_input_data[367 % IN_WIDTH];
                886 / IN_WIDTH: pong_storage_data_612 <= (fillup_transition == 1'b1) ? i_input_data[886 % IN_WIDTH] : pong_storage_data_612 ^ i_input_data[886 % IN_WIDTH];
                978 / IN_WIDTH: pong_storage_data_612 <= (fillup_transition == 1'b1) ? i_input_data[978 % IN_WIDTH] : pong_storage_data_612 ^ i_input_data[978 % IN_WIDTH];
                default: pong_storage_data_612 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_612;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_612 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_612;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_612 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_612;
            end
        end
    end
end

logic ping_storage_data_613;
logic pong_storage_data_613;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_613 <= 1'b0;
        pong_storage_data_613 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                230 / IN_WIDTH: ping_storage_data_613 <= (fillup_transition == 1'b1) ? i_input_data[230 % IN_WIDTH] : ping_storage_data_613 ^ i_input_data[230 % IN_WIDTH];
                368 / IN_WIDTH: ping_storage_data_613 <= (fillup_transition == 1'b1) ? i_input_data[368 % IN_WIDTH] : ping_storage_data_613 ^ i_input_data[368 % IN_WIDTH];
                887 / IN_WIDTH: ping_storage_data_613 <= (fillup_transition == 1'b1) ? i_input_data[887 % IN_WIDTH] : ping_storage_data_613 ^ i_input_data[887 % IN_WIDTH];
                979 / IN_WIDTH: ping_storage_data_613 <= (fillup_transition == 1'b1) ? i_input_data[979 % IN_WIDTH] : ping_storage_data_613 ^ i_input_data[979 % IN_WIDTH];
                default: ping_storage_data_613 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_613;
                endcase
            end else begin
                case (input_count)
                230 / IN_WIDTH: pong_storage_data_613 <= (fillup_transition == 1'b1) ? i_input_data[230 % IN_WIDTH] : pong_storage_data_613 ^ i_input_data[230 % IN_WIDTH];
                368 / IN_WIDTH: pong_storage_data_613 <= (fillup_transition == 1'b1) ? i_input_data[368 % IN_WIDTH] : pong_storage_data_613 ^ i_input_data[368 % IN_WIDTH];
                887 / IN_WIDTH: pong_storage_data_613 <= (fillup_transition == 1'b1) ? i_input_data[887 % IN_WIDTH] : pong_storage_data_613 ^ i_input_data[887 % IN_WIDTH];
                979 / IN_WIDTH: pong_storage_data_613 <= (fillup_transition == 1'b1) ? i_input_data[979 % IN_WIDTH] : pong_storage_data_613 ^ i_input_data[979 % IN_WIDTH];
                default: pong_storage_data_613 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_613;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_613 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_613;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_613 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_613;
            end
        end
    end
end

logic ping_storage_data_614;
logic pong_storage_data_614;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_614 <= 1'b0;
        pong_storage_data_614 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                231 / IN_WIDTH: ping_storage_data_614 <= (fillup_transition == 1'b1) ? i_input_data[231 % IN_WIDTH] : ping_storage_data_614 ^ i_input_data[231 % IN_WIDTH];
                369 / IN_WIDTH: ping_storage_data_614 <= (fillup_transition == 1'b1) ? i_input_data[369 % IN_WIDTH] : ping_storage_data_614 ^ i_input_data[369 % IN_WIDTH];
                888 / IN_WIDTH: ping_storage_data_614 <= (fillup_transition == 1'b1) ? i_input_data[888 % IN_WIDTH] : ping_storage_data_614 ^ i_input_data[888 % IN_WIDTH];
                980 / IN_WIDTH: ping_storage_data_614 <= (fillup_transition == 1'b1) ? i_input_data[980 % IN_WIDTH] : ping_storage_data_614 ^ i_input_data[980 % IN_WIDTH];
                default: ping_storage_data_614 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_614;
                endcase
            end else begin
                case (input_count)
                231 / IN_WIDTH: pong_storage_data_614 <= (fillup_transition == 1'b1) ? i_input_data[231 % IN_WIDTH] : pong_storage_data_614 ^ i_input_data[231 % IN_WIDTH];
                369 / IN_WIDTH: pong_storage_data_614 <= (fillup_transition == 1'b1) ? i_input_data[369 % IN_WIDTH] : pong_storage_data_614 ^ i_input_data[369 % IN_WIDTH];
                888 / IN_WIDTH: pong_storage_data_614 <= (fillup_transition == 1'b1) ? i_input_data[888 % IN_WIDTH] : pong_storage_data_614 ^ i_input_data[888 % IN_WIDTH];
                980 / IN_WIDTH: pong_storage_data_614 <= (fillup_transition == 1'b1) ? i_input_data[980 % IN_WIDTH] : pong_storage_data_614 ^ i_input_data[980 % IN_WIDTH];
                default: pong_storage_data_614 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_614;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_614 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_614;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_614 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_614;
            end
        end
    end
end

logic ping_storage_data_615;
logic pong_storage_data_615;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_615 <= 1'b0;
        pong_storage_data_615 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                232 / IN_WIDTH: ping_storage_data_615 <= (fillup_transition == 1'b1) ? i_input_data[232 % IN_WIDTH] : ping_storage_data_615 ^ i_input_data[232 % IN_WIDTH];
                370 / IN_WIDTH: ping_storage_data_615 <= (fillup_transition == 1'b1) ? i_input_data[370 % IN_WIDTH] : ping_storage_data_615 ^ i_input_data[370 % IN_WIDTH];
                889 / IN_WIDTH: ping_storage_data_615 <= (fillup_transition == 1'b1) ? i_input_data[889 % IN_WIDTH] : ping_storage_data_615 ^ i_input_data[889 % IN_WIDTH];
                981 / IN_WIDTH: ping_storage_data_615 <= (fillup_transition == 1'b1) ? i_input_data[981 % IN_WIDTH] : ping_storage_data_615 ^ i_input_data[981 % IN_WIDTH];
                default: ping_storage_data_615 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_615;
                endcase
            end else begin
                case (input_count)
                232 / IN_WIDTH: pong_storage_data_615 <= (fillup_transition == 1'b1) ? i_input_data[232 % IN_WIDTH] : pong_storage_data_615 ^ i_input_data[232 % IN_WIDTH];
                370 / IN_WIDTH: pong_storage_data_615 <= (fillup_transition == 1'b1) ? i_input_data[370 % IN_WIDTH] : pong_storage_data_615 ^ i_input_data[370 % IN_WIDTH];
                889 / IN_WIDTH: pong_storage_data_615 <= (fillup_transition == 1'b1) ? i_input_data[889 % IN_WIDTH] : pong_storage_data_615 ^ i_input_data[889 % IN_WIDTH];
                981 / IN_WIDTH: pong_storage_data_615 <= (fillup_transition == 1'b1) ? i_input_data[981 % IN_WIDTH] : pong_storage_data_615 ^ i_input_data[981 % IN_WIDTH];
                default: pong_storage_data_615 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_615;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_615 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_615;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_615 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_615;
            end
        end
    end
end

logic ping_storage_data_616;
logic pong_storage_data_616;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_616 <= 1'b0;
        pong_storage_data_616 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                233 / IN_WIDTH: ping_storage_data_616 <= (fillup_transition == 1'b1) ? i_input_data[233 % IN_WIDTH] : ping_storage_data_616 ^ i_input_data[233 % IN_WIDTH];
                371 / IN_WIDTH: ping_storage_data_616 <= (fillup_transition == 1'b1) ? i_input_data[371 % IN_WIDTH] : ping_storage_data_616 ^ i_input_data[371 % IN_WIDTH];
                890 / IN_WIDTH: ping_storage_data_616 <= (fillup_transition == 1'b1) ? i_input_data[890 % IN_WIDTH] : ping_storage_data_616 ^ i_input_data[890 % IN_WIDTH];
                982 / IN_WIDTH: ping_storage_data_616 <= (fillup_transition == 1'b1) ? i_input_data[982 % IN_WIDTH] : ping_storage_data_616 ^ i_input_data[982 % IN_WIDTH];
                default: ping_storage_data_616 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_616;
                endcase
            end else begin
                case (input_count)
                233 / IN_WIDTH: pong_storage_data_616 <= (fillup_transition == 1'b1) ? i_input_data[233 % IN_WIDTH] : pong_storage_data_616 ^ i_input_data[233 % IN_WIDTH];
                371 / IN_WIDTH: pong_storage_data_616 <= (fillup_transition == 1'b1) ? i_input_data[371 % IN_WIDTH] : pong_storage_data_616 ^ i_input_data[371 % IN_WIDTH];
                890 / IN_WIDTH: pong_storage_data_616 <= (fillup_transition == 1'b1) ? i_input_data[890 % IN_WIDTH] : pong_storage_data_616 ^ i_input_data[890 % IN_WIDTH];
                982 / IN_WIDTH: pong_storage_data_616 <= (fillup_transition == 1'b1) ? i_input_data[982 % IN_WIDTH] : pong_storage_data_616 ^ i_input_data[982 % IN_WIDTH];
                default: pong_storage_data_616 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_616;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_616 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_616;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_616 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_616;
            end
        end
    end
end

logic ping_storage_data_617;
logic pong_storage_data_617;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_617 <= 1'b0;
        pong_storage_data_617 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                234 / IN_WIDTH: ping_storage_data_617 <= (fillup_transition == 1'b1) ? i_input_data[234 % IN_WIDTH] : ping_storage_data_617 ^ i_input_data[234 % IN_WIDTH];
                372 / IN_WIDTH: ping_storage_data_617 <= (fillup_transition == 1'b1) ? i_input_data[372 % IN_WIDTH] : ping_storage_data_617 ^ i_input_data[372 % IN_WIDTH];
                891 / IN_WIDTH: ping_storage_data_617 <= (fillup_transition == 1'b1) ? i_input_data[891 % IN_WIDTH] : ping_storage_data_617 ^ i_input_data[891 % IN_WIDTH];
                983 / IN_WIDTH: ping_storage_data_617 <= (fillup_transition == 1'b1) ? i_input_data[983 % IN_WIDTH] : ping_storage_data_617 ^ i_input_data[983 % IN_WIDTH];
                default: ping_storage_data_617 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_617;
                endcase
            end else begin
                case (input_count)
                234 / IN_WIDTH: pong_storage_data_617 <= (fillup_transition == 1'b1) ? i_input_data[234 % IN_WIDTH] : pong_storage_data_617 ^ i_input_data[234 % IN_WIDTH];
                372 / IN_WIDTH: pong_storage_data_617 <= (fillup_transition == 1'b1) ? i_input_data[372 % IN_WIDTH] : pong_storage_data_617 ^ i_input_data[372 % IN_WIDTH];
                891 / IN_WIDTH: pong_storage_data_617 <= (fillup_transition == 1'b1) ? i_input_data[891 % IN_WIDTH] : pong_storage_data_617 ^ i_input_data[891 % IN_WIDTH];
                983 / IN_WIDTH: pong_storage_data_617 <= (fillup_transition == 1'b1) ? i_input_data[983 % IN_WIDTH] : pong_storage_data_617 ^ i_input_data[983 % IN_WIDTH];
                default: pong_storage_data_617 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_617;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_617 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_617;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_617 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_617;
            end
        end
    end
end

logic ping_storage_data_618;
logic pong_storage_data_618;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_618 <= 1'b0;
        pong_storage_data_618 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                235 / IN_WIDTH: ping_storage_data_618 <= (fillup_transition == 1'b1) ? i_input_data[235 % IN_WIDTH] : ping_storage_data_618 ^ i_input_data[235 % IN_WIDTH];
                373 / IN_WIDTH: ping_storage_data_618 <= (fillup_transition == 1'b1) ? i_input_data[373 % IN_WIDTH] : ping_storage_data_618 ^ i_input_data[373 % IN_WIDTH];
                892 / IN_WIDTH: ping_storage_data_618 <= (fillup_transition == 1'b1) ? i_input_data[892 % IN_WIDTH] : ping_storage_data_618 ^ i_input_data[892 % IN_WIDTH];
                984 / IN_WIDTH: ping_storage_data_618 <= (fillup_transition == 1'b1) ? i_input_data[984 % IN_WIDTH] : ping_storage_data_618 ^ i_input_data[984 % IN_WIDTH];
                default: ping_storage_data_618 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_618;
                endcase
            end else begin
                case (input_count)
                235 / IN_WIDTH: pong_storage_data_618 <= (fillup_transition == 1'b1) ? i_input_data[235 % IN_WIDTH] : pong_storage_data_618 ^ i_input_data[235 % IN_WIDTH];
                373 / IN_WIDTH: pong_storage_data_618 <= (fillup_transition == 1'b1) ? i_input_data[373 % IN_WIDTH] : pong_storage_data_618 ^ i_input_data[373 % IN_WIDTH];
                892 / IN_WIDTH: pong_storage_data_618 <= (fillup_transition == 1'b1) ? i_input_data[892 % IN_WIDTH] : pong_storage_data_618 ^ i_input_data[892 % IN_WIDTH];
                984 / IN_WIDTH: pong_storage_data_618 <= (fillup_transition == 1'b1) ? i_input_data[984 % IN_WIDTH] : pong_storage_data_618 ^ i_input_data[984 % IN_WIDTH];
                default: pong_storage_data_618 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_618;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_618 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_618;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_618 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_618;
            end
        end
    end
end

logic ping_storage_data_619;
logic pong_storage_data_619;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_619 <= 1'b0;
        pong_storage_data_619 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                236 / IN_WIDTH: ping_storage_data_619 <= (fillup_transition == 1'b1) ? i_input_data[236 % IN_WIDTH] : ping_storage_data_619 ^ i_input_data[236 % IN_WIDTH];
                374 / IN_WIDTH: ping_storage_data_619 <= (fillup_transition == 1'b1) ? i_input_data[374 % IN_WIDTH] : ping_storage_data_619 ^ i_input_data[374 % IN_WIDTH];
                893 / IN_WIDTH: ping_storage_data_619 <= (fillup_transition == 1'b1) ? i_input_data[893 % IN_WIDTH] : ping_storage_data_619 ^ i_input_data[893 % IN_WIDTH];
                985 / IN_WIDTH: ping_storage_data_619 <= (fillup_transition == 1'b1) ? i_input_data[985 % IN_WIDTH] : ping_storage_data_619 ^ i_input_data[985 % IN_WIDTH];
                default: ping_storage_data_619 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_619;
                endcase
            end else begin
                case (input_count)
                236 / IN_WIDTH: pong_storage_data_619 <= (fillup_transition == 1'b1) ? i_input_data[236 % IN_WIDTH] : pong_storage_data_619 ^ i_input_data[236 % IN_WIDTH];
                374 / IN_WIDTH: pong_storage_data_619 <= (fillup_transition == 1'b1) ? i_input_data[374 % IN_WIDTH] : pong_storage_data_619 ^ i_input_data[374 % IN_WIDTH];
                893 / IN_WIDTH: pong_storage_data_619 <= (fillup_transition == 1'b1) ? i_input_data[893 % IN_WIDTH] : pong_storage_data_619 ^ i_input_data[893 % IN_WIDTH];
                985 / IN_WIDTH: pong_storage_data_619 <= (fillup_transition == 1'b1) ? i_input_data[985 % IN_WIDTH] : pong_storage_data_619 ^ i_input_data[985 % IN_WIDTH];
                default: pong_storage_data_619 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_619;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_619 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_619;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_619 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_619;
            end
        end
    end
end

logic ping_storage_data_620;
logic pong_storage_data_620;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_620 <= 1'b0;
        pong_storage_data_620 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                237 / IN_WIDTH: ping_storage_data_620 <= (fillup_transition == 1'b1) ? i_input_data[237 % IN_WIDTH] : ping_storage_data_620 ^ i_input_data[237 % IN_WIDTH];
                375 / IN_WIDTH: ping_storage_data_620 <= (fillup_transition == 1'b1) ? i_input_data[375 % IN_WIDTH] : ping_storage_data_620 ^ i_input_data[375 % IN_WIDTH];
                894 / IN_WIDTH: ping_storage_data_620 <= (fillup_transition == 1'b1) ? i_input_data[894 % IN_WIDTH] : ping_storage_data_620 ^ i_input_data[894 % IN_WIDTH];
                986 / IN_WIDTH: ping_storage_data_620 <= (fillup_transition == 1'b1) ? i_input_data[986 % IN_WIDTH] : ping_storage_data_620 ^ i_input_data[986 % IN_WIDTH];
                default: ping_storage_data_620 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_620;
                endcase
            end else begin
                case (input_count)
                237 / IN_WIDTH: pong_storage_data_620 <= (fillup_transition == 1'b1) ? i_input_data[237 % IN_WIDTH] : pong_storage_data_620 ^ i_input_data[237 % IN_WIDTH];
                375 / IN_WIDTH: pong_storage_data_620 <= (fillup_transition == 1'b1) ? i_input_data[375 % IN_WIDTH] : pong_storage_data_620 ^ i_input_data[375 % IN_WIDTH];
                894 / IN_WIDTH: pong_storage_data_620 <= (fillup_transition == 1'b1) ? i_input_data[894 % IN_WIDTH] : pong_storage_data_620 ^ i_input_data[894 % IN_WIDTH];
                986 / IN_WIDTH: pong_storage_data_620 <= (fillup_transition == 1'b1) ? i_input_data[986 % IN_WIDTH] : pong_storage_data_620 ^ i_input_data[986 % IN_WIDTH];
                default: pong_storage_data_620 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_620;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_620 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_620;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_620 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_620;
            end
        end
    end
end

logic ping_storage_data_621;
logic pong_storage_data_621;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_621 <= 1'b0;
        pong_storage_data_621 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                238 / IN_WIDTH: ping_storage_data_621 <= (fillup_transition == 1'b1) ? i_input_data[238 % IN_WIDTH] : ping_storage_data_621 ^ i_input_data[238 % IN_WIDTH];
                376 / IN_WIDTH: ping_storage_data_621 <= (fillup_transition == 1'b1) ? i_input_data[376 % IN_WIDTH] : ping_storage_data_621 ^ i_input_data[376 % IN_WIDTH];
                895 / IN_WIDTH: ping_storage_data_621 <= (fillup_transition == 1'b1) ? i_input_data[895 % IN_WIDTH] : ping_storage_data_621 ^ i_input_data[895 % IN_WIDTH];
                987 / IN_WIDTH: ping_storage_data_621 <= (fillup_transition == 1'b1) ? i_input_data[987 % IN_WIDTH] : ping_storage_data_621 ^ i_input_data[987 % IN_WIDTH];
                default: ping_storage_data_621 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_621;
                endcase
            end else begin
                case (input_count)
                238 / IN_WIDTH: pong_storage_data_621 <= (fillup_transition == 1'b1) ? i_input_data[238 % IN_WIDTH] : pong_storage_data_621 ^ i_input_data[238 % IN_WIDTH];
                376 / IN_WIDTH: pong_storage_data_621 <= (fillup_transition == 1'b1) ? i_input_data[376 % IN_WIDTH] : pong_storage_data_621 ^ i_input_data[376 % IN_WIDTH];
                895 / IN_WIDTH: pong_storage_data_621 <= (fillup_transition == 1'b1) ? i_input_data[895 % IN_WIDTH] : pong_storage_data_621 ^ i_input_data[895 % IN_WIDTH];
                987 / IN_WIDTH: pong_storage_data_621 <= (fillup_transition == 1'b1) ? i_input_data[987 % IN_WIDTH] : pong_storage_data_621 ^ i_input_data[987 % IN_WIDTH];
                default: pong_storage_data_621 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_621;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_621 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_621;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_621 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_621;
            end
        end
    end
end

logic ping_storage_data_622;
logic pong_storage_data_622;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_622 <= 1'b0;
        pong_storage_data_622 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                239 / IN_WIDTH: ping_storage_data_622 <= (fillup_transition == 1'b1) ? i_input_data[239 % IN_WIDTH] : ping_storage_data_622 ^ i_input_data[239 % IN_WIDTH];
                377 / IN_WIDTH: ping_storage_data_622 <= (fillup_transition == 1'b1) ? i_input_data[377 % IN_WIDTH] : ping_storage_data_622 ^ i_input_data[377 % IN_WIDTH];
                896 / IN_WIDTH: ping_storage_data_622 <= (fillup_transition == 1'b1) ? i_input_data[896 % IN_WIDTH] : ping_storage_data_622 ^ i_input_data[896 % IN_WIDTH];
                988 / IN_WIDTH: ping_storage_data_622 <= (fillup_transition == 1'b1) ? i_input_data[988 % IN_WIDTH] : ping_storage_data_622 ^ i_input_data[988 % IN_WIDTH];
                default: ping_storage_data_622 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_622;
                endcase
            end else begin
                case (input_count)
                239 / IN_WIDTH: pong_storage_data_622 <= (fillup_transition == 1'b1) ? i_input_data[239 % IN_WIDTH] : pong_storage_data_622 ^ i_input_data[239 % IN_WIDTH];
                377 / IN_WIDTH: pong_storage_data_622 <= (fillup_transition == 1'b1) ? i_input_data[377 % IN_WIDTH] : pong_storage_data_622 ^ i_input_data[377 % IN_WIDTH];
                896 / IN_WIDTH: pong_storage_data_622 <= (fillup_transition == 1'b1) ? i_input_data[896 % IN_WIDTH] : pong_storage_data_622 ^ i_input_data[896 % IN_WIDTH];
                988 / IN_WIDTH: pong_storage_data_622 <= (fillup_transition == 1'b1) ? i_input_data[988 % IN_WIDTH] : pong_storage_data_622 ^ i_input_data[988 % IN_WIDTH];
                default: pong_storage_data_622 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_622;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_622 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_622;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_622 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_622;
            end
        end
    end
end

logic ping_storage_data_623;
logic pong_storage_data_623;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_623 <= 1'b0;
        pong_storage_data_623 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                240 / IN_WIDTH: ping_storage_data_623 <= (fillup_transition == 1'b1) ? i_input_data[240 % IN_WIDTH] : ping_storage_data_623 ^ i_input_data[240 % IN_WIDTH];
                378 / IN_WIDTH: ping_storage_data_623 <= (fillup_transition == 1'b1) ? i_input_data[378 % IN_WIDTH] : ping_storage_data_623 ^ i_input_data[378 % IN_WIDTH];
                897 / IN_WIDTH: ping_storage_data_623 <= (fillup_transition == 1'b1) ? i_input_data[897 % IN_WIDTH] : ping_storage_data_623 ^ i_input_data[897 % IN_WIDTH];
                989 / IN_WIDTH: ping_storage_data_623 <= (fillup_transition == 1'b1) ? i_input_data[989 % IN_WIDTH] : ping_storage_data_623 ^ i_input_data[989 % IN_WIDTH];
                default: ping_storage_data_623 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_623;
                endcase
            end else begin
                case (input_count)
                240 / IN_WIDTH: pong_storage_data_623 <= (fillup_transition == 1'b1) ? i_input_data[240 % IN_WIDTH] : pong_storage_data_623 ^ i_input_data[240 % IN_WIDTH];
                378 / IN_WIDTH: pong_storage_data_623 <= (fillup_transition == 1'b1) ? i_input_data[378 % IN_WIDTH] : pong_storage_data_623 ^ i_input_data[378 % IN_WIDTH];
                897 / IN_WIDTH: pong_storage_data_623 <= (fillup_transition == 1'b1) ? i_input_data[897 % IN_WIDTH] : pong_storage_data_623 ^ i_input_data[897 % IN_WIDTH];
                989 / IN_WIDTH: pong_storage_data_623 <= (fillup_transition == 1'b1) ? i_input_data[989 % IN_WIDTH] : pong_storage_data_623 ^ i_input_data[989 % IN_WIDTH];
                default: pong_storage_data_623 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_623;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_623 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_623;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_623 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_623;
            end
        end
    end
end

logic ping_storage_data_624;
logic pong_storage_data_624;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_624 <= 1'b0;
        pong_storage_data_624 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                241 / IN_WIDTH: ping_storage_data_624 <= (fillup_transition == 1'b1) ? i_input_data[241 % IN_WIDTH] : ping_storage_data_624 ^ i_input_data[241 % IN_WIDTH];
                379 / IN_WIDTH: ping_storage_data_624 <= (fillup_transition == 1'b1) ? i_input_data[379 % IN_WIDTH] : ping_storage_data_624 ^ i_input_data[379 % IN_WIDTH];
                898 / IN_WIDTH: ping_storage_data_624 <= (fillup_transition == 1'b1) ? i_input_data[898 % IN_WIDTH] : ping_storage_data_624 ^ i_input_data[898 % IN_WIDTH];
                990 / IN_WIDTH: ping_storage_data_624 <= (fillup_transition == 1'b1) ? i_input_data[990 % IN_WIDTH] : ping_storage_data_624 ^ i_input_data[990 % IN_WIDTH];
                default: ping_storage_data_624 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_624;
                endcase
            end else begin
                case (input_count)
                241 / IN_WIDTH: pong_storage_data_624 <= (fillup_transition == 1'b1) ? i_input_data[241 % IN_WIDTH] : pong_storage_data_624 ^ i_input_data[241 % IN_WIDTH];
                379 / IN_WIDTH: pong_storage_data_624 <= (fillup_transition == 1'b1) ? i_input_data[379 % IN_WIDTH] : pong_storage_data_624 ^ i_input_data[379 % IN_WIDTH];
                898 / IN_WIDTH: pong_storage_data_624 <= (fillup_transition == 1'b1) ? i_input_data[898 % IN_WIDTH] : pong_storage_data_624 ^ i_input_data[898 % IN_WIDTH];
                990 / IN_WIDTH: pong_storage_data_624 <= (fillup_transition == 1'b1) ? i_input_data[990 % IN_WIDTH] : pong_storage_data_624 ^ i_input_data[990 % IN_WIDTH];
                default: pong_storage_data_624 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_624;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_624 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_624;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_624 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_624;
            end
        end
    end
end

logic ping_storage_data_625;
logic pong_storage_data_625;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_625 <= 1'b0;
        pong_storage_data_625 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                242 / IN_WIDTH: ping_storage_data_625 <= (fillup_transition == 1'b1) ? i_input_data[242 % IN_WIDTH] : ping_storage_data_625 ^ i_input_data[242 % IN_WIDTH];
                380 / IN_WIDTH: ping_storage_data_625 <= (fillup_transition == 1'b1) ? i_input_data[380 % IN_WIDTH] : ping_storage_data_625 ^ i_input_data[380 % IN_WIDTH];
                899 / IN_WIDTH: ping_storage_data_625 <= (fillup_transition == 1'b1) ? i_input_data[899 % IN_WIDTH] : ping_storage_data_625 ^ i_input_data[899 % IN_WIDTH];
                991 / IN_WIDTH: ping_storage_data_625 <= (fillup_transition == 1'b1) ? i_input_data[991 % IN_WIDTH] : ping_storage_data_625 ^ i_input_data[991 % IN_WIDTH];
                default: ping_storage_data_625 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_625;
                endcase
            end else begin
                case (input_count)
                242 / IN_WIDTH: pong_storage_data_625 <= (fillup_transition == 1'b1) ? i_input_data[242 % IN_WIDTH] : pong_storage_data_625 ^ i_input_data[242 % IN_WIDTH];
                380 / IN_WIDTH: pong_storage_data_625 <= (fillup_transition == 1'b1) ? i_input_data[380 % IN_WIDTH] : pong_storage_data_625 ^ i_input_data[380 % IN_WIDTH];
                899 / IN_WIDTH: pong_storage_data_625 <= (fillup_transition == 1'b1) ? i_input_data[899 % IN_WIDTH] : pong_storage_data_625 ^ i_input_data[899 % IN_WIDTH];
                991 / IN_WIDTH: pong_storage_data_625 <= (fillup_transition == 1'b1) ? i_input_data[991 % IN_WIDTH] : pong_storage_data_625 ^ i_input_data[991 % IN_WIDTH];
                default: pong_storage_data_625 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_625;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_625 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_625;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_625 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_625;
            end
        end
    end
end

logic ping_storage_data_626;
logic pong_storage_data_626;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_626 <= 1'b0;
        pong_storage_data_626 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                243 / IN_WIDTH: ping_storage_data_626 <= (fillup_transition == 1'b1) ? i_input_data[243 % IN_WIDTH] : ping_storage_data_626 ^ i_input_data[243 % IN_WIDTH];
                381 / IN_WIDTH: ping_storage_data_626 <= (fillup_transition == 1'b1) ? i_input_data[381 % IN_WIDTH] : ping_storage_data_626 ^ i_input_data[381 % IN_WIDTH];
                900 / IN_WIDTH: ping_storage_data_626 <= (fillup_transition == 1'b1) ? i_input_data[900 % IN_WIDTH] : ping_storage_data_626 ^ i_input_data[900 % IN_WIDTH];
                992 / IN_WIDTH: ping_storage_data_626 <= (fillup_transition == 1'b1) ? i_input_data[992 % IN_WIDTH] : ping_storage_data_626 ^ i_input_data[992 % IN_WIDTH];
                default: ping_storage_data_626 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_626;
                endcase
            end else begin
                case (input_count)
                243 / IN_WIDTH: pong_storage_data_626 <= (fillup_transition == 1'b1) ? i_input_data[243 % IN_WIDTH] : pong_storage_data_626 ^ i_input_data[243 % IN_WIDTH];
                381 / IN_WIDTH: pong_storage_data_626 <= (fillup_transition == 1'b1) ? i_input_data[381 % IN_WIDTH] : pong_storage_data_626 ^ i_input_data[381 % IN_WIDTH];
                900 / IN_WIDTH: pong_storage_data_626 <= (fillup_transition == 1'b1) ? i_input_data[900 % IN_WIDTH] : pong_storage_data_626 ^ i_input_data[900 % IN_WIDTH];
                992 / IN_WIDTH: pong_storage_data_626 <= (fillup_transition == 1'b1) ? i_input_data[992 % IN_WIDTH] : pong_storage_data_626 ^ i_input_data[992 % IN_WIDTH];
                default: pong_storage_data_626 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_626;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_626 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_626;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_626 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_626;
            end
        end
    end
end

logic ping_storage_data_627;
logic pong_storage_data_627;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_627 <= 1'b0;
        pong_storage_data_627 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                244 / IN_WIDTH: ping_storage_data_627 <= (fillup_transition == 1'b1) ? i_input_data[244 % IN_WIDTH] : ping_storage_data_627 ^ i_input_data[244 % IN_WIDTH];
                382 / IN_WIDTH: ping_storage_data_627 <= (fillup_transition == 1'b1) ? i_input_data[382 % IN_WIDTH] : ping_storage_data_627 ^ i_input_data[382 % IN_WIDTH];
                901 / IN_WIDTH: ping_storage_data_627 <= (fillup_transition == 1'b1) ? i_input_data[901 % IN_WIDTH] : ping_storage_data_627 ^ i_input_data[901 % IN_WIDTH];
                993 / IN_WIDTH: ping_storage_data_627 <= (fillup_transition == 1'b1) ? i_input_data[993 % IN_WIDTH] : ping_storage_data_627 ^ i_input_data[993 % IN_WIDTH];
                default: ping_storage_data_627 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_627;
                endcase
            end else begin
                case (input_count)
                244 / IN_WIDTH: pong_storage_data_627 <= (fillup_transition == 1'b1) ? i_input_data[244 % IN_WIDTH] : pong_storage_data_627 ^ i_input_data[244 % IN_WIDTH];
                382 / IN_WIDTH: pong_storage_data_627 <= (fillup_transition == 1'b1) ? i_input_data[382 % IN_WIDTH] : pong_storage_data_627 ^ i_input_data[382 % IN_WIDTH];
                901 / IN_WIDTH: pong_storage_data_627 <= (fillup_transition == 1'b1) ? i_input_data[901 % IN_WIDTH] : pong_storage_data_627 ^ i_input_data[901 % IN_WIDTH];
                993 / IN_WIDTH: pong_storage_data_627 <= (fillup_transition == 1'b1) ? i_input_data[993 % IN_WIDTH] : pong_storage_data_627 ^ i_input_data[993 % IN_WIDTH];
                default: pong_storage_data_627 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_627;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_627 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_627;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_627 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_627;
            end
        end
    end
end

logic ping_storage_data_628;
logic pong_storage_data_628;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_628 <= 1'b0;
        pong_storage_data_628 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                245 / IN_WIDTH: ping_storage_data_628 <= (fillup_transition == 1'b1) ? i_input_data[245 % IN_WIDTH] : ping_storage_data_628 ^ i_input_data[245 % IN_WIDTH];
                383 / IN_WIDTH: ping_storage_data_628 <= (fillup_transition == 1'b1) ? i_input_data[383 % IN_WIDTH] : ping_storage_data_628 ^ i_input_data[383 % IN_WIDTH];
                902 / IN_WIDTH: ping_storage_data_628 <= (fillup_transition == 1'b1) ? i_input_data[902 % IN_WIDTH] : ping_storage_data_628 ^ i_input_data[902 % IN_WIDTH];
                994 / IN_WIDTH: ping_storage_data_628 <= (fillup_transition == 1'b1) ? i_input_data[994 % IN_WIDTH] : ping_storage_data_628 ^ i_input_data[994 % IN_WIDTH];
                default: ping_storage_data_628 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_628;
                endcase
            end else begin
                case (input_count)
                245 / IN_WIDTH: pong_storage_data_628 <= (fillup_transition == 1'b1) ? i_input_data[245 % IN_WIDTH] : pong_storage_data_628 ^ i_input_data[245 % IN_WIDTH];
                383 / IN_WIDTH: pong_storage_data_628 <= (fillup_transition == 1'b1) ? i_input_data[383 % IN_WIDTH] : pong_storage_data_628 ^ i_input_data[383 % IN_WIDTH];
                902 / IN_WIDTH: pong_storage_data_628 <= (fillup_transition == 1'b1) ? i_input_data[902 % IN_WIDTH] : pong_storage_data_628 ^ i_input_data[902 % IN_WIDTH];
                994 / IN_WIDTH: pong_storage_data_628 <= (fillup_transition == 1'b1) ? i_input_data[994 % IN_WIDTH] : pong_storage_data_628 ^ i_input_data[994 % IN_WIDTH];
                default: pong_storage_data_628 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_628;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_628 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_628;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_628 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_628;
            end
        end
    end
end

logic ping_storage_data_629;
logic pong_storage_data_629;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_629 <= 1'b0;
        pong_storage_data_629 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                246 / IN_WIDTH: ping_storage_data_629 <= (fillup_transition == 1'b1) ? i_input_data[246 % IN_WIDTH] : ping_storage_data_629 ^ i_input_data[246 % IN_WIDTH];
                288 / IN_WIDTH: ping_storage_data_629 <= (fillup_transition == 1'b1) ? i_input_data[288 % IN_WIDTH] : ping_storage_data_629 ^ i_input_data[288 % IN_WIDTH];
                903 / IN_WIDTH: ping_storage_data_629 <= (fillup_transition == 1'b1) ? i_input_data[903 % IN_WIDTH] : ping_storage_data_629 ^ i_input_data[903 % IN_WIDTH];
                995 / IN_WIDTH: ping_storage_data_629 <= (fillup_transition == 1'b1) ? i_input_data[995 % IN_WIDTH] : ping_storage_data_629 ^ i_input_data[995 % IN_WIDTH];
                default: ping_storage_data_629 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_629;
                endcase
            end else begin
                case (input_count)
                246 / IN_WIDTH: pong_storage_data_629 <= (fillup_transition == 1'b1) ? i_input_data[246 % IN_WIDTH] : pong_storage_data_629 ^ i_input_data[246 % IN_WIDTH];
                288 / IN_WIDTH: pong_storage_data_629 <= (fillup_transition == 1'b1) ? i_input_data[288 % IN_WIDTH] : pong_storage_data_629 ^ i_input_data[288 % IN_WIDTH];
                903 / IN_WIDTH: pong_storage_data_629 <= (fillup_transition == 1'b1) ? i_input_data[903 % IN_WIDTH] : pong_storage_data_629 ^ i_input_data[903 % IN_WIDTH];
                995 / IN_WIDTH: pong_storage_data_629 <= (fillup_transition == 1'b1) ? i_input_data[995 % IN_WIDTH] : pong_storage_data_629 ^ i_input_data[995 % IN_WIDTH];
                default: pong_storage_data_629 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_629;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_629 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_629;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_629 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_629;
            end
        end
    end
end

logic ping_storage_data_630;
logic pong_storage_data_630;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_630 <= 1'b0;
        pong_storage_data_630 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                247 / IN_WIDTH: ping_storage_data_630 <= (fillup_transition == 1'b1) ? i_input_data[247 % IN_WIDTH] : ping_storage_data_630 ^ i_input_data[247 % IN_WIDTH];
                289 / IN_WIDTH: ping_storage_data_630 <= (fillup_transition == 1'b1) ? i_input_data[289 % IN_WIDTH] : ping_storage_data_630 ^ i_input_data[289 % IN_WIDTH];
                904 / IN_WIDTH: ping_storage_data_630 <= (fillup_transition == 1'b1) ? i_input_data[904 % IN_WIDTH] : ping_storage_data_630 ^ i_input_data[904 % IN_WIDTH];
                996 / IN_WIDTH: ping_storage_data_630 <= (fillup_transition == 1'b1) ? i_input_data[996 % IN_WIDTH] : ping_storage_data_630 ^ i_input_data[996 % IN_WIDTH];
                default: ping_storage_data_630 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_630;
                endcase
            end else begin
                case (input_count)
                247 / IN_WIDTH: pong_storage_data_630 <= (fillup_transition == 1'b1) ? i_input_data[247 % IN_WIDTH] : pong_storage_data_630 ^ i_input_data[247 % IN_WIDTH];
                289 / IN_WIDTH: pong_storage_data_630 <= (fillup_transition == 1'b1) ? i_input_data[289 % IN_WIDTH] : pong_storage_data_630 ^ i_input_data[289 % IN_WIDTH];
                904 / IN_WIDTH: pong_storage_data_630 <= (fillup_transition == 1'b1) ? i_input_data[904 % IN_WIDTH] : pong_storage_data_630 ^ i_input_data[904 % IN_WIDTH];
                996 / IN_WIDTH: pong_storage_data_630 <= (fillup_transition == 1'b1) ? i_input_data[996 % IN_WIDTH] : pong_storage_data_630 ^ i_input_data[996 % IN_WIDTH];
                default: pong_storage_data_630 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_630;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_630 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_630;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_630 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_630;
            end
        end
    end
end

logic ping_storage_data_631;
logic pong_storage_data_631;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_631 <= 1'b0;
        pong_storage_data_631 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                248 / IN_WIDTH: ping_storage_data_631 <= (fillup_transition == 1'b1) ? i_input_data[248 % IN_WIDTH] : ping_storage_data_631 ^ i_input_data[248 % IN_WIDTH];
                290 / IN_WIDTH: ping_storage_data_631 <= (fillup_transition == 1'b1) ? i_input_data[290 % IN_WIDTH] : ping_storage_data_631 ^ i_input_data[290 % IN_WIDTH];
                905 / IN_WIDTH: ping_storage_data_631 <= (fillup_transition == 1'b1) ? i_input_data[905 % IN_WIDTH] : ping_storage_data_631 ^ i_input_data[905 % IN_WIDTH];
                997 / IN_WIDTH: ping_storage_data_631 <= (fillup_transition == 1'b1) ? i_input_data[997 % IN_WIDTH] : ping_storage_data_631 ^ i_input_data[997 % IN_WIDTH];
                default: ping_storage_data_631 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_631;
                endcase
            end else begin
                case (input_count)
                248 / IN_WIDTH: pong_storage_data_631 <= (fillup_transition == 1'b1) ? i_input_data[248 % IN_WIDTH] : pong_storage_data_631 ^ i_input_data[248 % IN_WIDTH];
                290 / IN_WIDTH: pong_storage_data_631 <= (fillup_transition == 1'b1) ? i_input_data[290 % IN_WIDTH] : pong_storage_data_631 ^ i_input_data[290 % IN_WIDTH];
                905 / IN_WIDTH: pong_storage_data_631 <= (fillup_transition == 1'b1) ? i_input_data[905 % IN_WIDTH] : pong_storage_data_631 ^ i_input_data[905 % IN_WIDTH];
                997 / IN_WIDTH: pong_storage_data_631 <= (fillup_transition == 1'b1) ? i_input_data[997 % IN_WIDTH] : pong_storage_data_631 ^ i_input_data[997 % IN_WIDTH];
                default: pong_storage_data_631 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_631;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_631 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_631;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_631 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_631;
            end
        end
    end
end

logic ping_storage_data_632;
logic pong_storage_data_632;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_632 <= 1'b0;
        pong_storage_data_632 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                249 / IN_WIDTH: ping_storage_data_632 <= (fillup_transition == 1'b1) ? i_input_data[249 % IN_WIDTH] : ping_storage_data_632 ^ i_input_data[249 % IN_WIDTH];
                291 / IN_WIDTH: ping_storage_data_632 <= (fillup_transition == 1'b1) ? i_input_data[291 % IN_WIDTH] : ping_storage_data_632 ^ i_input_data[291 % IN_WIDTH];
                906 / IN_WIDTH: ping_storage_data_632 <= (fillup_transition == 1'b1) ? i_input_data[906 % IN_WIDTH] : ping_storage_data_632 ^ i_input_data[906 % IN_WIDTH];
                998 / IN_WIDTH: ping_storage_data_632 <= (fillup_transition == 1'b1) ? i_input_data[998 % IN_WIDTH] : ping_storage_data_632 ^ i_input_data[998 % IN_WIDTH];
                default: ping_storage_data_632 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_632;
                endcase
            end else begin
                case (input_count)
                249 / IN_WIDTH: pong_storage_data_632 <= (fillup_transition == 1'b1) ? i_input_data[249 % IN_WIDTH] : pong_storage_data_632 ^ i_input_data[249 % IN_WIDTH];
                291 / IN_WIDTH: pong_storage_data_632 <= (fillup_transition == 1'b1) ? i_input_data[291 % IN_WIDTH] : pong_storage_data_632 ^ i_input_data[291 % IN_WIDTH];
                906 / IN_WIDTH: pong_storage_data_632 <= (fillup_transition == 1'b1) ? i_input_data[906 % IN_WIDTH] : pong_storage_data_632 ^ i_input_data[906 % IN_WIDTH];
                998 / IN_WIDTH: pong_storage_data_632 <= (fillup_transition == 1'b1) ? i_input_data[998 % IN_WIDTH] : pong_storage_data_632 ^ i_input_data[998 % IN_WIDTH];
                default: pong_storage_data_632 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_632;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_632 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_632;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_632 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_632;
            end
        end
    end
end

logic ping_storage_data_633;
logic pong_storage_data_633;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_633 <= 1'b0;
        pong_storage_data_633 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                250 / IN_WIDTH: ping_storage_data_633 <= (fillup_transition == 1'b1) ? i_input_data[250 % IN_WIDTH] : ping_storage_data_633 ^ i_input_data[250 % IN_WIDTH];
                292 / IN_WIDTH: ping_storage_data_633 <= (fillup_transition == 1'b1) ? i_input_data[292 % IN_WIDTH] : ping_storage_data_633 ^ i_input_data[292 % IN_WIDTH];
                907 / IN_WIDTH: ping_storage_data_633 <= (fillup_transition == 1'b1) ? i_input_data[907 % IN_WIDTH] : ping_storage_data_633 ^ i_input_data[907 % IN_WIDTH];
                999 / IN_WIDTH: ping_storage_data_633 <= (fillup_transition == 1'b1) ? i_input_data[999 % IN_WIDTH] : ping_storage_data_633 ^ i_input_data[999 % IN_WIDTH];
                default: ping_storage_data_633 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_633;
                endcase
            end else begin
                case (input_count)
                250 / IN_WIDTH: pong_storage_data_633 <= (fillup_transition == 1'b1) ? i_input_data[250 % IN_WIDTH] : pong_storage_data_633 ^ i_input_data[250 % IN_WIDTH];
                292 / IN_WIDTH: pong_storage_data_633 <= (fillup_transition == 1'b1) ? i_input_data[292 % IN_WIDTH] : pong_storage_data_633 ^ i_input_data[292 % IN_WIDTH];
                907 / IN_WIDTH: pong_storage_data_633 <= (fillup_transition == 1'b1) ? i_input_data[907 % IN_WIDTH] : pong_storage_data_633 ^ i_input_data[907 % IN_WIDTH];
                999 / IN_WIDTH: pong_storage_data_633 <= (fillup_transition == 1'b1) ? i_input_data[999 % IN_WIDTH] : pong_storage_data_633 ^ i_input_data[999 % IN_WIDTH];
                default: pong_storage_data_633 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_633;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_633 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_633;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_633 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_633;
            end
        end
    end
end

logic ping_storage_data_634;
logic pong_storage_data_634;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_634 <= 1'b0;
        pong_storage_data_634 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                251 / IN_WIDTH: ping_storage_data_634 <= (fillup_transition == 1'b1) ? i_input_data[251 % IN_WIDTH] : ping_storage_data_634 ^ i_input_data[251 % IN_WIDTH];
                293 / IN_WIDTH: ping_storage_data_634 <= (fillup_transition == 1'b1) ? i_input_data[293 % IN_WIDTH] : ping_storage_data_634 ^ i_input_data[293 % IN_WIDTH];
                908 / IN_WIDTH: ping_storage_data_634 <= (fillup_transition == 1'b1) ? i_input_data[908 % IN_WIDTH] : ping_storage_data_634 ^ i_input_data[908 % IN_WIDTH];
                1000 / IN_WIDTH: ping_storage_data_634 <= (fillup_transition == 1'b1) ? i_input_data[1000 % IN_WIDTH] : ping_storage_data_634 ^ i_input_data[1000 % IN_WIDTH];
                default: ping_storage_data_634 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_634;
                endcase
            end else begin
                case (input_count)
                251 / IN_WIDTH: pong_storage_data_634 <= (fillup_transition == 1'b1) ? i_input_data[251 % IN_WIDTH] : pong_storage_data_634 ^ i_input_data[251 % IN_WIDTH];
                293 / IN_WIDTH: pong_storage_data_634 <= (fillup_transition == 1'b1) ? i_input_data[293 % IN_WIDTH] : pong_storage_data_634 ^ i_input_data[293 % IN_WIDTH];
                908 / IN_WIDTH: pong_storage_data_634 <= (fillup_transition == 1'b1) ? i_input_data[908 % IN_WIDTH] : pong_storage_data_634 ^ i_input_data[908 % IN_WIDTH];
                1000 / IN_WIDTH: pong_storage_data_634 <= (fillup_transition == 1'b1) ? i_input_data[1000 % IN_WIDTH] : pong_storage_data_634 ^ i_input_data[1000 % IN_WIDTH];
                default: pong_storage_data_634 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_634;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_634 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_634;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_634 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_634;
            end
        end
    end
end

logic ping_storage_data_635;
logic pong_storage_data_635;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_635 <= 1'b0;
        pong_storage_data_635 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                252 / IN_WIDTH: ping_storage_data_635 <= (fillup_transition == 1'b1) ? i_input_data[252 % IN_WIDTH] : ping_storage_data_635 ^ i_input_data[252 % IN_WIDTH];
                294 / IN_WIDTH: ping_storage_data_635 <= (fillup_transition == 1'b1) ? i_input_data[294 % IN_WIDTH] : ping_storage_data_635 ^ i_input_data[294 % IN_WIDTH];
                909 / IN_WIDTH: ping_storage_data_635 <= (fillup_transition == 1'b1) ? i_input_data[909 % IN_WIDTH] : ping_storage_data_635 ^ i_input_data[909 % IN_WIDTH];
                1001 / IN_WIDTH: ping_storage_data_635 <= (fillup_transition == 1'b1) ? i_input_data[1001 % IN_WIDTH] : ping_storage_data_635 ^ i_input_data[1001 % IN_WIDTH];
                default: ping_storage_data_635 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_635;
                endcase
            end else begin
                case (input_count)
                252 / IN_WIDTH: pong_storage_data_635 <= (fillup_transition == 1'b1) ? i_input_data[252 % IN_WIDTH] : pong_storage_data_635 ^ i_input_data[252 % IN_WIDTH];
                294 / IN_WIDTH: pong_storage_data_635 <= (fillup_transition == 1'b1) ? i_input_data[294 % IN_WIDTH] : pong_storage_data_635 ^ i_input_data[294 % IN_WIDTH];
                909 / IN_WIDTH: pong_storage_data_635 <= (fillup_transition == 1'b1) ? i_input_data[909 % IN_WIDTH] : pong_storage_data_635 ^ i_input_data[909 % IN_WIDTH];
                1001 / IN_WIDTH: pong_storage_data_635 <= (fillup_transition == 1'b1) ? i_input_data[1001 % IN_WIDTH] : pong_storage_data_635 ^ i_input_data[1001 % IN_WIDTH];
                default: pong_storage_data_635 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_635;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_635 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_635;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_635 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_635;
            end
        end
    end
end

logic ping_storage_data_636;
logic pong_storage_data_636;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_636 <= 1'b0;
        pong_storage_data_636 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                253 / IN_WIDTH: ping_storage_data_636 <= (fillup_transition == 1'b1) ? i_input_data[253 % IN_WIDTH] : ping_storage_data_636 ^ i_input_data[253 % IN_WIDTH];
                295 / IN_WIDTH: ping_storage_data_636 <= (fillup_transition == 1'b1) ? i_input_data[295 % IN_WIDTH] : ping_storage_data_636 ^ i_input_data[295 % IN_WIDTH];
                910 / IN_WIDTH: ping_storage_data_636 <= (fillup_transition == 1'b1) ? i_input_data[910 % IN_WIDTH] : ping_storage_data_636 ^ i_input_data[910 % IN_WIDTH];
                1002 / IN_WIDTH: ping_storage_data_636 <= (fillup_transition == 1'b1) ? i_input_data[1002 % IN_WIDTH] : ping_storage_data_636 ^ i_input_data[1002 % IN_WIDTH];
                default: ping_storage_data_636 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_636;
                endcase
            end else begin
                case (input_count)
                253 / IN_WIDTH: pong_storage_data_636 <= (fillup_transition == 1'b1) ? i_input_data[253 % IN_WIDTH] : pong_storage_data_636 ^ i_input_data[253 % IN_WIDTH];
                295 / IN_WIDTH: pong_storage_data_636 <= (fillup_transition == 1'b1) ? i_input_data[295 % IN_WIDTH] : pong_storage_data_636 ^ i_input_data[295 % IN_WIDTH];
                910 / IN_WIDTH: pong_storage_data_636 <= (fillup_transition == 1'b1) ? i_input_data[910 % IN_WIDTH] : pong_storage_data_636 ^ i_input_data[910 % IN_WIDTH];
                1002 / IN_WIDTH: pong_storage_data_636 <= (fillup_transition == 1'b1) ? i_input_data[1002 % IN_WIDTH] : pong_storage_data_636 ^ i_input_data[1002 % IN_WIDTH];
                default: pong_storage_data_636 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_636;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_636 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_636;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_636 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_636;
            end
        end
    end
end

logic ping_storage_data_637;
logic pong_storage_data_637;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_637 <= 1'b0;
        pong_storage_data_637 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                254 / IN_WIDTH: ping_storage_data_637 <= (fillup_transition == 1'b1) ? i_input_data[254 % IN_WIDTH] : ping_storage_data_637 ^ i_input_data[254 % IN_WIDTH];
                296 / IN_WIDTH: ping_storage_data_637 <= (fillup_transition == 1'b1) ? i_input_data[296 % IN_WIDTH] : ping_storage_data_637 ^ i_input_data[296 % IN_WIDTH];
                911 / IN_WIDTH: ping_storage_data_637 <= (fillup_transition == 1'b1) ? i_input_data[911 % IN_WIDTH] : ping_storage_data_637 ^ i_input_data[911 % IN_WIDTH];
                1003 / IN_WIDTH: ping_storage_data_637 <= (fillup_transition == 1'b1) ? i_input_data[1003 % IN_WIDTH] : ping_storage_data_637 ^ i_input_data[1003 % IN_WIDTH];
                default: ping_storage_data_637 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_637;
                endcase
            end else begin
                case (input_count)
                254 / IN_WIDTH: pong_storage_data_637 <= (fillup_transition == 1'b1) ? i_input_data[254 % IN_WIDTH] : pong_storage_data_637 ^ i_input_data[254 % IN_WIDTH];
                296 / IN_WIDTH: pong_storage_data_637 <= (fillup_transition == 1'b1) ? i_input_data[296 % IN_WIDTH] : pong_storage_data_637 ^ i_input_data[296 % IN_WIDTH];
                911 / IN_WIDTH: pong_storage_data_637 <= (fillup_transition == 1'b1) ? i_input_data[911 % IN_WIDTH] : pong_storage_data_637 ^ i_input_data[911 % IN_WIDTH];
                1003 / IN_WIDTH: pong_storage_data_637 <= (fillup_transition == 1'b1) ? i_input_data[1003 % IN_WIDTH] : pong_storage_data_637 ^ i_input_data[1003 % IN_WIDTH];
                default: pong_storage_data_637 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_637;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_637 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_637;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_637 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_637;
            end
        end
    end
end

logic ping_storage_data_638;
logic pong_storage_data_638;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_638 <= 1'b0;
        pong_storage_data_638 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                255 / IN_WIDTH: ping_storage_data_638 <= (fillup_transition == 1'b1) ? i_input_data[255 % IN_WIDTH] : ping_storage_data_638 ^ i_input_data[255 % IN_WIDTH];
                297 / IN_WIDTH: ping_storage_data_638 <= (fillup_transition == 1'b1) ? i_input_data[297 % IN_WIDTH] : ping_storage_data_638 ^ i_input_data[297 % IN_WIDTH];
                912 / IN_WIDTH: ping_storage_data_638 <= (fillup_transition == 1'b1) ? i_input_data[912 % IN_WIDTH] : ping_storage_data_638 ^ i_input_data[912 % IN_WIDTH];
                1004 / IN_WIDTH: ping_storage_data_638 <= (fillup_transition == 1'b1) ? i_input_data[1004 % IN_WIDTH] : ping_storage_data_638 ^ i_input_data[1004 % IN_WIDTH];
                default: ping_storage_data_638 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_638;
                endcase
            end else begin
                case (input_count)
                255 / IN_WIDTH: pong_storage_data_638 <= (fillup_transition == 1'b1) ? i_input_data[255 % IN_WIDTH] : pong_storage_data_638 ^ i_input_data[255 % IN_WIDTH];
                297 / IN_WIDTH: pong_storage_data_638 <= (fillup_transition == 1'b1) ? i_input_data[297 % IN_WIDTH] : pong_storage_data_638 ^ i_input_data[297 % IN_WIDTH];
                912 / IN_WIDTH: pong_storage_data_638 <= (fillup_transition == 1'b1) ? i_input_data[912 % IN_WIDTH] : pong_storage_data_638 ^ i_input_data[912 % IN_WIDTH];
                1004 / IN_WIDTH: pong_storage_data_638 <= (fillup_transition == 1'b1) ? i_input_data[1004 % IN_WIDTH] : pong_storage_data_638 ^ i_input_data[1004 % IN_WIDTH];
                default: pong_storage_data_638 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_638;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_638 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_638;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_638 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_638;
            end
        end
    end
end

logic ping_storage_data_639;
logic pong_storage_data_639;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_639 <= 1'b0;
        pong_storage_data_639 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                256 / IN_WIDTH: ping_storage_data_639 <= (fillup_transition == 1'b1) ? i_input_data[256 % IN_WIDTH] : ping_storage_data_639 ^ i_input_data[256 % IN_WIDTH];
                298 / IN_WIDTH: ping_storage_data_639 <= (fillup_transition == 1'b1) ? i_input_data[298 % IN_WIDTH] : ping_storage_data_639 ^ i_input_data[298 % IN_WIDTH];
                913 / IN_WIDTH: ping_storage_data_639 <= (fillup_transition == 1'b1) ? i_input_data[913 % IN_WIDTH] : ping_storage_data_639 ^ i_input_data[913 % IN_WIDTH];
                1005 / IN_WIDTH: ping_storage_data_639 <= (fillup_transition == 1'b1) ? i_input_data[1005 % IN_WIDTH] : ping_storage_data_639 ^ i_input_data[1005 % IN_WIDTH];
                default: ping_storage_data_639 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_639;
                endcase
            end else begin
                case (input_count)
                256 / IN_WIDTH: pong_storage_data_639 <= (fillup_transition == 1'b1) ? i_input_data[256 % IN_WIDTH] : pong_storage_data_639 ^ i_input_data[256 % IN_WIDTH];
                298 / IN_WIDTH: pong_storage_data_639 <= (fillup_transition == 1'b1) ? i_input_data[298 % IN_WIDTH] : pong_storage_data_639 ^ i_input_data[298 % IN_WIDTH];
                913 / IN_WIDTH: pong_storage_data_639 <= (fillup_transition == 1'b1) ? i_input_data[913 % IN_WIDTH] : pong_storage_data_639 ^ i_input_data[913 % IN_WIDTH];
                1005 / IN_WIDTH: pong_storage_data_639 <= (fillup_transition == 1'b1) ? i_input_data[1005 % IN_WIDTH] : pong_storage_data_639 ^ i_input_data[1005 % IN_WIDTH];
                default: pong_storage_data_639 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_639;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_639 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_639;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_639 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_639;
            end
        end
    end
end

logic ping_storage_data_640;
logic pong_storage_data_640;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_640 <= 1'b0;
        pong_storage_data_640 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                257 / IN_WIDTH: ping_storage_data_640 <= (fillup_transition == 1'b1) ? i_input_data[257 % IN_WIDTH] : ping_storage_data_640 ^ i_input_data[257 % IN_WIDTH];
                299 / IN_WIDTH: ping_storage_data_640 <= (fillup_transition == 1'b1) ? i_input_data[299 % IN_WIDTH] : ping_storage_data_640 ^ i_input_data[299 % IN_WIDTH];
                914 / IN_WIDTH: ping_storage_data_640 <= (fillup_transition == 1'b1) ? i_input_data[914 % IN_WIDTH] : ping_storage_data_640 ^ i_input_data[914 % IN_WIDTH];
                1006 / IN_WIDTH: ping_storage_data_640 <= (fillup_transition == 1'b1) ? i_input_data[1006 % IN_WIDTH] : ping_storage_data_640 ^ i_input_data[1006 % IN_WIDTH];
                default: ping_storage_data_640 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_640;
                endcase
            end else begin
                case (input_count)
                257 / IN_WIDTH: pong_storage_data_640 <= (fillup_transition == 1'b1) ? i_input_data[257 % IN_WIDTH] : pong_storage_data_640 ^ i_input_data[257 % IN_WIDTH];
                299 / IN_WIDTH: pong_storage_data_640 <= (fillup_transition == 1'b1) ? i_input_data[299 % IN_WIDTH] : pong_storage_data_640 ^ i_input_data[299 % IN_WIDTH];
                914 / IN_WIDTH: pong_storage_data_640 <= (fillup_transition == 1'b1) ? i_input_data[914 % IN_WIDTH] : pong_storage_data_640 ^ i_input_data[914 % IN_WIDTH];
                1006 / IN_WIDTH: pong_storage_data_640 <= (fillup_transition == 1'b1) ? i_input_data[1006 % IN_WIDTH] : pong_storage_data_640 ^ i_input_data[1006 % IN_WIDTH];
                default: pong_storage_data_640 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_640;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_640 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_640;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_640 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_640;
            end
        end
    end
end

logic ping_storage_data_641;
logic pong_storage_data_641;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_641 <= 1'b0;
        pong_storage_data_641 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                258 / IN_WIDTH: ping_storage_data_641 <= (fillup_transition == 1'b1) ? i_input_data[258 % IN_WIDTH] : ping_storage_data_641 ^ i_input_data[258 % IN_WIDTH];
                300 / IN_WIDTH: ping_storage_data_641 <= (fillup_transition == 1'b1) ? i_input_data[300 % IN_WIDTH] : ping_storage_data_641 ^ i_input_data[300 % IN_WIDTH];
                915 / IN_WIDTH: ping_storage_data_641 <= (fillup_transition == 1'b1) ? i_input_data[915 % IN_WIDTH] : ping_storage_data_641 ^ i_input_data[915 % IN_WIDTH];
                1007 / IN_WIDTH: ping_storage_data_641 <= (fillup_transition == 1'b1) ? i_input_data[1007 % IN_WIDTH] : ping_storage_data_641 ^ i_input_data[1007 % IN_WIDTH];
                default: ping_storage_data_641 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_641;
                endcase
            end else begin
                case (input_count)
                258 / IN_WIDTH: pong_storage_data_641 <= (fillup_transition == 1'b1) ? i_input_data[258 % IN_WIDTH] : pong_storage_data_641 ^ i_input_data[258 % IN_WIDTH];
                300 / IN_WIDTH: pong_storage_data_641 <= (fillup_transition == 1'b1) ? i_input_data[300 % IN_WIDTH] : pong_storage_data_641 ^ i_input_data[300 % IN_WIDTH];
                915 / IN_WIDTH: pong_storage_data_641 <= (fillup_transition == 1'b1) ? i_input_data[915 % IN_WIDTH] : pong_storage_data_641 ^ i_input_data[915 % IN_WIDTH];
                1007 / IN_WIDTH: pong_storage_data_641 <= (fillup_transition == 1'b1) ? i_input_data[1007 % IN_WIDTH] : pong_storage_data_641 ^ i_input_data[1007 % IN_WIDTH];
                default: pong_storage_data_641 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_641;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_641 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_641;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_641 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_641;
            end
        end
    end
end

logic ping_storage_data_642;
logic pong_storage_data_642;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_642 <= 1'b0;
        pong_storage_data_642 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                259 / IN_WIDTH: ping_storage_data_642 <= (fillup_transition == 1'b1) ? i_input_data[259 % IN_WIDTH] : ping_storage_data_642 ^ i_input_data[259 % IN_WIDTH];
                301 / IN_WIDTH: ping_storage_data_642 <= (fillup_transition == 1'b1) ? i_input_data[301 % IN_WIDTH] : ping_storage_data_642 ^ i_input_data[301 % IN_WIDTH];
                916 / IN_WIDTH: ping_storage_data_642 <= (fillup_transition == 1'b1) ? i_input_data[916 % IN_WIDTH] : ping_storage_data_642 ^ i_input_data[916 % IN_WIDTH];
                1008 / IN_WIDTH: ping_storage_data_642 <= (fillup_transition == 1'b1) ? i_input_data[1008 % IN_WIDTH] : ping_storage_data_642 ^ i_input_data[1008 % IN_WIDTH];
                default: ping_storage_data_642 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_642;
                endcase
            end else begin
                case (input_count)
                259 / IN_WIDTH: pong_storage_data_642 <= (fillup_transition == 1'b1) ? i_input_data[259 % IN_WIDTH] : pong_storage_data_642 ^ i_input_data[259 % IN_WIDTH];
                301 / IN_WIDTH: pong_storage_data_642 <= (fillup_transition == 1'b1) ? i_input_data[301 % IN_WIDTH] : pong_storage_data_642 ^ i_input_data[301 % IN_WIDTH];
                916 / IN_WIDTH: pong_storage_data_642 <= (fillup_transition == 1'b1) ? i_input_data[916 % IN_WIDTH] : pong_storage_data_642 ^ i_input_data[916 % IN_WIDTH];
                1008 / IN_WIDTH: pong_storage_data_642 <= (fillup_transition == 1'b1) ? i_input_data[1008 % IN_WIDTH] : pong_storage_data_642 ^ i_input_data[1008 % IN_WIDTH];
                default: pong_storage_data_642 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_642;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_642 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_642;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_642 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_642;
            end
        end
    end
end

logic ping_storage_data_643;
logic pong_storage_data_643;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_643 <= 1'b0;
        pong_storage_data_643 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                260 / IN_WIDTH: ping_storage_data_643 <= (fillup_transition == 1'b1) ? i_input_data[260 % IN_WIDTH] : ping_storage_data_643 ^ i_input_data[260 % IN_WIDTH];
                302 / IN_WIDTH: ping_storage_data_643 <= (fillup_transition == 1'b1) ? i_input_data[302 % IN_WIDTH] : ping_storage_data_643 ^ i_input_data[302 % IN_WIDTH];
                917 / IN_WIDTH: ping_storage_data_643 <= (fillup_transition == 1'b1) ? i_input_data[917 % IN_WIDTH] : ping_storage_data_643 ^ i_input_data[917 % IN_WIDTH];
                1009 / IN_WIDTH: ping_storage_data_643 <= (fillup_transition == 1'b1) ? i_input_data[1009 % IN_WIDTH] : ping_storage_data_643 ^ i_input_data[1009 % IN_WIDTH];
                default: ping_storage_data_643 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_643;
                endcase
            end else begin
                case (input_count)
                260 / IN_WIDTH: pong_storage_data_643 <= (fillup_transition == 1'b1) ? i_input_data[260 % IN_WIDTH] : pong_storage_data_643 ^ i_input_data[260 % IN_WIDTH];
                302 / IN_WIDTH: pong_storage_data_643 <= (fillup_transition == 1'b1) ? i_input_data[302 % IN_WIDTH] : pong_storage_data_643 ^ i_input_data[302 % IN_WIDTH];
                917 / IN_WIDTH: pong_storage_data_643 <= (fillup_transition == 1'b1) ? i_input_data[917 % IN_WIDTH] : pong_storage_data_643 ^ i_input_data[917 % IN_WIDTH];
                1009 / IN_WIDTH: pong_storage_data_643 <= (fillup_transition == 1'b1) ? i_input_data[1009 % IN_WIDTH] : pong_storage_data_643 ^ i_input_data[1009 % IN_WIDTH];
                default: pong_storage_data_643 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_643;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_643 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_643;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_643 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_643;
            end
        end
    end
end

logic ping_storage_data_644;
logic pong_storage_data_644;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_644 <= 1'b0;
        pong_storage_data_644 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                261 / IN_WIDTH: ping_storage_data_644 <= (fillup_transition == 1'b1) ? i_input_data[261 % IN_WIDTH] : ping_storage_data_644 ^ i_input_data[261 % IN_WIDTH];
                303 / IN_WIDTH: ping_storage_data_644 <= (fillup_transition == 1'b1) ? i_input_data[303 % IN_WIDTH] : ping_storage_data_644 ^ i_input_data[303 % IN_WIDTH];
                918 / IN_WIDTH: ping_storage_data_644 <= (fillup_transition == 1'b1) ? i_input_data[918 % IN_WIDTH] : ping_storage_data_644 ^ i_input_data[918 % IN_WIDTH];
                1010 / IN_WIDTH: ping_storage_data_644 <= (fillup_transition == 1'b1) ? i_input_data[1010 % IN_WIDTH] : ping_storage_data_644 ^ i_input_data[1010 % IN_WIDTH];
                default: ping_storage_data_644 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_644;
                endcase
            end else begin
                case (input_count)
                261 / IN_WIDTH: pong_storage_data_644 <= (fillup_transition == 1'b1) ? i_input_data[261 % IN_WIDTH] : pong_storage_data_644 ^ i_input_data[261 % IN_WIDTH];
                303 / IN_WIDTH: pong_storage_data_644 <= (fillup_transition == 1'b1) ? i_input_data[303 % IN_WIDTH] : pong_storage_data_644 ^ i_input_data[303 % IN_WIDTH];
                918 / IN_WIDTH: pong_storage_data_644 <= (fillup_transition == 1'b1) ? i_input_data[918 % IN_WIDTH] : pong_storage_data_644 ^ i_input_data[918 % IN_WIDTH];
                1010 / IN_WIDTH: pong_storage_data_644 <= (fillup_transition == 1'b1) ? i_input_data[1010 % IN_WIDTH] : pong_storage_data_644 ^ i_input_data[1010 % IN_WIDTH];
                default: pong_storage_data_644 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_644;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_644 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_644;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_644 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_644;
            end
        end
    end
end

logic ping_storage_data_645;
logic pong_storage_data_645;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_645 <= 1'b0;
        pong_storage_data_645 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                262 / IN_WIDTH: ping_storage_data_645 <= (fillup_transition == 1'b1) ? i_input_data[262 % IN_WIDTH] : ping_storage_data_645 ^ i_input_data[262 % IN_WIDTH];
                304 / IN_WIDTH: ping_storage_data_645 <= (fillup_transition == 1'b1) ? i_input_data[304 % IN_WIDTH] : ping_storage_data_645 ^ i_input_data[304 % IN_WIDTH];
                919 / IN_WIDTH: ping_storage_data_645 <= (fillup_transition == 1'b1) ? i_input_data[919 % IN_WIDTH] : ping_storage_data_645 ^ i_input_data[919 % IN_WIDTH];
                1011 / IN_WIDTH: ping_storage_data_645 <= (fillup_transition == 1'b1) ? i_input_data[1011 % IN_WIDTH] : ping_storage_data_645 ^ i_input_data[1011 % IN_WIDTH];
                default: ping_storage_data_645 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_645;
                endcase
            end else begin
                case (input_count)
                262 / IN_WIDTH: pong_storage_data_645 <= (fillup_transition == 1'b1) ? i_input_data[262 % IN_WIDTH] : pong_storage_data_645 ^ i_input_data[262 % IN_WIDTH];
                304 / IN_WIDTH: pong_storage_data_645 <= (fillup_transition == 1'b1) ? i_input_data[304 % IN_WIDTH] : pong_storage_data_645 ^ i_input_data[304 % IN_WIDTH];
                919 / IN_WIDTH: pong_storage_data_645 <= (fillup_transition == 1'b1) ? i_input_data[919 % IN_WIDTH] : pong_storage_data_645 ^ i_input_data[919 % IN_WIDTH];
                1011 / IN_WIDTH: pong_storage_data_645 <= (fillup_transition == 1'b1) ? i_input_data[1011 % IN_WIDTH] : pong_storage_data_645 ^ i_input_data[1011 % IN_WIDTH];
                default: pong_storage_data_645 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_645;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_645 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_645;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_645 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_645;
            end
        end
    end
end

logic ping_storage_data_646;
logic pong_storage_data_646;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_646 <= 1'b0;
        pong_storage_data_646 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                263 / IN_WIDTH: ping_storage_data_646 <= (fillup_transition == 1'b1) ? i_input_data[263 % IN_WIDTH] : ping_storage_data_646 ^ i_input_data[263 % IN_WIDTH];
                305 / IN_WIDTH: ping_storage_data_646 <= (fillup_transition == 1'b1) ? i_input_data[305 % IN_WIDTH] : ping_storage_data_646 ^ i_input_data[305 % IN_WIDTH];
                920 / IN_WIDTH: ping_storage_data_646 <= (fillup_transition == 1'b1) ? i_input_data[920 % IN_WIDTH] : ping_storage_data_646 ^ i_input_data[920 % IN_WIDTH];
                1012 / IN_WIDTH: ping_storage_data_646 <= (fillup_transition == 1'b1) ? i_input_data[1012 % IN_WIDTH] : ping_storage_data_646 ^ i_input_data[1012 % IN_WIDTH];
                default: ping_storage_data_646 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_646;
                endcase
            end else begin
                case (input_count)
                263 / IN_WIDTH: pong_storage_data_646 <= (fillup_transition == 1'b1) ? i_input_data[263 % IN_WIDTH] : pong_storage_data_646 ^ i_input_data[263 % IN_WIDTH];
                305 / IN_WIDTH: pong_storage_data_646 <= (fillup_transition == 1'b1) ? i_input_data[305 % IN_WIDTH] : pong_storage_data_646 ^ i_input_data[305 % IN_WIDTH];
                920 / IN_WIDTH: pong_storage_data_646 <= (fillup_transition == 1'b1) ? i_input_data[920 % IN_WIDTH] : pong_storage_data_646 ^ i_input_data[920 % IN_WIDTH];
                1012 / IN_WIDTH: pong_storage_data_646 <= (fillup_transition == 1'b1) ? i_input_data[1012 % IN_WIDTH] : pong_storage_data_646 ^ i_input_data[1012 % IN_WIDTH];
                default: pong_storage_data_646 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_646;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_646 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_646;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_646 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_646;
            end
        end
    end
end

logic ping_storage_data_647;
logic pong_storage_data_647;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_647 <= 1'b0;
        pong_storage_data_647 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                264 / IN_WIDTH: ping_storage_data_647 <= (fillup_transition == 1'b1) ? i_input_data[264 % IN_WIDTH] : ping_storage_data_647 ^ i_input_data[264 % IN_WIDTH];
                306 / IN_WIDTH: ping_storage_data_647 <= (fillup_transition == 1'b1) ? i_input_data[306 % IN_WIDTH] : ping_storage_data_647 ^ i_input_data[306 % IN_WIDTH];
                921 / IN_WIDTH: ping_storage_data_647 <= (fillup_transition == 1'b1) ? i_input_data[921 % IN_WIDTH] : ping_storage_data_647 ^ i_input_data[921 % IN_WIDTH];
                1013 / IN_WIDTH: ping_storage_data_647 <= (fillup_transition == 1'b1) ? i_input_data[1013 % IN_WIDTH] : ping_storage_data_647 ^ i_input_data[1013 % IN_WIDTH];
                default: ping_storage_data_647 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_647;
                endcase
            end else begin
                case (input_count)
                264 / IN_WIDTH: pong_storage_data_647 <= (fillup_transition == 1'b1) ? i_input_data[264 % IN_WIDTH] : pong_storage_data_647 ^ i_input_data[264 % IN_WIDTH];
                306 / IN_WIDTH: pong_storage_data_647 <= (fillup_transition == 1'b1) ? i_input_data[306 % IN_WIDTH] : pong_storage_data_647 ^ i_input_data[306 % IN_WIDTH];
                921 / IN_WIDTH: pong_storage_data_647 <= (fillup_transition == 1'b1) ? i_input_data[921 % IN_WIDTH] : pong_storage_data_647 ^ i_input_data[921 % IN_WIDTH];
                1013 / IN_WIDTH: pong_storage_data_647 <= (fillup_transition == 1'b1) ? i_input_data[1013 % IN_WIDTH] : pong_storage_data_647 ^ i_input_data[1013 % IN_WIDTH];
                default: pong_storage_data_647 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_647;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_647 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_647;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_647 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_647;
            end
        end
    end
end

logic ping_storage_data_648;
logic pong_storage_data_648;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_648 <= 1'b0;
        pong_storage_data_648 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                265 / IN_WIDTH: ping_storage_data_648 <= (fillup_transition == 1'b1) ? i_input_data[265 % IN_WIDTH] : ping_storage_data_648 ^ i_input_data[265 % IN_WIDTH];
                307 / IN_WIDTH: ping_storage_data_648 <= (fillup_transition == 1'b1) ? i_input_data[307 % IN_WIDTH] : ping_storage_data_648 ^ i_input_data[307 % IN_WIDTH];
                922 / IN_WIDTH: ping_storage_data_648 <= (fillup_transition == 1'b1) ? i_input_data[922 % IN_WIDTH] : ping_storage_data_648 ^ i_input_data[922 % IN_WIDTH];
                1014 / IN_WIDTH: ping_storage_data_648 <= (fillup_transition == 1'b1) ? i_input_data[1014 % IN_WIDTH] : ping_storage_data_648 ^ i_input_data[1014 % IN_WIDTH];
                default: ping_storage_data_648 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_648;
                endcase
            end else begin
                case (input_count)
                265 / IN_WIDTH: pong_storage_data_648 <= (fillup_transition == 1'b1) ? i_input_data[265 % IN_WIDTH] : pong_storage_data_648 ^ i_input_data[265 % IN_WIDTH];
                307 / IN_WIDTH: pong_storage_data_648 <= (fillup_transition == 1'b1) ? i_input_data[307 % IN_WIDTH] : pong_storage_data_648 ^ i_input_data[307 % IN_WIDTH];
                922 / IN_WIDTH: pong_storage_data_648 <= (fillup_transition == 1'b1) ? i_input_data[922 % IN_WIDTH] : pong_storage_data_648 ^ i_input_data[922 % IN_WIDTH];
                1014 / IN_WIDTH: pong_storage_data_648 <= (fillup_transition == 1'b1) ? i_input_data[1014 % IN_WIDTH] : pong_storage_data_648 ^ i_input_data[1014 % IN_WIDTH];
                default: pong_storage_data_648 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_648;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_648 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_648;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_648 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_648;
            end
        end
    end
end

logic ping_storage_data_649;
logic pong_storage_data_649;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_649 <= 1'b0;
        pong_storage_data_649 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                266 / IN_WIDTH: ping_storage_data_649 <= (fillup_transition == 1'b1) ? i_input_data[266 % IN_WIDTH] : ping_storage_data_649 ^ i_input_data[266 % IN_WIDTH];
                308 / IN_WIDTH: ping_storage_data_649 <= (fillup_transition == 1'b1) ? i_input_data[308 % IN_WIDTH] : ping_storage_data_649 ^ i_input_data[308 % IN_WIDTH];
                923 / IN_WIDTH: ping_storage_data_649 <= (fillup_transition == 1'b1) ? i_input_data[923 % IN_WIDTH] : ping_storage_data_649 ^ i_input_data[923 % IN_WIDTH];
                1015 / IN_WIDTH: ping_storage_data_649 <= (fillup_transition == 1'b1) ? i_input_data[1015 % IN_WIDTH] : ping_storage_data_649 ^ i_input_data[1015 % IN_WIDTH];
                default: ping_storage_data_649 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_649;
                endcase
            end else begin
                case (input_count)
                266 / IN_WIDTH: pong_storage_data_649 <= (fillup_transition == 1'b1) ? i_input_data[266 % IN_WIDTH] : pong_storage_data_649 ^ i_input_data[266 % IN_WIDTH];
                308 / IN_WIDTH: pong_storage_data_649 <= (fillup_transition == 1'b1) ? i_input_data[308 % IN_WIDTH] : pong_storage_data_649 ^ i_input_data[308 % IN_WIDTH];
                923 / IN_WIDTH: pong_storage_data_649 <= (fillup_transition == 1'b1) ? i_input_data[923 % IN_WIDTH] : pong_storage_data_649 ^ i_input_data[923 % IN_WIDTH];
                1015 / IN_WIDTH: pong_storage_data_649 <= (fillup_transition == 1'b1) ? i_input_data[1015 % IN_WIDTH] : pong_storage_data_649 ^ i_input_data[1015 % IN_WIDTH];
                default: pong_storage_data_649 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_649;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_649 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_649;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_649 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_649;
            end
        end
    end
end

logic ping_storage_data_650;
logic pong_storage_data_650;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_650 <= 1'b0;
        pong_storage_data_650 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                267 / IN_WIDTH: ping_storage_data_650 <= (fillup_transition == 1'b1) ? i_input_data[267 % IN_WIDTH] : ping_storage_data_650 ^ i_input_data[267 % IN_WIDTH];
                309 / IN_WIDTH: ping_storage_data_650 <= (fillup_transition == 1'b1) ? i_input_data[309 % IN_WIDTH] : ping_storage_data_650 ^ i_input_data[309 % IN_WIDTH];
                924 / IN_WIDTH: ping_storage_data_650 <= (fillup_transition == 1'b1) ? i_input_data[924 % IN_WIDTH] : ping_storage_data_650 ^ i_input_data[924 % IN_WIDTH];
                1016 / IN_WIDTH: ping_storage_data_650 <= (fillup_transition == 1'b1) ? i_input_data[1016 % IN_WIDTH] : ping_storage_data_650 ^ i_input_data[1016 % IN_WIDTH];
                default: ping_storage_data_650 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_650;
                endcase
            end else begin
                case (input_count)
                267 / IN_WIDTH: pong_storage_data_650 <= (fillup_transition == 1'b1) ? i_input_data[267 % IN_WIDTH] : pong_storage_data_650 ^ i_input_data[267 % IN_WIDTH];
                309 / IN_WIDTH: pong_storage_data_650 <= (fillup_transition == 1'b1) ? i_input_data[309 % IN_WIDTH] : pong_storage_data_650 ^ i_input_data[309 % IN_WIDTH];
                924 / IN_WIDTH: pong_storage_data_650 <= (fillup_transition == 1'b1) ? i_input_data[924 % IN_WIDTH] : pong_storage_data_650 ^ i_input_data[924 % IN_WIDTH];
                1016 / IN_WIDTH: pong_storage_data_650 <= (fillup_transition == 1'b1) ? i_input_data[1016 % IN_WIDTH] : pong_storage_data_650 ^ i_input_data[1016 % IN_WIDTH];
                default: pong_storage_data_650 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_650;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_650 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_650;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_650 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_650;
            end
        end
    end
end

logic ping_storage_data_651;
logic pong_storage_data_651;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_651 <= 1'b0;
        pong_storage_data_651 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                268 / IN_WIDTH: ping_storage_data_651 <= (fillup_transition == 1'b1) ? i_input_data[268 % IN_WIDTH] : ping_storage_data_651 ^ i_input_data[268 % IN_WIDTH];
                310 / IN_WIDTH: ping_storage_data_651 <= (fillup_transition == 1'b1) ? i_input_data[310 % IN_WIDTH] : ping_storage_data_651 ^ i_input_data[310 % IN_WIDTH];
                925 / IN_WIDTH: ping_storage_data_651 <= (fillup_transition == 1'b1) ? i_input_data[925 % IN_WIDTH] : ping_storage_data_651 ^ i_input_data[925 % IN_WIDTH];
                1017 / IN_WIDTH: ping_storage_data_651 <= (fillup_transition == 1'b1) ? i_input_data[1017 % IN_WIDTH] : ping_storage_data_651 ^ i_input_data[1017 % IN_WIDTH];
                default: ping_storage_data_651 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_651;
                endcase
            end else begin
                case (input_count)
                268 / IN_WIDTH: pong_storage_data_651 <= (fillup_transition == 1'b1) ? i_input_data[268 % IN_WIDTH] : pong_storage_data_651 ^ i_input_data[268 % IN_WIDTH];
                310 / IN_WIDTH: pong_storage_data_651 <= (fillup_transition == 1'b1) ? i_input_data[310 % IN_WIDTH] : pong_storage_data_651 ^ i_input_data[310 % IN_WIDTH];
                925 / IN_WIDTH: pong_storage_data_651 <= (fillup_transition == 1'b1) ? i_input_data[925 % IN_WIDTH] : pong_storage_data_651 ^ i_input_data[925 % IN_WIDTH];
                1017 / IN_WIDTH: pong_storage_data_651 <= (fillup_transition == 1'b1) ? i_input_data[1017 % IN_WIDTH] : pong_storage_data_651 ^ i_input_data[1017 % IN_WIDTH];
                default: pong_storage_data_651 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_651;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_651 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_651;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_651 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_651;
            end
        end
    end
end

logic ping_storage_data_652;
logic pong_storage_data_652;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_652 <= 1'b0;
        pong_storage_data_652 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                269 / IN_WIDTH: ping_storage_data_652 <= (fillup_transition == 1'b1) ? i_input_data[269 % IN_WIDTH] : ping_storage_data_652 ^ i_input_data[269 % IN_WIDTH];
                311 / IN_WIDTH: ping_storage_data_652 <= (fillup_transition == 1'b1) ? i_input_data[311 % IN_WIDTH] : ping_storage_data_652 ^ i_input_data[311 % IN_WIDTH];
                926 / IN_WIDTH: ping_storage_data_652 <= (fillup_transition == 1'b1) ? i_input_data[926 % IN_WIDTH] : ping_storage_data_652 ^ i_input_data[926 % IN_WIDTH];
                1018 / IN_WIDTH: ping_storage_data_652 <= (fillup_transition == 1'b1) ? i_input_data[1018 % IN_WIDTH] : ping_storage_data_652 ^ i_input_data[1018 % IN_WIDTH];
                default: ping_storage_data_652 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_652;
                endcase
            end else begin
                case (input_count)
                269 / IN_WIDTH: pong_storage_data_652 <= (fillup_transition == 1'b1) ? i_input_data[269 % IN_WIDTH] : pong_storage_data_652 ^ i_input_data[269 % IN_WIDTH];
                311 / IN_WIDTH: pong_storage_data_652 <= (fillup_transition == 1'b1) ? i_input_data[311 % IN_WIDTH] : pong_storage_data_652 ^ i_input_data[311 % IN_WIDTH];
                926 / IN_WIDTH: pong_storage_data_652 <= (fillup_transition == 1'b1) ? i_input_data[926 % IN_WIDTH] : pong_storage_data_652 ^ i_input_data[926 % IN_WIDTH];
                1018 / IN_WIDTH: pong_storage_data_652 <= (fillup_transition == 1'b1) ? i_input_data[1018 % IN_WIDTH] : pong_storage_data_652 ^ i_input_data[1018 % IN_WIDTH];
                default: pong_storage_data_652 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_652;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_652 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_652;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_652 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_652;
            end
        end
    end
end

logic ping_storage_data_653;
logic pong_storage_data_653;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_653 <= 1'b0;
        pong_storage_data_653 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                270 / IN_WIDTH: ping_storage_data_653 <= (fillup_transition == 1'b1) ? i_input_data[270 % IN_WIDTH] : ping_storage_data_653 ^ i_input_data[270 % IN_WIDTH];
                312 / IN_WIDTH: ping_storage_data_653 <= (fillup_transition == 1'b1) ? i_input_data[312 % IN_WIDTH] : ping_storage_data_653 ^ i_input_data[312 % IN_WIDTH];
                927 / IN_WIDTH: ping_storage_data_653 <= (fillup_transition == 1'b1) ? i_input_data[927 % IN_WIDTH] : ping_storage_data_653 ^ i_input_data[927 % IN_WIDTH];
                1019 / IN_WIDTH: ping_storage_data_653 <= (fillup_transition == 1'b1) ? i_input_data[1019 % IN_WIDTH] : ping_storage_data_653 ^ i_input_data[1019 % IN_WIDTH];
                default: ping_storage_data_653 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_653;
                endcase
            end else begin
                case (input_count)
                270 / IN_WIDTH: pong_storage_data_653 <= (fillup_transition == 1'b1) ? i_input_data[270 % IN_WIDTH] : pong_storage_data_653 ^ i_input_data[270 % IN_WIDTH];
                312 / IN_WIDTH: pong_storage_data_653 <= (fillup_transition == 1'b1) ? i_input_data[312 % IN_WIDTH] : pong_storage_data_653 ^ i_input_data[312 % IN_WIDTH];
                927 / IN_WIDTH: pong_storage_data_653 <= (fillup_transition == 1'b1) ? i_input_data[927 % IN_WIDTH] : pong_storage_data_653 ^ i_input_data[927 % IN_WIDTH];
                1019 / IN_WIDTH: pong_storage_data_653 <= (fillup_transition == 1'b1) ? i_input_data[1019 % IN_WIDTH] : pong_storage_data_653 ^ i_input_data[1019 % IN_WIDTH];
                default: pong_storage_data_653 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_653;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_653 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_653;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_653 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_653;
            end
        end
    end
end

logic ping_storage_data_654;
logic pong_storage_data_654;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_654 <= 1'b0;
        pong_storage_data_654 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                271 / IN_WIDTH: ping_storage_data_654 <= (fillup_transition == 1'b1) ? i_input_data[271 % IN_WIDTH] : ping_storage_data_654 ^ i_input_data[271 % IN_WIDTH];
                313 / IN_WIDTH: ping_storage_data_654 <= (fillup_transition == 1'b1) ? i_input_data[313 % IN_WIDTH] : ping_storage_data_654 ^ i_input_data[313 % IN_WIDTH];
                928 / IN_WIDTH: ping_storage_data_654 <= (fillup_transition == 1'b1) ? i_input_data[928 % IN_WIDTH] : ping_storage_data_654 ^ i_input_data[928 % IN_WIDTH];
                1020 / IN_WIDTH: ping_storage_data_654 <= (fillup_transition == 1'b1) ? i_input_data[1020 % IN_WIDTH] : ping_storage_data_654 ^ i_input_data[1020 % IN_WIDTH];
                default: ping_storage_data_654 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_654;
                endcase
            end else begin
                case (input_count)
                271 / IN_WIDTH: pong_storage_data_654 <= (fillup_transition == 1'b1) ? i_input_data[271 % IN_WIDTH] : pong_storage_data_654 ^ i_input_data[271 % IN_WIDTH];
                313 / IN_WIDTH: pong_storage_data_654 <= (fillup_transition == 1'b1) ? i_input_data[313 % IN_WIDTH] : pong_storage_data_654 ^ i_input_data[313 % IN_WIDTH];
                928 / IN_WIDTH: pong_storage_data_654 <= (fillup_transition == 1'b1) ? i_input_data[928 % IN_WIDTH] : pong_storage_data_654 ^ i_input_data[928 % IN_WIDTH];
                1020 / IN_WIDTH: pong_storage_data_654 <= (fillup_transition == 1'b1) ? i_input_data[1020 % IN_WIDTH] : pong_storage_data_654 ^ i_input_data[1020 % IN_WIDTH];
                default: pong_storage_data_654 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_654;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_654 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_654;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_654 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_654;
            end
        end
    end
end

logic ping_storage_data_655;
logic pong_storage_data_655;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_655 <= 1'b0;
        pong_storage_data_655 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                272 / IN_WIDTH: ping_storage_data_655 <= (fillup_transition == 1'b1) ? i_input_data[272 % IN_WIDTH] : ping_storage_data_655 ^ i_input_data[272 % IN_WIDTH];
                314 / IN_WIDTH: ping_storage_data_655 <= (fillup_transition == 1'b1) ? i_input_data[314 % IN_WIDTH] : ping_storage_data_655 ^ i_input_data[314 % IN_WIDTH];
                929 / IN_WIDTH: ping_storage_data_655 <= (fillup_transition == 1'b1) ? i_input_data[929 % IN_WIDTH] : ping_storage_data_655 ^ i_input_data[929 % IN_WIDTH];
                1021 / IN_WIDTH: ping_storage_data_655 <= (fillup_transition == 1'b1) ? i_input_data[1021 % IN_WIDTH] : ping_storage_data_655 ^ i_input_data[1021 % IN_WIDTH];
                default: ping_storage_data_655 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_655;
                endcase
            end else begin
                case (input_count)
                272 / IN_WIDTH: pong_storage_data_655 <= (fillup_transition == 1'b1) ? i_input_data[272 % IN_WIDTH] : pong_storage_data_655 ^ i_input_data[272 % IN_WIDTH];
                314 / IN_WIDTH: pong_storage_data_655 <= (fillup_transition == 1'b1) ? i_input_data[314 % IN_WIDTH] : pong_storage_data_655 ^ i_input_data[314 % IN_WIDTH];
                929 / IN_WIDTH: pong_storage_data_655 <= (fillup_transition == 1'b1) ? i_input_data[929 % IN_WIDTH] : pong_storage_data_655 ^ i_input_data[929 % IN_WIDTH];
                1021 / IN_WIDTH: pong_storage_data_655 <= (fillup_transition == 1'b1) ? i_input_data[1021 % IN_WIDTH] : pong_storage_data_655 ^ i_input_data[1021 % IN_WIDTH];
                default: pong_storage_data_655 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_655;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_655 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_655;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_655 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_655;
            end
        end
    end
end

logic ping_storage_data_656;
logic pong_storage_data_656;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_656 <= 1'b0;
        pong_storage_data_656 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                273 / IN_WIDTH: ping_storage_data_656 <= (fillup_transition == 1'b1) ? i_input_data[273 % IN_WIDTH] : ping_storage_data_656 ^ i_input_data[273 % IN_WIDTH];
                315 / IN_WIDTH: ping_storage_data_656 <= (fillup_transition == 1'b1) ? i_input_data[315 % IN_WIDTH] : ping_storage_data_656 ^ i_input_data[315 % IN_WIDTH];
                930 / IN_WIDTH: ping_storage_data_656 <= (fillup_transition == 1'b1) ? i_input_data[930 % IN_WIDTH] : ping_storage_data_656 ^ i_input_data[930 % IN_WIDTH];
                1022 / IN_WIDTH: ping_storage_data_656 <= (fillup_transition == 1'b1) ? i_input_data[1022 % IN_WIDTH] : ping_storage_data_656 ^ i_input_data[1022 % IN_WIDTH];
                default: ping_storage_data_656 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_656;
                endcase
            end else begin
                case (input_count)
                273 / IN_WIDTH: pong_storage_data_656 <= (fillup_transition == 1'b1) ? i_input_data[273 % IN_WIDTH] : pong_storage_data_656 ^ i_input_data[273 % IN_WIDTH];
                315 / IN_WIDTH: pong_storage_data_656 <= (fillup_transition == 1'b1) ? i_input_data[315 % IN_WIDTH] : pong_storage_data_656 ^ i_input_data[315 % IN_WIDTH];
                930 / IN_WIDTH: pong_storage_data_656 <= (fillup_transition == 1'b1) ? i_input_data[930 % IN_WIDTH] : pong_storage_data_656 ^ i_input_data[930 % IN_WIDTH];
                1022 / IN_WIDTH: pong_storage_data_656 <= (fillup_transition == 1'b1) ? i_input_data[1022 % IN_WIDTH] : pong_storage_data_656 ^ i_input_data[1022 % IN_WIDTH];
                default: pong_storage_data_656 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_656;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_656 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_656;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_656 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_656;
            end
        end
    end
end

logic ping_storage_data_657;
logic pong_storage_data_657;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_657 <= 1'b0;
        pong_storage_data_657 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                274 / IN_WIDTH: ping_storage_data_657 <= (fillup_transition == 1'b1) ? i_input_data[274 % IN_WIDTH] : ping_storage_data_657 ^ i_input_data[274 % IN_WIDTH];
                316 / IN_WIDTH: ping_storage_data_657 <= (fillup_transition == 1'b1) ? i_input_data[316 % IN_WIDTH] : ping_storage_data_657 ^ i_input_data[316 % IN_WIDTH];
                931 / IN_WIDTH: ping_storage_data_657 <= (fillup_transition == 1'b1) ? i_input_data[931 % IN_WIDTH] : ping_storage_data_657 ^ i_input_data[931 % IN_WIDTH];
                1023 / IN_WIDTH: ping_storage_data_657 <= (fillup_transition == 1'b1) ? i_input_data[1023 % IN_WIDTH] : ping_storage_data_657 ^ i_input_data[1023 % IN_WIDTH];
                default: ping_storage_data_657 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_657;
                endcase
            end else begin
                case (input_count)
                274 / IN_WIDTH: pong_storage_data_657 <= (fillup_transition == 1'b1) ? i_input_data[274 % IN_WIDTH] : pong_storage_data_657 ^ i_input_data[274 % IN_WIDTH];
                316 / IN_WIDTH: pong_storage_data_657 <= (fillup_transition == 1'b1) ? i_input_data[316 % IN_WIDTH] : pong_storage_data_657 ^ i_input_data[316 % IN_WIDTH];
                931 / IN_WIDTH: pong_storage_data_657 <= (fillup_transition == 1'b1) ? i_input_data[931 % IN_WIDTH] : pong_storage_data_657 ^ i_input_data[931 % IN_WIDTH];
                1023 / IN_WIDTH: pong_storage_data_657 <= (fillup_transition == 1'b1) ? i_input_data[1023 % IN_WIDTH] : pong_storage_data_657 ^ i_input_data[1023 % IN_WIDTH];
                default: pong_storage_data_657 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_657;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_657 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_657;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_657 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_657;
            end
        end
    end
end

logic ping_storage_data_658;
logic pong_storage_data_658;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_658 <= 1'b0;
        pong_storage_data_658 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                275 / IN_WIDTH: ping_storage_data_658 <= (fillup_transition == 1'b1) ? i_input_data[275 % IN_WIDTH] : ping_storage_data_658 ^ i_input_data[275 % IN_WIDTH];
                317 / IN_WIDTH: ping_storage_data_658 <= (fillup_transition == 1'b1) ? i_input_data[317 % IN_WIDTH] : ping_storage_data_658 ^ i_input_data[317 % IN_WIDTH];
                932 / IN_WIDTH: ping_storage_data_658 <= (fillup_transition == 1'b1) ? i_input_data[932 % IN_WIDTH] : ping_storage_data_658 ^ i_input_data[932 % IN_WIDTH];
                1024 / IN_WIDTH: ping_storage_data_658 <= (fillup_transition == 1'b1) ? i_input_data[1024 % IN_WIDTH] : ping_storage_data_658 ^ i_input_data[1024 % IN_WIDTH];
                default: ping_storage_data_658 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_658;
                endcase
            end else begin
                case (input_count)
                275 / IN_WIDTH: pong_storage_data_658 <= (fillup_transition == 1'b1) ? i_input_data[275 % IN_WIDTH] : pong_storage_data_658 ^ i_input_data[275 % IN_WIDTH];
                317 / IN_WIDTH: pong_storage_data_658 <= (fillup_transition == 1'b1) ? i_input_data[317 % IN_WIDTH] : pong_storage_data_658 ^ i_input_data[317 % IN_WIDTH];
                932 / IN_WIDTH: pong_storage_data_658 <= (fillup_transition == 1'b1) ? i_input_data[932 % IN_WIDTH] : pong_storage_data_658 ^ i_input_data[932 % IN_WIDTH];
                1024 / IN_WIDTH: pong_storage_data_658 <= (fillup_transition == 1'b1) ? i_input_data[1024 % IN_WIDTH] : pong_storage_data_658 ^ i_input_data[1024 % IN_WIDTH];
                default: pong_storage_data_658 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_658;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_658 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_658;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_658 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_658;
            end
        end
    end
end

logic ping_storage_data_659;
logic pong_storage_data_659;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_659 <= 1'b0;
        pong_storage_data_659 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                276 / IN_WIDTH: ping_storage_data_659 <= (fillup_transition == 1'b1) ? i_input_data[276 % IN_WIDTH] : ping_storage_data_659 ^ i_input_data[276 % IN_WIDTH];
                318 / IN_WIDTH: ping_storage_data_659 <= (fillup_transition == 1'b1) ? i_input_data[318 % IN_WIDTH] : ping_storage_data_659 ^ i_input_data[318 % IN_WIDTH];
                933 / IN_WIDTH: ping_storage_data_659 <= (fillup_transition == 1'b1) ? i_input_data[933 % IN_WIDTH] : ping_storage_data_659 ^ i_input_data[933 % IN_WIDTH];
                1025 / IN_WIDTH: ping_storage_data_659 <= (fillup_transition == 1'b1) ? i_input_data[1025 % IN_WIDTH] : ping_storage_data_659 ^ i_input_data[1025 % IN_WIDTH];
                default: ping_storage_data_659 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_659;
                endcase
            end else begin
                case (input_count)
                276 / IN_WIDTH: pong_storage_data_659 <= (fillup_transition == 1'b1) ? i_input_data[276 % IN_WIDTH] : pong_storage_data_659 ^ i_input_data[276 % IN_WIDTH];
                318 / IN_WIDTH: pong_storage_data_659 <= (fillup_transition == 1'b1) ? i_input_data[318 % IN_WIDTH] : pong_storage_data_659 ^ i_input_data[318 % IN_WIDTH];
                933 / IN_WIDTH: pong_storage_data_659 <= (fillup_transition == 1'b1) ? i_input_data[933 % IN_WIDTH] : pong_storage_data_659 ^ i_input_data[933 % IN_WIDTH];
                1025 / IN_WIDTH: pong_storage_data_659 <= (fillup_transition == 1'b1) ? i_input_data[1025 % IN_WIDTH] : pong_storage_data_659 ^ i_input_data[1025 % IN_WIDTH];
                default: pong_storage_data_659 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_659;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_659 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_659;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_659 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_659;
            end
        end
    end
end

logic ping_storage_data_660;
logic pong_storage_data_660;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_660 <= 1'b0;
        pong_storage_data_660 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                277 / IN_WIDTH: ping_storage_data_660 <= (fillup_transition == 1'b1) ? i_input_data[277 % IN_WIDTH] : ping_storage_data_660 ^ i_input_data[277 % IN_WIDTH];
                319 / IN_WIDTH: ping_storage_data_660 <= (fillup_transition == 1'b1) ? i_input_data[319 % IN_WIDTH] : ping_storage_data_660 ^ i_input_data[319 % IN_WIDTH];
                934 / IN_WIDTH: ping_storage_data_660 <= (fillup_transition == 1'b1) ? i_input_data[934 % IN_WIDTH] : ping_storage_data_660 ^ i_input_data[934 % IN_WIDTH];
                1026 / IN_WIDTH: ping_storage_data_660 <= (fillup_transition == 1'b1) ? i_input_data[1026 % IN_WIDTH] : ping_storage_data_660 ^ i_input_data[1026 % IN_WIDTH];
                default: ping_storage_data_660 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_660;
                endcase
            end else begin
                case (input_count)
                277 / IN_WIDTH: pong_storage_data_660 <= (fillup_transition == 1'b1) ? i_input_data[277 % IN_WIDTH] : pong_storage_data_660 ^ i_input_data[277 % IN_WIDTH];
                319 / IN_WIDTH: pong_storage_data_660 <= (fillup_transition == 1'b1) ? i_input_data[319 % IN_WIDTH] : pong_storage_data_660 ^ i_input_data[319 % IN_WIDTH];
                934 / IN_WIDTH: pong_storage_data_660 <= (fillup_transition == 1'b1) ? i_input_data[934 % IN_WIDTH] : pong_storage_data_660 ^ i_input_data[934 % IN_WIDTH];
                1026 / IN_WIDTH: pong_storage_data_660 <= (fillup_transition == 1'b1) ? i_input_data[1026 % IN_WIDTH] : pong_storage_data_660 ^ i_input_data[1026 % IN_WIDTH];
                default: pong_storage_data_660 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_660;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_660 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_660;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_660 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_660;
            end
        end
    end
end

logic ping_storage_data_661;
logic pong_storage_data_661;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_661 <= 1'b0;
        pong_storage_data_661 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                278 / IN_WIDTH: ping_storage_data_661 <= (fillup_transition == 1'b1) ? i_input_data[278 % IN_WIDTH] : ping_storage_data_661 ^ i_input_data[278 % IN_WIDTH];
                320 / IN_WIDTH: ping_storage_data_661 <= (fillup_transition == 1'b1) ? i_input_data[320 % IN_WIDTH] : ping_storage_data_661 ^ i_input_data[320 % IN_WIDTH];
                935 / IN_WIDTH: ping_storage_data_661 <= (fillup_transition == 1'b1) ? i_input_data[935 % IN_WIDTH] : ping_storage_data_661 ^ i_input_data[935 % IN_WIDTH];
                1027 / IN_WIDTH: ping_storage_data_661 <= (fillup_transition == 1'b1) ? i_input_data[1027 % IN_WIDTH] : ping_storage_data_661 ^ i_input_data[1027 % IN_WIDTH];
                default: ping_storage_data_661 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_661;
                endcase
            end else begin
                case (input_count)
                278 / IN_WIDTH: pong_storage_data_661 <= (fillup_transition == 1'b1) ? i_input_data[278 % IN_WIDTH] : pong_storage_data_661 ^ i_input_data[278 % IN_WIDTH];
                320 / IN_WIDTH: pong_storage_data_661 <= (fillup_transition == 1'b1) ? i_input_data[320 % IN_WIDTH] : pong_storage_data_661 ^ i_input_data[320 % IN_WIDTH];
                935 / IN_WIDTH: pong_storage_data_661 <= (fillup_transition == 1'b1) ? i_input_data[935 % IN_WIDTH] : pong_storage_data_661 ^ i_input_data[935 % IN_WIDTH];
                1027 / IN_WIDTH: pong_storage_data_661 <= (fillup_transition == 1'b1) ? i_input_data[1027 % IN_WIDTH] : pong_storage_data_661 ^ i_input_data[1027 % IN_WIDTH];
                default: pong_storage_data_661 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_661;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_661 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_661;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_661 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_661;
            end
        end
    end
end

logic ping_storage_data_662;
logic pong_storage_data_662;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_662 <= 1'b0;
        pong_storage_data_662 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                279 / IN_WIDTH: ping_storage_data_662 <= (fillup_transition == 1'b1) ? i_input_data[279 % IN_WIDTH] : ping_storage_data_662 ^ i_input_data[279 % IN_WIDTH];
                321 / IN_WIDTH: ping_storage_data_662 <= (fillup_transition == 1'b1) ? i_input_data[321 % IN_WIDTH] : ping_storage_data_662 ^ i_input_data[321 % IN_WIDTH];
                936 / IN_WIDTH: ping_storage_data_662 <= (fillup_transition == 1'b1) ? i_input_data[936 % IN_WIDTH] : ping_storage_data_662 ^ i_input_data[936 % IN_WIDTH];
                1028 / IN_WIDTH: ping_storage_data_662 <= (fillup_transition == 1'b1) ? i_input_data[1028 % IN_WIDTH] : ping_storage_data_662 ^ i_input_data[1028 % IN_WIDTH];
                default: ping_storage_data_662 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_662;
                endcase
            end else begin
                case (input_count)
                279 / IN_WIDTH: pong_storage_data_662 <= (fillup_transition == 1'b1) ? i_input_data[279 % IN_WIDTH] : pong_storage_data_662 ^ i_input_data[279 % IN_WIDTH];
                321 / IN_WIDTH: pong_storage_data_662 <= (fillup_transition == 1'b1) ? i_input_data[321 % IN_WIDTH] : pong_storage_data_662 ^ i_input_data[321 % IN_WIDTH];
                936 / IN_WIDTH: pong_storage_data_662 <= (fillup_transition == 1'b1) ? i_input_data[936 % IN_WIDTH] : pong_storage_data_662 ^ i_input_data[936 % IN_WIDTH];
                1028 / IN_WIDTH: pong_storage_data_662 <= (fillup_transition == 1'b1) ? i_input_data[1028 % IN_WIDTH] : pong_storage_data_662 ^ i_input_data[1028 % IN_WIDTH];
                default: pong_storage_data_662 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_662;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_662 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_662;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_662 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_662;
            end
        end
    end
end

logic ping_storage_data_663;
logic pong_storage_data_663;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_663 <= 1'b0;
        pong_storage_data_663 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                280 / IN_WIDTH: ping_storage_data_663 <= (fillup_transition == 1'b1) ? i_input_data[280 % IN_WIDTH] : ping_storage_data_663 ^ i_input_data[280 % IN_WIDTH];
                322 / IN_WIDTH: ping_storage_data_663 <= (fillup_transition == 1'b1) ? i_input_data[322 % IN_WIDTH] : ping_storage_data_663 ^ i_input_data[322 % IN_WIDTH];
                937 / IN_WIDTH: ping_storage_data_663 <= (fillup_transition == 1'b1) ? i_input_data[937 % IN_WIDTH] : ping_storage_data_663 ^ i_input_data[937 % IN_WIDTH];
                1029 / IN_WIDTH: ping_storage_data_663 <= (fillup_transition == 1'b1) ? i_input_data[1029 % IN_WIDTH] : ping_storage_data_663 ^ i_input_data[1029 % IN_WIDTH];
                default: ping_storage_data_663 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_663;
                endcase
            end else begin
                case (input_count)
                280 / IN_WIDTH: pong_storage_data_663 <= (fillup_transition == 1'b1) ? i_input_data[280 % IN_WIDTH] : pong_storage_data_663 ^ i_input_data[280 % IN_WIDTH];
                322 / IN_WIDTH: pong_storage_data_663 <= (fillup_transition == 1'b1) ? i_input_data[322 % IN_WIDTH] : pong_storage_data_663 ^ i_input_data[322 % IN_WIDTH];
                937 / IN_WIDTH: pong_storage_data_663 <= (fillup_transition == 1'b1) ? i_input_data[937 % IN_WIDTH] : pong_storage_data_663 ^ i_input_data[937 % IN_WIDTH];
                1029 / IN_WIDTH: pong_storage_data_663 <= (fillup_transition == 1'b1) ? i_input_data[1029 % IN_WIDTH] : pong_storage_data_663 ^ i_input_data[1029 % IN_WIDTH];
                default: pong_storage_data_663 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_663;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_663 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_663;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_663 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_663;
            end
        end
    end
end

logic ping_storage_data_664;
logic pong_storage_data_664;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_664 <= 1'b0;
        pong_storage_data_664 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                281 / IN_WIDTH: ping_storage_data_664 <= (fillup_transition == 1'b1) ? i_input_data[281 % IN_WIDTH] : ping_storage_data_664 ^ i_input_data[281 % IN_WIDTH];
                323 / IN_WIDTH: ping_storage_data_664 <= (fillup_transition == 1'b1) ? i_input_data[323 % IN_WIDTH] : ping_storage_data_664 ^ i_input_data[323 % IN_WIDTH];
                938 / IN_WIDTH: ping_storage_data_664 <= (fillup_transition == 1'b1) ? i_input_data[938 % IN_WIDTH] : ping_storage_data_664 ^ i_input_data[938 % IN_WIDTH];
                1030 / IN_WIDTH: ping_storage_data_664 <= (fillup_transition == 1'b1) ? i_input_data[1030 % IN_WIDTH] : ping_storage_data_664 ^ i_input_data[1030 % IN_WIDTH];
                default: ping_storage_data_664 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_664;
                endcase
            end else begin
                case (input_count)
                281 / IN_WIDTH: pong_storage_data_664 <= (fillup_transition == 1'b1) ? i_input_data[281 % IN_WIDTH] : pong_storage_data_664 ^ i_input_data[281 % IN_WIDTH];
                323 / IN_WIDTH: pong_storage_data_664 <= (fillup_transition == 1'b1) ? i_input_data[323 % IN_WIDTH] : pong_storage_data_664 ^ i_input_data[323 % IN_WIDTH];
                938 / IN_WIDTH: pong_storage_data_664 <= (fillup_transition == 1'b1) ? i_input_data[938 % IN_WIDTH] : pong_storage_data_664 ^ i_input_data[938 % IN_WIDTH];
                1030 / IN_WIDTH: pong_storage_data_664 <= (fillup_transition == 1'b1) ? i_input_data[1030 % IN_WIDTH] : pong_storage_data_664 ^ i_input_data[1030 % IN_WIDTH];
                default: pong_storage_data_664 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_664;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_664 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_664;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_664 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_664;
            end
        end
    end
end

logic ping_storage_data_665;
logic pong_storage_data_665;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_665 <= 1'b0;
        pong_storage_data_665 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                282 / IN_WIDTH: ping_storage_data_665 <= (fillup_transition == 1'b1) ? i_input_data[282 % IN_WIDTH] : ping_storage_data_665 ^ i_input_data[282 % IN_WIDTH];
                324 / IN_WIDTH: ping_storage_data_665 <= (fillup_transition == 1'b1) ? i_input_data[324 % IN_WIDTH] : ping_storage_data_665 ^ i_input_data[324 % IN_WIDTH];
                939 / IN_WIDTH: ping_storage_data_665 <= (fillup_transition == 1'b1) ? i_input_data[939 % IN_WIDTH] : ping_storage_data_665 ^ i_input_data[939 % IN_WIDTH];
                1031 / IN_WIDTH: ping_storage_data_665 <= (fillup_transition == 1'b1) ? i_input_data[1031 % IN_WIDTH] : ping_storage_data_665 ^ i_input_data[1031 % IN_WIDTH];
                default: ping_storage_data_665 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_665;
                endcase
            end else begin
                case (input_count)
                282 / IN_WIDTH: pong_storage_data_665 <= (fillup_transition == 1'b1) ? i_input_data[282 % IN_WIDTH] : pong_storage_data_665 ^ i_input_data[282 % IN_WIDTH];
                324 / IN_WIDTH: pong_storage_data_665 <= (fillup_transition == 1'b1) ? i_input_data[324 % IN_WIDTH] : pong_storage_data_665 ^ i_input_data[324 % IN_WIDTH];
                939 / IN_WIDTH: pong_storage_data_665 <= (fillup_transition == 1'b1) ? i_input_data[939 % IN_WIDTH] : pong_storage_data_665 ^ i_input_data[939 % IN_WIDTH];
                1031 / IN_WIDTH: pong_storage_data_665 <= (fillup_transition == 1'b1) ? i_input_data[1031 % IN_WIDTH] : pong_storage_data_665 ^ i_input_data[1031 % IN_WIDTH];
                default: pong_storage_data_665 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_665;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_665 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_665;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_665 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_665;
            end
        end
    end
end

logic ping_storage_data_666;
logic pong_storage_data_666;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_666 <= 1'b0;
        pong_storage_data_666 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                283 / IN_WIDTH: ping_storage_data_666 <= (fillup_transition == 1'b1) ? i_input_data[283 % IN_WIDTH] : ping_storage_data_666 ^ i_input_data[283 % IN_WIDTH];
                325 / IN_WIDTH: ping_storage_data_666 <= (fillup_transition == 1'b1) ? i_input_data[325 % IN_WIDTH] : ping_storage_data_666 ^ i_input_data[325 % IN_WIDTH];
                940 / IN_WIDTH: ping_storage_data_666 <= (fillup_transition == 1'b1) ? i_input_data[940 % IN_WIDTH] : ping_storage_data_666 ^ i_input_data[940 % IN_WIDTH];
                1032 / IN_WIDTH: ping_storage_data_666 <= (fillup_transition == 1'b1) ? i_input_data[1032 % IN_WIDTH] : ping_storage_data_666 ^ i_input_data[1032 % IN_WIDTH];
                default: ping_storage_data_666 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_666;
                endcase
            end else begin
                case (input_count)
                283 / IN_WIDTH: pong_storage_data_666 <= (fillup_transition == 1'b1) ? i_input_data[283 % IN_WIDTH] : pong_storage_data_666 ^ i_input_data[283 % IN_WIDTH];
                325 / IN_WIDTH: pong_storage_data_666 <= (fillup_transition == 1'b1) ? i_input_data[325 % IN_WIDTH] : pong_storage_data_666 ^ i_input_data[325 % IN_WIDTH];
                940 / IN_WIDTH: pong_storage_data_666 <= (fillup_transition == 1'b1) ? i_input_data[940 % IN_WIDTH] : pong_storage_data_666 ^ i_input_data[940 % IN_WIDTH];
                1032 / IN_WIDTH: pong_storage_data_666 <= (fillup_transition == 1'b1) ? i_input_data[1032 % IN_WIDTH] : pong_storage_data_666 ^ i_input_data[1032 % IN_WIDTH];
                default: pong_storage_data_666 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_666;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_666 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_666;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_666 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_666;
            end
        end
    end
end

logic ping_storage_data_667;
logic pong_storage_data_667;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_667 <= 1'b0;
        pong_storage_data_667 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                284 / IN_WIDTH: ping_storage_data_667 <= (fillup_transition == 1'b1) ? i_input_data[284 % IN_WIDTH] : ping_storage_data_667 ^ i_input_data[284 % IN_WIDTH];
                326 / IN_WIDTH: ping_storage_data_667 <= (fillup_transition == 1'b1) ? i_input_data[326 % IN_WIDTH] : ping_storage_data_667 ^ i_input_data[326 % IN_WIDTH];
                941 / IN_WIDTH: ping_storage_data_667 <= (fillup_transition == 1'b1) ? i_input_data[941 % IN_WIDTH] : ping_storage_data_667 ^ i_input_data[941 % IN_WIDTH];
                1033 / IN_WIDTH: ping_storage_data_667 <= (fillup_transition == 1'b1) ? i_input_data[1033 % IN_WIDTH] : ping_storage_data_667 ^ i_input_data[1033 % IN_WIDTH];
                default: ping_storage_data_667 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_667;
                endcase
            end else begin
                case (input_count)
                284 / IN_WIDTH: pong_storage_data_667 <= (fillup_transition == 1'b1) ? i_input_data[284 % IN_WIDTH] : pong_storage_data_667 ^ i_input_data[284 % IN_WIDTH];
                326 / IN_WIDTH: pong_storage_data_667 <= (fillup_transition == 1'b1) ? i_input_data[326 % IN_WIDTH] : pong_storage_data_667 ^ i_input_data[326 % IN_WIDTH];
                941 / IN_WIDTH: pong_storage_data_667 <= (fillup_transition == 1'b1) ? i_input_data[941 % IN_WIDTH] : pong_storage_data_667 ^ i_input_data[941 % IN_WIDTH];
                1033 / IN_WIDTH: pong_storage_data_667 <= (fillup_transition == 1'b1) ? i_input_data[1033 % IN_WIDTH] : pong_storage_data_667 ^ i_input_data[1033 % IN_WIDTH];
                default: pong_storage_data_667 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_667;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_667 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_667;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_667 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_667;
            end
        end
    end
end

logic ping_storage_data_668;
logic pong_storage_data_668;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_668 <= 1'b0;
        pong_storage_data_668 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                285 / IN_WIDTH: ping_storage_data_668 <= (fillup_transition == 1'b1) ? i_input_data[285 % IN_WIDTH] : ping_storage_data_668 ^ i_input_data[285 % IN_WIDTH];
                327 / IN_WIDTH: ping_storage_data_668 <= (fillup_transition == 1'b1) ? i_input_data[327 % IN_WIDTH] : ping_storage_data_668 ^ i_input_data[327 % IN_WIDTH];
                942 / IN_WIDTH: ping_storage_data_668 <= (fillup_transition == 1'b1) ? i_input_data[942 % IN_WIDTH] : ping_storage_data_668 ^ i_input_data[942 % IN_WIDTH];
                1034 / IN_WIDTH: ping_storage_data_668 <= (fillup_transition == 1'b1) ? i_input_data[1034 % IN_WIDTH] : ping_storage_data_668 ^ i_input_data[1034 % IN_WIDTH];
                default: ping_storage_data_668 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_668;
                endcase
            end else begin
                case (input_count)
                285 / IN_WIDTH: pong_storage_data_668 <= (fillup_transition == 1'b1) ? i_input_data[285 % IN_WIDTH] : pong_storage_data_668 ^ i_input_data[285 % IN_WIDTH];
                327 / IN_WIDTH: pong_storage_data_668 <= (fillup_transition == 1'b1) ? i_input_data[327 % IN_WIDTH] : pong_storage_data_668 ^ i_input_data[327 % IN_WIDTH];
                942 / IN_WIDTH: pong_storage_data_668 <= (fillup_transition == 1'b1) ? i_input_data[942 % IN_WIDTH] : pong_storage_data_668 ^ i_input_data[942 % IN_WIDTH];
                1034 / IN_WIDTH: pong_storage_data_668 <= (fillup_transition == 1'b1) ? i_input_data[1034 % IN_WIDTH] : pong_storage_data_668 ^ i_input_data[1034 % IN_WIDTH];
                default: pong_storage_data_668 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_668;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_668 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_668;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_668 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_668;
            end
        end
    end
end

logic ping_storage_data_669;
logic pong_storage_data_669;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_669 <= 1'b0;
        pong_storage_data_669 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                286 / IN_WIDTH: ping_storage_data_669 <= (fillup_transition == 1'b1) ? i_input_data[286 % IN_WIDTH] : ping_storage_data_669 ^ i_input_data[286 % IN_WIDTH];
                328 / IN_WIDTH: ping_storage_data_669 <= (fillup_transition == 1'b1) ? i_input_data[328 % IN_WIDTH] : ping_storage_data_669 ^ i_input_data[328 % IN_WIDTH];
                943 / IN_WIDTH: ping_storage_data_669 <= (fillup_transition == 1'b1) ? i_input_data[943 % IN_WIDTH] : ping_storage_data_669 ^ i_input_data[943 % IN_WIDTH];
                1035 / IN_WIDTH: ping_storage_data_669 <= (fillup_transition == 1'b1) ? i_input_data[1035 % IN_WIDTH] : ping_storage_data_669 ^ i_input_data[1035 % IN_WIDTH];
                default: ping_storage_data_669 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_669;
                endcase
            end else begin
                case (input_count)
                286 / IN_WIDTH: pong_storage_data_669 <= (fillup_transition == 1'b1) ? i_input_data[286 % IN_WIDTH] : pong_storage_data_669 ^ i_input_data[286 % IN_WIDTH];
                328 / IN_WIDTH: pong_storage_data_669 <= (fillup_transition == 1'b1) ? i_input_data[328 % IN_WIDTH] : pong_storage_data_669 ^ i_input_data[328 % IN_WIDTH];
                943 / IN_WIDTH: pong_storage_data_669 <= (fillup_transition == 1'b1) ? i_input_data[943 % IN_WIDTH] : pong_storage_data_669 ^ i_input_data[943 % IN_WIDTH];
                1035 / IN_WIDTH: pong_storage_data_669 <= (fillup_transition == 1'b1) ? i_input_data[1035 % IN_WIDTH] : pong_storage_data_669 ^ i_input_data[1035 % IN_WIDTH];
                default: pong_storage_data_669 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_669;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_669 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_669;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_669 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_669;
            end
        end
    end
end

logic ping_storage_data_670;
logic pong_storage_data_670;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_670 <= 1'b0;
        pong_storage_data_670 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                287 / IN_WIDTH: ping_storage_data_670 <= (fillup_transition == 1'b1) ? i_input_data[287 % IN_WIDTH] : ping_storage_data_670 ^ i_input_data[287 % IN_WIDTH];
                329 / IN_WIDTH: ping_storage_data_670 <= (fillup_transition == 1'b1) ? i_input_data[329 % IN_WIDTH] : ping_storage_data_670 ^ i_input_data[329 % IN_WIDTH];
                944 / IN_WIDTH: ping_storage_data_670 <= (fillup_transition == 1'b1) ? i_input_data[944 % IN_WIDTH] : ping_storage_data_670 ^ i_input_data[944 % IN_WIDTH];
                1036 / IN_WIDTH: ping_storage_data_670 <= (fillup_transition == 1'b1) ? i_input_data[1036 % IN_WIDTH] : ping_storage_data_670 ^ i_input_data[1036 % IN_WIDTH];
                default: ping_storage_data_670 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_670;
                endcase
            end else begin
                case (input_count)
                287 / IN_WIDTH: pong_storage_data_670 <= (fillup_transition == 1'b1) ? i_input_data[287 % IN_WIDTH] : pong_storage_data_670 ^ i_input_data[287 % IN_WIDTH];
                329 / IN_WIDTH: pong_storage_data_670 <= (fillup_transition == 1'b1) ? i_input_data[329 % IN_WIDTH] : pong_storage_data_670 ^ i_input_data[329 % IN_WIDTH];
                944 / IN_WIDTH: pong_storage_data_670 <= (fillup_transition == 1'b1) ? i_input_data[944 % IN_WIDTH] : pong_storage_data_670 ^ i_input_data[944 % IN_WIDTH];
                1036 / IN_WIDTH: pong_storage_data_670 <= (fillup_transition == 1'b1) ? i_input_data[1036 % IN_WIDTH] : pong_storage_data_670 ^ i_input_data[1036 % IN_WIDTH];
                default: pong_storage_data_670 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_670;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_670 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_670;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_670 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_670;
            end
        end
    end
end

logic ping_storage_data_671;
logic pong_storage_data_671;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_671 <= 1'b0;
        pong_storage_data_671 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                192 / IN_WIDTH: ping_storage_data_671 <= (fillup_transition == 1'b1) ? i_input_data[192 % IN_WIDTH] : ping_storage_data_671 ^ i_input_data[192 % IN_WIDTH];
                330 / IN_WIDTH: ping_storage_data_671 <= (fillup_transition == 1'b1) ? i_input_data[330 % IN_WIDTH] : ping_storage_data_671 ^ i_input_data[330 % IN_WIDTH];
                945 / IN_WIDTH: ping_storage_data_671 <= (fillup_transition == 1'b1) ? i_input_data[945 % IN_WIDTH] : ping_storage_data_671 ^ i_input_data[945 % IN_WIDTH];
                1037 / IN_WIDTH: ping_storage_data_671 <= (fillup_transition == 1'b1) ? i_input_data[1037 % IN_WIDTH] : ping_storage_data_671 ^ i_input_data[1037 % IN_WIDTH];
                default: ping_storage_data_671 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_671;
                endcase
            end else begin
                case (input_count)
                192 / IN_WIDTH: pong_storage_data_671 <= (fillup_transition == 1'b1) ? i_input_data[192 % IN_WIDTH] : pong_storage_data_671 ^ i_input_data[192 % IN_WIDTH];
                330 / IN_WIDTH: pong_storage_data_671 <= (fillup_transition == 1'b1) ? i_input_data[330 % IN_WIDTH] : pong_storage_data_671 ^ i_input_data[330 % IN_WIDTH];
                945 / IN_WIDTH: pong_storage_data_671 <= (fillup_transition == 1'b1) ? i_input_data[945 % IN_WIDTH] : pong_storage_data_671 ^ i_input_data[945 % IN_WIDTH];
                1037 / IN_WIDTH: pong_storage_data_671 <= (fillup_transition == 1'b1) ? i_input_data[1037 % IN_WIDTH] : pong_storage_data_671 ^ i_input_data[1037 % IN_WIDTH];
                default: pong_storage_data_671 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_671;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_671 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_671;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_671 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_671;
            end
        end
    end
end

logic ping_storage_data_672;
logic pong_storage_data_672;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_672 <= 1'b0;
        pong_storage_data_672 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                181 / IN_WIDTH: ping_storage_data_672 <= (fillup_transition == 1'b1) ? i_input_data[181 % IN_WIDTH] : ping_storage_data_672 ^ i_input_data[181 % IN_WIDTH];
                215 / IN_WIDTH: ping_storage_data_672 <= (fillup_transition == 1'b1) ? i_input_data[215 % IN_WIDTH] : ping_storage_data_672 ^ i_input_data[215 % IN_WIDTH];
                670 / IN_WIDTH: ping_storage_data_672 <= (fillup_transition == 1'b1) ? i_input_data[670 % IN_WIDTH] : ping_storage_data_672 ^ i_input_data[670 % IN_WIDTH];
                913 / IN_WIDTH: ping_storage_data_672 <= (fillup_transition == 1'b1) ? i_input_data[913 % IN_WIDTH] : ping_storage_data_672 ^ i_input_data[913 % IN_WIDTH];
                default: ping_storage_data_672 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_672;
                endcase
            end else begin
                case (input_count)
                181 / IN_WIDTH: pong_storage_data_672 <= (fillup_transition == 1'b1) ? i_input_data[181 % IN_WIDTH] : pong_storage_data_672 ^ i_input_data[181 % IN_WIDTH];
                215 / IN_WIDTH: pong_storage_data_672 <= (fillup_transition == 1'b1) ? i_input_data[215 % IN_WIDTH] : pong_storage_data_672 ^ i_input_data[215 % IN_WIDTH];
                670 / IN_WIDTH: pong_storage_data_672 <= (fillup_transition == 1'b1) ? i_input_data[670 % IN_WIDTH] : pong_storage_data_672 ^ i_input_data[670 % IN_WIDTH];
                913 / IN_WIDTH: pong_storage_data_672 <= (fillup_transition == 1'b1) ? i_input_data[913 % IN_WIDTH] : pong_storage_data_672 ^ i_input_data[913 % IN_WIDTH];
                default: pong_storage_data_672 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_672;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_672 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_672;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_672 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_672;
            end
        end
    end
end

logic ping_storage_data_673;
logic pong_storage_data_673;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_673 <= 1'b0;
        pong_storage_data_673 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                182 / IN_WIDTH: ping_storage_data_673 <= (fillup_transition == 1'b1) ? i_input_data[182 % IN_WIDTH] : ping_storage_data_673 ^ i_input_data[182 % IN_WIDTH];
                216 / IN_WIDTH: ping_storage_data_673 <= (fillup_transition == 1'b1) ? i_input_data[216 % IN_WIDTH] : ping_storage_data_673 ^ i_input_data[216 % IN_WIDTH];
                671 / IN_WIDTH: ping_storage_data_673 <= (fillup_transition == 1'b1) ? i_input_data[671 % IN_WIDTH] : ping_storage_data_673 ^ i_input_data[671 % IN_WIDTH];
                914 / IN_WIDTH: ping_storage_data_673 <= (fillup_transition == 1'b1) ? i_input_data[914 % IN_WIDTH] : ping_storage_data_673 ^ i_input_data[914 % IN_WIDTH];
                default: ping_storage_data_673 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_673;
                endcase
            end else begin
                case (input_count)
                182 / IN_WIDTH: pong_storage_data_673 <= (fillup_transition == 1'b1) ? i_input_data[182 % IN_WIDTH] : pong_storage_data_673 ^ i_input_data[182 % IN_WIDTH];
                216 / IN_WIDTH: pong_storage_data_673 <= (fillup_transition == 1'b1) ? i_input_data[216 % IN_WIDTH] : pong_storage_data_673 ^ i_input_data[216 % IN_WIDTH];
                671 / IN_WIDTH: pong_storage_data_673 <= (fillup_transition == 1'b1) ? i_input_data[671 % IN_WIDTH] : pong_storage_data_673 ^ i_input_data[671 % IN_WIDTH];
                914 / IN_WIDTH: pong_storage_data_673 <= (fillup_transition == 1'b1) ? i_input_data[914 % IN_WIDTH] : pong_storage_data_673 ^ i_input_data[914 % IN_WIDTH];
                default: pong_storage_data_673 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_673;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_673 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_673;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_673 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_673;
            end
        end
    end
end

logic ping_storage_data_674;
logic pong_storage_data_674;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_674 <= 1'b0;
        pong_storage_data_674 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                183 / IN_WIDTH: ping_storage_data_674 <= (fillup_transition == 1'b1) ? i_input_data[183 % IN_WIDTH] : ping_storage_data_674 ^ i_input_data[183 % IN_WIDTH];
                217 / IN_WIDTH: ping_storage_data_674 <= (fillup_transition == 1'b1) ? i_input_data[217 % IN_WIDTH] : ping_storage_data_674 ^ i_input_data[217 % IN_WIDTH];
                576 / IN_WIDTH: ping_storage_data_674 <= (fillup_transition == 1'b1) ? i_input_data[576 % IN_WIDTH] : ping_storage_data_674 ^ i_input_data[576 % IN_WIDTH];
                915 / IN_WIDTH: ping_storage_data_674 <= (fillup_transition == 1'b1) ? i_input_data[915 % IN_WIDTH] : ping_storage_data_674 ^ i_input_data[915 % IN_WIDTH];
                default: ping_storage_data_674 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_674;
                endcase
            end else begin
                case (input_count)
                183 / IN_WIDTH: pong_storage_data_674 <= (fillup_transition == 1'b1) ? i_input_data[183 % IN_WIDTH] : pong_storage_data_674 ^ i_input_data[183 % IN_WIDTH];
                217 / IN_WIDTH: pong_storage_data_674 <= (fillup_transition == 1'b1) ? i_input_data[217 % IN_WIDTH] : pong_storage_data_674 ^ i_input_data[217 % IN_WIDTH];
                576 / IN_WIDTH: pong_storage_data_674 <= (fillup_transition == 1'b1) ? i_input_data[576 % IN_WIDTH] : pong_storage_data_674 ^ i_input_data[576 % IN_WIDTH];
                915 / IN_WIDTH: pong_storage_data_674 <= (fillup_transition == 1'b1) ? i_input_data[915 % IN_WIDTH] : pong_storage_data_674 ^ i_input_data[915 % IN_WIDTH];
                default: pong_storage_data_674 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_674;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_674 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_674;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_674 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_674;
            end
        end
    end
end

logic ping_storage_data_675;
logic pong_storage_data_675;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_675 <= 1'b0;
        pong_storage_data_675 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                184 / IN_WIDTH: ping_storage_data_675 <= (fillup_transition == 1'b1) ? i_input_data[184 % IN_WIDTH] : ping_storage_data_675 ^ i_input_data[184 % IN_WIDTH];
                218 / IN_WIDTH: ping_storage_data_675 <= (fillup_transition == 1'b1) ? i_input_data[218 % IN_WIDTH] : ping_storage_data_675 ^ i_input_data[218 % IN_WIDTH];
                577 / IN_WIDTH: ping_storage_data_675 <= (fillup_transition == 1'b1) ? i_input_data[577 % IN_WIDTH] : ping_storage_data_675 ^ i_input_data[577 % IN_WIDTH];
                916 / IN_WIDTH: ping_storage_data_675 <= (fillup_transition == 1'b1) ? i_input_data[916 % IN_WIDTH] : ping_storage_data_675 ^ i_input_data[916 % IN_WIDTH];
                default: ping_storage_data_675 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_675;
                endcase
            end else begin
                case (input_count)
                184 / IN_WIDTH: pong_storage_data_675 <= (fillup_transition == 1'b1) ? i_input_data[184 % IN_WIDTH] : pong_storage_data_675 ^ i_input_data[184 % IN_WIDTH];
                218 / IN_WIDTH: pong_storage_data_675 <= (fillup_transition == 1'b1) ? i_input_data[218 % IN_WIDTH] : pong_storage_data_675 ^ i_input_data[218 % IN_WIDTH];
                577 / IN_WIDTH: pong_storage_data_675 <= (fillup_transition == 1'b1) ? i_input_data[577 % IN_WIDTH] : pong_storage_data_675 ^ i_input_data[577 % IN_WIDTH];
                916 / IN_WIDTH: pong_storage_data_675 <= (fillup_transition == 1'b1) ? i_input_data[916 % IN_WIDTH] : pong_storage_data_675 ^ i_input_data[916 % IN_WIDTH];
                default: pong_storage_data_675 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_675;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_675 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_675;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_675 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_675;
            end
        end
    end
end

logic ping_storage_data_676;
logic pong_storage_data_676;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_676 <= 1'b0;
        pong_storage_data_676 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                185 / IN_WIDTH: ping_storage_data_676 <= (fillup_transition == 1'b1) ? i_input_data[185 % IN_WIDTH] : ping_storage_data_676 ^ i_input_data[185 % IN_WIDTH];
                219 / IN_WIDTH: ping_storage_data_676 <= (fillup_transition == 1'b1) ? i_input_data[219 % IN_WIDTH] : ping_storage_data_676 ^ i_input_data[219 % IN_WIDTH];
                578 / IN_WIDTH: ping_storage_data_676 <= (fillup_transition == 1'b1) ? i_input_data[578 % IN_WIDTH] : ping_storage_data_676 ^ i_input_data[578 % IN_WIDTH];
                917 / IN_WIDTH: ping_storage_data_676 <= (fillup_transition == 1'b1) ? i_input_data[917 % IN_WIDTH] : ping_storage_data_676 ^ i_input_data[917 % IN_WIDTH];
                default: ping_storage_data_676 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_676;
                endcase
            end else begin
                case (input_count)
                185 / IN_WIDTH: pong_storage_data_676 <= (fillup_transition == 1'b1) ? i_input_data[185 % IN_WIDTH] : pong_storage_data_676 ^ i_input_data[185 % IN_WIDTH];
                219 / IN_WIDTH: pong_storage_data_676 <= (fillup_transition == 1'b1) ? i_input_data[219 % IN_WIDTH] : pong_storage_data_676 ^ i_input_data[219 % IN_WIDTH];
                578 / IN_WIDTH: pong_storage_data_676 <= (fillup_transition == 1'b1) ? i_input_data[578 % IN_WIDTH] : pong_storage_data_676 ^ i_input_data[578 % IN_WIDTH];
                917 / IN_WIDTH: pong_storage_data_676 <= (fillup_transition == 1'b1) ? i_input_data[917 % IN_WIDTH] : pong_storage_data_676 ^ i_input_data[917 % IN_WIDTH];
                default: pong_storage_data_676 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_676;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_676 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_676;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_676 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_676;
            end
        end
    end
end

logic ping_storage_data_677;
logic pong_storage_data_677;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_677 <= 1'b0;
        pong_storage_data_677 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                186 / IN_WIDTH: ping_storage_data_677 <= (fillup_transition == 1'b1) ? i_input_data[186 % IN_WIDTH] : ping_storage_data_677 ^ i_input_data[186 % IN_WIDTH];
                220 / IN_WIDTH: ping_storage_data_677 <= (fillup_transition == 1'b1) ? i_input_data[220 % IN_WIDTH] : ping_storage_data_677 ^ i_input_data[220 % IN_WIDTH];
                579 / IN_WIDTH: ping_storage_data_677 <= (fillup_transition == 1'b1) ? i_input_data[579 % IN_WIDTH] : ping_storage_data_677 ^ i_input_data[579 % IN_WIDTH];
                918 / IN_WIDTH: ping_storage_data_677 <= (fillup_transition == 1'b1) ? i_input_data[918 % IN_WIDTH] : ping_storage_data_677 ^ i_input_data[918 % IN_WIDTH];
                default: ping_storage_data_677 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_677;
                endcase
            end else begin
                case (input_count)
                186 / IN_WIDTH: pong_storage_data_677 <= (fillup_transition == 1'b1) ? i_input_data[186 % IN_WIDTH] : pong_storage_data_677 ^ i_input_data[186 % IN_WIDTH];
                220 / IN_WIDTH: pong_storage_data_677 <= (fillup_transition == 1'b1) ? i_input_data[220 % IN_WIDTH] : pong_storage_data_677 ^ i_input_data[220 % IN_WIDTH];
                579 / IN_WIDTH: pong_storage_data_677 <= (fillup_transition == 1'b1) ? i_input_data[579 % IN_WIDTH] : pong_storage_data_677 ^ i_input_data[579 % IN_WIDTH];
                918 / IN_WIDTH: pong_storage_data_677 <= (fillup_transition == 1'b1) ? i_input_data[918 % IN_WIDTH] : pong_storage_data_677 ^ i_input_data[918 % IN_WIDTH];
                default: pong_storage_data_677 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_677;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_677 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_677;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_677 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_677;
            end
        end
    end
end

logic ping_storage_data_678;
logic pong_storage_data_678;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_678 <= 1'b0;
        pong_storage_data_678 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                187 / IN_WIDTH: ping_storage_data_678 <= (fillup_transition == 1'b1) ? i_input_data[187 % IN_WIDTH] : ping_storage_data_678 ^ i_input_data[187 % IN_WIDTH];
                221 / IN_WIDTH: ping_storage_data_678 <= (fillup_transition == 1'b1) ? i_input_data[221 % IN_WIDTH] : ping_storage_data_678 ^ i_input_data[221 % IN_WIDTH];
                580 / IN_WIDTH: ping_storage_data_678 <= (fillup_transition == 1'b1) ? i_input_data[580 % IN_WIDTH] : ping_storage_data_678 ^ i_input_data[580 % IN_WIDTH];
                919 / IN_WIDTH: ping_storage_data_678 <= (fillup_transition == 1'b1) ? i_input_data[919 % IN_WIDTH] : ping_storage_data_678 ^ i_input_data[919 % IN_WIDTH];
                default: ping_storage_data_678 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_678;
                endcase
            end else begin
                case (input_count)
                187 / IN_WIDTH: pong_storage_data_678 <= (fillup_transition == 1'b1) ? i_input_data[187 % IN_WIDTH] : pong_storage_data_678 ^ i_input_data[187 % IN_WIDTH];
                221 / IN_WIDTH: pong_storage_data_678 <= (fillup_transition == 1'b1) ? i_input_data[221 % IN_WIDTH] : pong_storage_data_678 ^ i_input_data[221 % IN_WIDTH];
                580 / IN_WIDTH: pong_storage_data_678 <= (fillup_transition == 1'b1) ? i_input_data[580 % IN_WIDTH] : pong_storage_data_678 ^ i_input_data[580 % IN_WIDTH];
                919 / IN_WIDTH: pong_storage_data_678 <= (fillup_transition == 1'b1) ? i_input_data[919 % IN_WIDTH] : pong_storage_data_678 ^ i_input_data[919 % IN_WIDTH];
                default: pong_storage_data_678 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_678;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_678 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_678;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_678 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_678;
            end
        end
    end
end

logic ping_storage_data_679;
logic pong_storage_data_679;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_679 <= 1'b0;
        pong_storage_data_679 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                188 / IN_WIDTH: ping_storage_data_679 <= (fillup_transition == 1'b1) ? i_input_data[188 % IN_WIDTH] : ping_storage_data_679 ^ i_input_data[188 % IN_WIDTH];
                222 / IN_WIDTH: ping_storage_data_679 <= (fillup_transition == 1'b1) ? i_input_data[222 % IN_WIDTH] : ping_storage_data_679 ^ i_input_data[222 % IN_WIDTH];
                581 / IN_WIDTH: ping_storage_data_679 <= (fillup_transition == 1'b1) ? i_input_data[581 % IN_WIDTH] : ping_storage_data_679 ^ i_input_data[581 % IN_WIDTH];
                920 / IN_WIDTH: ping_storage_data_679 <= (fillup_transition == 1'b1) ? i_input_data[920 % IN_WIDTH] : ping_storage_data_679 ^ i_input_data[920 % IN_WIDTH];
                default: ping_storage_data_679 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_679;
                endcase
            end else begin
                case (input_count)
                188 / IN_WIDTH: pong_storage_data_679 <= (fillup_transition == 1'b1) ? i_input_data[188 % IN_WIDTH] : pong_storage_data_679 ^ i_input_data[188 % IN_WIDTH];
                222 / IN_WIDTH: pong_storage_data_679 <= (fillup_transition == 1'b1) ? i_input_data[222 % IN_WIDTH] : pong_storage_data_679 ^ i_input_data[222 % IN_WIDTH];
                581 / IN_WIDTH: pong_storage_data_679 <= (fillup_transition == 1'b1) ? i_input_data[581 % IN_WIDTH] : pong_storage_data_679 ^ i_input_data[581 % IN_WIDTH];
                920 / IN_WIDTH: pong_storage_data_679 <= (fillup_transition == 1'b1) ? i_input_data[920 % IN_WIDTH] : pong_storage_data_679 ^ i_input_data[920 % IN_WIDTH];
                default: pong_storage_data_679 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_679;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_679 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_679;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_679 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_679;
            end
        end
    end
end

logic ping_storage_data_680;
logic pong_storage_data_680;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_680 <= 1'b0;
        pong_storage_data_680 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                189 / IN_WIDTH: ping_storage_data_680 <= (fillup_transition == 1'b1) ? i_input_data[189 % IN_WIDTH] : ping_storage_data_680 ^ i_input_data[189 % IN_WIDTH];
                223 / IN_WIDTH: ping_storage_data_680 <= (fillup_transition == 1'b1) ? i_input_data[223 % IN_WIDTH] : ping_storage_data_680 ^ i_input_data[223 % IN_WIDTH];
                582 / IN_WIDTH: ping_storage_data_680 <= (fillup_transition == 1'b1) ? i_input_data[582 % IN_WIDTH] : ping_storage_data_680 ^ i_input_data[582 % IN_WIDTH];
                921 / IN_WIDTH: ping_storage_data_680 <= (fillup_transition == 1'b1) ? i_input_data[921 % IN_WIDTH] : ping_storage_data_680 ^ i_input_data[921 % IN_WIDTH];
                default: ping_storage_data_680 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_680;
                endcase
            end else begin
                case (input_count)
                189 / IN_WIDTH: pong_storage_data_680 <= (fillup_transition == 1'b1) ? i_input_data[189 % IN_WIDTH] : pong_storage_data_680 ^ i_input_data[189 % IN_WIDTH];
                223 / IN_WIDTH: pong_storage_data_680 <= (fillup_transition == 1'b1) ? i_input_data[223 % IN_WIDTH] : pong_storage_data_680 ^ i_input_data[223 % IN_WIDTH];
                582 / IN_WIDTH: pong_storage_data_680 <= (fillup_transition == 1'b1) ? i_input_data[582 % IN_WIDTH] : pong_storage_data_680 ^ i_input_data[582 % IN_WIDTH];
                921 / IN_WIDTH: pong_storage_data_680 <= (fillup_transition == 1'b1) ? i_input_data[921 % IN_WIDTH] : pong_storage_data_680 ^ i_input_data[921 % IN_WIDTH];
                default: pong_storage_data_680 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_680;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_680 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_680;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_680 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_680;
            end
        end
    end
end

logic ping_storage_data_681;
logic pong_storage_data_681;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_681 <= 1'b0;
        pong_storage_data_681 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                190 / IN_WIDTH: ping_storage_data_681 <= (fillup_transition == 1'b1) ? i_input_data[190 % IN_WIDTH] : ping_storage_data_681 ^ i_input_data[190 % IN_WIDTH];
                224 / IN_WIDTH: ping_storage_data_681 <= (fillup_transition == 1'b1) ? i_input_data[224 % IN_WIDTH] : ping_storage_data_681 ^ i_input_data[224 % IN_WIDTH];
                583 / IN_WIDTH: ping_storage_data_681 <= (fillup_transition == 1'b1) ? i_input_data[583 % IN_WIDTH] : ping_storage_data_681 ^ i_input_data[583 % IN_WIDTH];
                922 / IN_WIDTH: ping_storage_data_681 <= (fillup_transition == 1'b1) ? i_input_data[922 % IN_WIDTH] : ping_storage_data_681 ^ i_input_data[922 % IN_WIDTH];
                default: ping_storage_data_681 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_681;
                endcase
            end else begin
                case (input_count)
                190 / IN_WIDTH: pong_storage_data_681 <= (fillup_transition == 1'b1) ? i_input_data[190 % IN_WIDTH] : pong_storage_data_681 ^ i_input_data[190 % IN_WIDTH];
                224 / IN_WIDTH: pong_storage_data_681 <= (fillup_transition == 1'b1) ? i_input_data[224 % IN_WIDTH] : pong_storage_data_681 ^ i_input_data[224 % IN_WIDTH];
                583 / IN_WIDTH: pong_storage_data_681 <= (fillup_transition == 1'b1) ? i_input_data[583 % IN_WIDTH] : pong_storage_data_681 ^ i_input_data[583 % IN_WIDTH];
                922 / IN_WIDTH: pong_storage_data_681 <= (fillup_transition == 1'b1) ? i_input_data[922 % IN_WIDTH] : pong_storage_data_681 ^ i_input_data[922 % IN_WIDTH];
                default: pong_storage_data_681 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_681;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_681 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_681;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_681 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_681;
            end
        end
    end
end

logic ping_storage_data_682;
logic pong_storage_data_682;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_682 <= 1'b0;
        pong_storage_data_682 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                191 / IN_WIDTH: ping_storage_data_682 <= (fillup_transition == 1'b1) ? i_input_data[191 % IN_WIDTH] : ping_storage_data_682 ^ i_input_data[191 % IN_WIDTH];
                225 / IN_WIDTH: ping_storage_data_682 <= (fillup_transition == 1'b1) ? i_input_data[225 % IN_WIDTH] : ping_storage_data_682 ^ i_input_data[225 % IN_WIDTH];
                584 / IN_WIDTH: ping_storage_data_682 <= (fillup_transition == 1'b1) ? i_input_data[584 % IN_WIDTH] : ping_storage_data_682 ^ i_input_data[584 % IN_WIDTH];
                923 / IN_WIDTH: ping_storage_data_682 <= (fillup_transition == 1'b1) ? i_input_data[923 % IN_WIDTH] : ping_storage_data_682 ^ i_input_data[923 % IN_WIDTH];
                default: ping_storage_data_682 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_682;
                endcase
            end else begin
                case (input_count)
                191 / IN_WIDTH: pong_storage_data_682 <= (fillup_transition == 1'b1) ? i_input_data[191 % IN_WIDTH] : pong_storage_data_682 ^ i_input_data[191 % IN_WIDTH];
                225 / IN_WIDTH: pong_storage_data_682 <= (fillup_transition == 1'b1) ? i_input_data[225 % IN_WIDTH] : pong_storage_data_682 ^ i_input_data[225 % IN_WIDTH];
                584 / IN_WIDTH: pong_storage_data_682 <= (fillup_transition == 1'b1) ? i_input_data[584 % IN_WIDTH] : pong_storage_data_682 ^ i_input_data[584 % IN_WIDTH];
                923 / IN_WIDTH: pong_storage_data_682 <= (fillup_transition == 1'b1) ? i_input_data[923 % IN_WIDTH] : pong_storage_data_682 ^ i_input_data[923 % IN_WIDTH];
                default: pong_storage_data_682 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_682;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_682 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_682;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_682 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_682;
            end
        end
    end
end

logic ping_storage_data_683;
logic pong_storage_data_683;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_683 <= 1'b0;
        pong_storage_data_683 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                96 / IN_WIDTH: ping_storage_data_683 <= (fillup_transition == 1'b1) ? i_input_data[96 % IN_WIDTH] : ping_storage_data_683 ^ i_input_data[96 % IN_WIDTH];
                226 / IN_WIDTH: ping_storage_data_683 <= (fillup_transition == 1'b1) ? i_input_data[226 % IN_WIDTH] : ping_storage_data_683 ^ i_input_data[226 % IN_WIDTH];
                585 / IN_WIDTH: ping_storage_data_683 <= (fillup_transition == 1'b1) ? i_input_data[585 % IN_WIDTH] : ping_storage_data_683 ^ i_input_data[585 % IN_WIDTH];
                924 / IN_WIDTH: ping_storage_data_683 <= (fillup_transition == 1'b1) ? i_input_data[924 % IN_WIDTH] : ping_storage_data_683 ^ i_input_data[924 % IN_WIDTH];
                default: ping_storage_data_683 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_683;
                endcase
            end else begin
                case (input_count)
                96 / IN_WIDTH: pong_storage_data_683 <= (fillup_transition == 1'b1) ? i_input_data[96 % IN_WIDTH] : pong_storage_data_683 ^ i_input_data[96 % IN_WIDTH];
                226 / IN_WIDTH: pong_storage_data_683 <= (fillup_transition == 1'b1) ? i_input_data[226 % IN_WIDTH] : pong_storage_data_683 ^ i_input_data[226 % IN_WIDTH];
                585 / IN_WIDTH: pong_storage_data_683 <= (fillup_transition == 1'b1) ? i_input_data[585 % IN_WIDTH] : pong_storage_data_683 ^ i_input_data[585 % IN_WIDTH];
                924 / IN_WIDTH: pong_storage_data_683 <= (fillup_transition == 1'b1) ? i_input_data[924 % IN_WIDTH] : pong_storage_data_683 ^ i_input_data[924 % IN_WIDTH];
                default: pong_storage_data_683 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_683;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_683 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_683;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_683 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_683;
            end
        end
    end
end

logic ping_storage_data_684;
logic pong_storage_data_684;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_684 <= 1'b0;
        pong_storage_data_684 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                97 / IN_WIDTH: ping_storage_data_684 <= (fillup_transition == 1'b1) ? i_input_data[97 % IN_WIDTH] : ping_storage_data_684 ^ i_input_data[97 % IN_WIDTH];
                227 / IN_WIDTH: ping_storage_data_684 <= (fillup_transition == 1'b1) ? i_input_data[227 % IN_WIDTH] : ping_storage_data_684 ^ i_input_data[227 % IN_WIDTH];
                586 / IN_WIDTH: ping_storage_data_684 <= (fillup_transition == 1'b1) ? i_input_data[586 % IN_WIDTH] : ping_storage_data_684 ^ i_input_data[586 % IN_WIDTH];
                925 / IN_WIDTH: ping_storage_data_684 <= (fillup_transition == 1'b1) ? i_input_data[925 % IN_WIDTH] : ping_storage_data_684 ^ i_input_data[925 % IN_WIDTH];
                default: ping_storage_data_684 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_684;
                endcase
            end else begin
                case (input_count)
                97 / IN_WIDTH: pong_storage_data_684 <= (fillup_transition == 1'b1) ? i_input_data[97 % IN_WIDTH] : pong_storage_data_684 ^ i_input_data[97 % IN_WIDTH];
                227 / IN_WIDTH: pong_storage_data_684 <= (fillup_transition == 1'b1) ? i_input_data[227 % IN_WIDTH] : pong_storage_data_684 ^ i_input_data[227 % IN_WIDTH];
                586 / IN_WIDTH: pong_storage_data_684 <= (fillup_transition == 1'b1) ? i_input_data[586 % IN_WIDTH] : pong_storage_data_684 ^ i_input_data[586 % IN_WIDTH];
                925 / IN_WIDTH: pong_storage_data_684 <= (fillup_transition == 1'b1) ? i_input_data[925 % IN_WIDTH] : pong_storage_data_684 ^ i_input_data[925 % IN_WIDTH];
                default: pong_storage_data_684 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_684;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_684 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_684;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_684 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_684;
            end
        end
    end
end

logic ping_storage_data_685;
logic pong_storage_data_685;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_685 <= 1'b0;
        pong_storage_data_685 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                98 / IN_WIDTH: ping_storage_data_685 <= (fillup_transition == 1'b1) ? i_input_data[98 % IN_WIDTH] : ping_storage_data_685 ^ i_input_data[98 % IN_WIDTH];
                228 / IN_WIDTH: ping_storage_data_685 <= (fillup_transition == 1'b1) ? i_input_data[228 % IN_WIDTH] : ping_storage_data_685 ^ i_input_data[228 % IN_WIDTH];
                587 / IN_WIDTH: ping_storage_data_685 <= (fillup_transition == 1'b1) ? i_input_data[587 % IN_WIDTH] : ping_storage_data_685 ^ i_input_data[587 % IN_WIDTH];
                926 / IN_WIDTH: ping_storage_data_685 <= (fillup_transition == 1'b1) ? i_input_data[926 % IN_WIDTH] : ping_storage_data_685 ^ i_input_data[926 % IN_WIDTH];
                default: ping_storage_data_685 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_685;
                endcase
            end else begin
                case (input_count)
                98 / IN_WIDTH: pong_storage_data_685 <= (fillup_transition == 1'b1) ? i_input_data[98 % IN_WIDTH] : pong_storage_data_685 ^ i_input_data[98 % IN_WIDTH];
                228 / IN_WIDTH: pong_storage_data_685 <= (fillup_transition == 1'b1) ? i_input_data[228 % IN_WIDTH] : pong_storage_data_685 ^ i_input_data[228 % IN_WIDTH];
                587 / IN_WIDTH: pong_storage_data_685 <= (fillup_transition == 1'b1) ? i_input_data[587 % IN_WIDTH] : pong_storage_data_685 ^ i_input_data[587 % IN_WIDTH];
                926 / IN_WIDTH: pong_storage_data_685 <= (fillup_transition == 1'b1) ? i_input_data[926 % IN_WIDTH] : pong_storage_data_685 ^ i_input_data[926 % IN_WIDTH];
                default: pong_storage_data_685 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_685;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_685 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_685;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_685 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_685;
            end
        end
    end
end

logic ping_storage_data_686;
logic pong_storage_data_686;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_686 <= 1'b0;
        pong_storage_data_686 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                99 / IN_WIDTH: ping_storage_data_686 <= (fillup_transition == 1'b1) ? i_input_data[99 % IN_WIDTH] : ping_storage_data_686 ^ i_input_data[99 % IN_WIDTH];
                229 / IN_WIDTH: ping_storage_data_686 <= (fillup_transition == 1'b1) ? i_input_data[229 % IN_WIDTH] : ping_storage_data_686 ^ i_input_data[229 % IN_WIDTH];
                588 / IN_WIDTH: ping_storage_data_686 <= (fillup_transition == 1'b1) ? i_input_data[588 % IN_WIDTH] : ping_storage_data_686 ^ i_input_data[588 % IN_WIDTH];
                927 / IN_WIDTH: ping_storage_data_686 <= (fillup_transition == 1'b1) ? i_input_data[927 % IN_WIDTH] : ping_storage_data_686 ^ i_input_data[927 % IN_WIDTH];
                default: ping_storage_data_686 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_686;
                endcase
            end else begin
                case (input_count)
                99 / IN_WIDTH: pong_storage_data_686 <= (fillup_transition == 1'b1) ? i_input_data[99 % IN_WIDTH] : pong_storage_data_686 ^ i_input_data[99 % IN_WIDTH];
                229 / IN_WIDTH: pong_storage_data_686 <= (fillup_transition == 1'b1) ? i_input_data[229 % IN_WIDTH] : pong_storage_data_686 ^ i_input_data[229 % IN_WIDTH];
                588 / IN_WIDTH: pong_storage_data_686 <= (fillup_transition == 1'b1) ? i_input_data[588 % IN_WIDTH] : pong_storage_data_686 ^ i_input_data[588 % IN_WIDTH];
                927 / IN_WIDTH: pong_storage_data_686 <= (fillup_transition == 1'b1) ? i_input_data[927 % IN_WIDTH] : pong_storage_data_686 ^ i_input_data[927 % IN_WIDTH];
                default: pong_storage_data_686 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_686;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_686 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_686;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_686 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_686;
            end
        end
    end
end

logic ping_storage_data_687;
logic pong_storage_data_687;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_687 <= 1'b0;
        pong_storage_data_687 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                100 / IN_WIDTH: ping_storage_data_687 <= (fillup_transition == 1'b1) ? i_input_data[100 % IN_WIDTH] : ping_storage_data_687 ^ i_input_data[100 % IN_WIDTH];
                230 / IN_WIDTH: ping_storage_data_687 <= (fillup_transition == 1'b1) ? i_input_data[230 % IN_WIDTH] : ping_storage_data_687 ^ i_input_data[230 % IN_WIDTH];
                589 / IN_WIDTH: ping_storage_data_687 <= (fillup_transition == 1'b1) ? i_input_data[589 % IN_WIDTH] : ping_storage_data_687 ^ i_input_data[589 % IN_WIDTH];
                928 / IN_WIDTH: ping_storage_data_687 <= (fillup_transition == 1'b1) ? i_input_data[928 % IN_WIDTH] : ping_storage_data_687 ^ i_input_data[928 % IN_WIDTH];
                default: ping_storage_data_687 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_687;
                endcase
            end else begin
                case (input_count)
                100 / IN_WIDTH: pong_storage_data_687 <= (fillup_transition == 1'b1) ? i_input_data[100 % IN_WIDTH] : pong_storage_data_687 ^ i_input_data[100 % IN_WIDTH];
                230 / IN_WIDTH: pong_storage_data_687 <= (fillup_transition == 1'b1) ? i_input_data[230 % IN_WIDTH] : pong_storage_data_687 ^ i_input_data[230 % IN_WIDTH];
                589 / IN_WIDTH: pong_storage_data_687 <= (fillup_transition == 1'b1) ? i_input_data[589 % IN_WIDTH] : pong_storage_data_687 ^ i_input_data[589 % IN_WIDTH];
                928 / IN_WIDTH: pong_storage_data_687 <= (fillup_transition == 1'b1) ? i_input_data[928 % IN_WIDTH] : pong_storage_data_687 ^ i_input_data[928 % IN_WIDTH];
                default: pong_storage_data_687 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_687;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_687 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_687;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_687 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_687;
            end
        end
    end
end

logic ping_storage_data_688;
logic pong_storage_data_688;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_688 <= 1'b0;
        pong_storage_data_688 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                101 / IN_WIDTH: ping_storage_data_688 <= (fillup_transition == 1'b1) ? i_input_data[101 % IN_WIDTH] : ping_storage_data_688 ^ i_input_data[101 % IN_WIDTH];
                231 / IN_WIDTH: ping_storage_data_688 <= (fillup_transition == 1'b1) ? i_input_data[231 % IN_WIDTH] : ping_storage_data_688 ^ i_input_data[231 % IN_WIDTH];
                590 / IN_WIDTH: ping_storage_data_688 <= (fillup_transition == 1'b1) ? i_input_data[590 % IN_WIDTH] : ping_storage_data_688 ^ i_input_data[590 % IN_WIDTH];
                929 / IN_WIDTH: ping_storage_data_688 <= (fillup_transition == 1'b1) ? i_input_data[929 % IN_WIDTH] : ping_storage_data_688 ^ i_input_data[929 % IN_WIDTH];
                default: ping_storage_data_688 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_688;
                endcase
            end else begin
                case (input_count)
                101 / IN_WIDTH: pong_storage_data_688 <= (fillup_transition == 1'b1) ? i_input_data[101 % IN_WIDTH] : pong_storage_data_688 ^ i_input_data[101 % IN_WIDTH];
                231 / IN_WIDTH: pong_storage_data_688 <= (fillup_transition == 1'b1) ? i_input_data[231 % IN_WIDTH] : pong_storage_data_688 ^ i_input_data[231 % IN_WIDTH];
                590 / IN_WIDTH: pong_storage_data_688 <= (fillup_transition == 1'b1) ? i_input_data[590 % IN_WIDTH] : pong_storage_data_688 ^ i_input_data[590 % IN_WIDTH];
                929 / IN_WIDTH: pong_storage_data_688 <= (fillup_transition == 1'b1) ? i_input_data[929 % IN_WIDTH] : pong_storage_data_688 ^ i_input_data[929 % IN_WIDTH];
                default: pong_storage_data_688 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_688;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_688 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_688;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_688 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_688;
            end
        end
    end
end

logic ping_storage_data_689;
logic pong_storage_data_689;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_689 <= 1'b0;
        pong_storage_data_689 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                102 / IN_WIDTH: ping_storage_data_689 <= (fillup_transition == 1'b1) ? i_input_data[102 % IN_WIDTH] : ping_storage_data_689 ^ i_input_data[102 % IN_WIDTH];
                232 / IN_WIDTH: ping_storage_data_689 <= (fillup_transition == 1'b1) ? i_input_data[232 % IN_WIDTH] : ping_storage_data_689 ^ i_input_data[232 % IN_WIDTH];
                591 / IN_WIDTH: ping_storage_data_689 <= (fillup_transition == 1'b1) ? i_input_data[591 % IN_WIDTH] : ping_storage_data_689 ^ i_input_data[591 % IN_WIDTH];
                930 / IN_WIDTH: ping_storage_data_689 <= (fillup_transition == 1'b1) ? i_input_data[930 % IN_WIDTH] : ping_storage_data_689 ^ i_input_data[930 % IN_WIDTH];
                default: ping_storage_data_689 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_689;
                endcase
            end else begin
                case (input_count)
                102 / IN_WIDTH: pong_storage_data_689 <= (fillup_transition == 1'b1) ? i_input_data[102 % IN_WIDTH] : pong_storage_data_689 ^ i_input_data[102 % IN_WIDTH];
                232 / IN_WIDTH: pong_storage_data_689 <= (fillup_transition == 1'b1) ? i_input_data[232 % IN_WIDTH] : pong_storage_data_689 ^ i_input_data[232 % IN_WIDTH];
                591 / IN_WIDTH: pong_storage_data_689 <= (fillup_transition == 1'b1) ? i_input_data[591 % IN_WIDTH] : pong_storage_data_689 ^ i_input_data[591 % IN_WIDTH];
                930 / IN_WIDTH: pong_storage_data_689 <= (fillup_transition == 1'b1) ? i_input_data[930 % IN_WIDTH] : pong_storage_data_689 ^ i_input_data[930 % IN_WIDTH];
                default: pong_storage_data_689 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_689;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_689 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_689;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_689 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_689;
            end
        end
    end
end

logic ping_storage_data_690;
logic pong_storage_data_690;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_690 <= 1'b0;
        pong_storage_data_690 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                103 / IN_WIDTH: ping_storage_data_690 <= (fillup_transition == 1'b1) ? i_input_data[103 % IN_WIDTH] : ping_storage_data_690 ^ i_input_data[103 % IN_WIDTH];
                233 / IN_WIDTH: ping_storage_data_690 <= (fillup_transition == 1'b1) ? i_input_data[233 % IN_WIDTH] : ping_storage_data_690 ^ i_input_data[233 % IN_WIDTH];
                592 / IN_WIDTH: ping_storage_data_690 <= (fillup_transition == 1'b1) ? i_input_data[592 % IN_WIDTH] : ping_storage_data_690 ^ i_input_data[592 % IN_WIDTH];
                931 / IN_WIDTH: ping_storage_data_690 <= (fillup_transition == 1'b1) ? i_input_data[931 % IN_WIDTH] : ping_storage_data_690 ^ i_input_data[931 % IN_WIDTH];
                default: ping_storage_data_690 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_690;
                endcase
            end else begin
                case (input_count)
                103 / IN_WIDTH: pong_storage_data_690 <= (fillup_transition == 1'b1) ? i_input_data[103 % IN_WIDTH] : pong_storage_data_690 ^ i_input_data[103 % IN_WIDTH];
                233 / IN_WIDTH: pong_storage_data_690 <= (fillup_transition == 1'b1) ? i_input_data[233 % IN_WIDTH] : pong_storage_data_690 ^ i_input_data[233 % IN_WIDTH];
                592 / IN_WIDTH: pong_storage_data_690 <= (fillup_transition == 1'b1) ? i_input_data[592 % IN_WIDTH] : pong_storage_data_690 ^ i_input_data[592 % IN_WIDTH];
                931 / IN_WIDTH: pong_storage_data_690 <= (fillup_transition == 1'b1) ? i_input_data[931 % IN_WIDTH] : pong_storage_data_690 ^ i_input_data[931 % IN_WIDTH];
                default: pong_storage_data_690 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_690;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_690 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_690;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_690 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_690;
            end
        end
    end
end

logic ping_storage_data_691;
logic pong_storage_data_691;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_691 <= 1'b0;
        pong_storage_data_691 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                104 / IN_WIDTH: ping_storage_data_691 <= (fillup_transition == 1'b1) ? i_input_data[104 % IN_WIDTH] : ping_storage_data_691 ^ i_input_data[104 % IN_WIDTH];
                234 / IN_WIDTH: ping_storage_data_691 <= (fillup_transition == 1'b1) ? i_input_data[234 % IN_WIDTH] : ping_storage_data_691 ^ i_input_data[234 % IN_WIDTH];
                593 / IN_WIDTH: ping_storage_data_691 <= (fillup_transition == 1'b1) ? i_input_data[593 % IN_WIDTH] : ping_storage_data_691 ^ i_input_data[593 % IN_WIDTH];
                932 / IN_WIDTH: ping_storage_data_691 <= (fillup_transition == 1'b1) ? i_input_data[932 % IN_WIDTH] : ping_storage_data_691 ^ i_input_data[932 % IN_WIDTH];
                default: ping_storage_data_691 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_691;
                endcase
            end else begin
                case (input_count)
                104 / IN_WIDTH: pong_storage_data_691 <= (fillup_transition == 1'b1) ? i_input_data[104 % IN_WIDTH] : pong_storage_data_691 ^ i_input_data[104 % IN_WIDTH];
                234 / IN_WIDTH: pong_storage_data_691 <= (fillup_transition == 1'b1) ? i_input_data[234 % IN_WIDTH] : pong_storage_data_691 ^ i_input_data[234 % IN_WIDTH];
                593 / IN_WIDTH: pong_storage_data_691 <= (fillup_transition == 1'b1) ? i_input_data[593 % IN_WIDTH] : pong_storage_data_691 ^ i_input_data[593 % IN_WIDTH];
                932 / IN_WIDTH: pong_storage_data_691 <= (fillup_transition == 1'b1) ? i_input_data[932 % IN_WIDTH] : pong_storage_data_691 ^ i_input_data[932 % IN_WIDTH];
                default: pong_storage_data_691 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_691;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_691 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_691;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_691 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_691;
            end
        end
    end
end

logic ping_storage_data_692;
logic pong_storage_data_692;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_692 <= 1'b0;
        pong_storage_data_692 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                105 / IN_WIDTH: ping_storage_data_692 <= (fillup_transition == 1'b1) ? i_input_data[105 % IN_WIDTH] : ping_storage_data_692 ^ i_input_data[105 % IN_WIDTH];
                235 / IN_WIDTH: ping_storage_data_692 <= (fillup_transition == 1'b1) ? i_input_data[235 % IN_WIDTH] : ping_storage_data_692 ^ i_input_data[235 % IN_WIDTH];
                594 / IN_WIDTH: ping_storage_data_692 <= (fillup_transition == 1'b1) ? i_input_data[594 % IN_WIDTH] : ping_storage_data_692 ^ i_input_data[594 % IN_WIDTH];
                933 / IN_WIDTH: ping_storage_data_692 <= (fillup_transition == 1'b1) ? i_input_data[933 % IN_WIDTH] : ping_storage_data_692 ^ i_input_data[933 % IN_WIDTH];
                default: ping_storage_data_692 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_692;
                endcase
            end else begin
                case (input_count)
                105 / IN_WIDTH: pong_storage_data_692 <= (fillup_transition == 1'b1) ? i_input_data[105 % IN_WIDTH] : pong_storage_data_692 ^ i_input_data[105 % IN_WIDTH];
                235 / IN_WIDTH: pong_storage_data_692 <= (fillup_transition == 1'b1) ? i_input_data[235 % IN_WIDTH] : pong_storage_data_692 ^ i_input_data[235 % IN_WIDTH];
                594 / IN_WIDTH: pong_storage_data_692 <= (fillup_transition == 1'b1) ? i_input_data[594 % IN_WIDTH] : pong_storage_data_692 ^ i_input_data[594 % IN_WIDTH];
                933 / IN_WIDTH: pong_storage_data_692 <= (fillup_transition == 1'b1) ? i_input_data[933 % IN_WIDTH] : pong_storage_data_692 ^ i_input_data[933 % IN_WIDTH];
                default: pong_storage_data_692 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_692;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_692 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_692;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_692 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_692;
            end
        end
    end
end

logic ping_storage_data_693;
logic pong_storage_data_693;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_693 <= 1'b0;
        pong_storage_data_693 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                106 / IN_WIDTH: ping_storage_data_693 <= (fillup_transition == 1'b1) ? i_input_data[106 % IN_WIDTH] : ping_storage_data_693 ^ i_input_data[106 % IN_WIDTH];
                236 / IN_WIDTH: ping_storage_data_693 <= (fillup_transition == 1'b1) ? i_input_data[236 % IN_WIDTH] : ping_storage_data_693 ^ i_input_data[236 % IN_WIDTH];
                595 / IN_WIDTH: ping_storage_data_693 <= (fillup_transition == 1'b1) ? i_input_data[595 % IN_WIDTH] : ping_storage_data_693 ^ i_input_data[595 % IN_WIDTH];
                934 / IN_WIDTH: ping_storage_data_693 <= (fillup_transition == 1'b1) ? i_input_data[934 % IN_WIDTH] : ping_storage_data_693 ^ i_input_data[934 % IN_WIDTH];
                default: ping_storage_data_693 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_693;
                endcase
            end else begin
                case (input_count)
                106 / IN_WIDTH: pong_storage_data_693 <= (fillup_transition == 1'b1) ? i_input_data[106 % IN_WIDTH] : pong_storage_data_693 ^ i_input_data[106 % IN_WIDTH];
                236 / IN_WIDTH: pong_storage_data_693 <= (fillup_transition == 1'b1) ? i_input_data[236 % IN_WIDTH] : pong_storage_data_693 ^ i_input_data[236 % IN_WIDTH];
                595 / IN_WIDTH: pong_storage_data_693 <= (fillup_transition == 1'b1) ? i_input_data[595 % IN_WIDTH] : pong_storage_data_693 ^ i_input_data[595 % IN_WIDTH];
                934 / IN_WIDTH: pong_storage_data_693 <= (fillup_transition == 1'b1) ? i_input_data[934 % IN_WIDTH] : pong_storage_data_693 ^ i_input_data[934 % IN_WIDTH];
                default: pong_storage_data_693 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_693;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_693 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_693;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_693 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_693;
            end
        end
    end
end

logic ping_storage_data_694;
logic pong_storage_data_694;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_694 <= 1'b0;
        pong_storage_data_694 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                107 / IN_WIDTH: ping_storage_data_694 <= (fillup_transition == 1'b1) ? i_input_data[107 % IN_WIDTH] : ping_storage_data_694 ^ i_input_data[107 % IN_WIDTH];
                237 / IN_WIDTH: ping_storage_data_694 <= (fillup_transition == 1'b1) ? i_input_data[237 % IN_WIDTH] : ping_storage_data_694 ^ i_input_data[237 % IN_WIDTH];
                596 / IN_WIDTH: ping_storage_data_694 <= (fillup_transition == 1'b1) ? i_input_data[596 % IN_WIDTH] : ping_storage_data_694 ^ i_input_data[596 % IN_WIDTH];
                935 / IN_WIDTH: ping_storage_data_694 <= (fillup_transition == 1'b1) ? i_input_data[935 % IN_WIDTH] : ping_storage_data_694 ^ i_input_data[935 % IN_WIDTH];
                default: ping_storage_data_694 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_694;
                endcase
            end else begin
                case (input_count)
                107 / IN_WIDTH: pong_storage_data_694 <= (fillup_transition == 1'b1) ? i_input_data[107 % IN_WIDTH] : pong_storage_data_694 ^ i_input_data[107 % IN_WIDTH];
                237 / IN_WIDTH: pong_storage_data_694 <= (fillup_transition == 1'b1) ? i_input_data[237 % IN_WIDTH] : pong_storage_data_694 ^ i_input_data[237 % IN_WIDTH];
                596 / IN_WIDTH: pong_storage_data_694 <= (fillup_transition == 1'b1) ? i_input_data[596 % IN_WIDTH] : pong_storage_data_694 ^ i_input_data[596 % IN_WIDTH];
                935 / IN_WIDTH: pong_storage_data_694 <= (fillup_transition == 1'b1) ? i_input_data[935 % IN_WIDTH] : pong_storage_data_694 ^ i_input_data[935 % IN_WIDTH];
                default: pong_storage_data_694 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_694;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_694 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_694;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_694 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_694;
            end
        end
    end
end

logic ping_storage_data_695;
logic pong_storage_data_695;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_695 <= 1'b0;
        pong_storage_data_695 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                108 / IN_WIDTH: ping_storage_data_695 <= (fillup_transition == 1'b1) ? i_input_data[108 % IN_WIDTH] : ping_storage_data_695 ^ i_input_data[108 % IN_WIDTH];
                238 / IN_WIDTH: ping_storage_data_695 <= (fillup_transition == 1'b1) ? i_input_data[238 % IN_WIDTH] : ping_storage_data_695 ^ i_input_data[238 % IN_WIDTH];
                597 / IN_WIDTH: ping_storage_data_695 <= (fillup_transition == 1'b1) ? i_input_data[597 % IN_WIDTH] : ping_storage_data_695 ^ i_input_data[597 % IN_WIDTH];
                936 / IN_WIDTH: ping_storage_data_695 <= (fillup_transition == 1'b1) ? i_input_data[936 % IN_WIDTH] : ping_storage_data_695 ^ i_input_data[936 % IN_WIDTH];
                default: ping_storage_data_695 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_695;
                endcase
            end else begin
                case (input_count)
                108 / IN_WIDTH: pong_storage_data_695 <= (fillup_transition == 1'b1) ? i_input_data[108 % IN_WIDTH] : pong_storage_data_695 ^ i_input_data[108 % IN_WIDTH];
                238 / IN_WIDTH: pong_storage_data_695 <= (fillup_transition == 1'b1) ? i_input_data[238 % IN_WIDTH] : pong_storage_data_695 ^ i_input_data[238 % IN_WIDTH];
                597 / IN_WIDTH: pong_storage_data_695 <= (fillup_transition == 1'b1) ? i_input_data[597 % IN_WIDTH] : pong_storage_data_695 ^ i_input_data[597 % IN_WIDTH];
                936 / IN_WIDTH: pong_storage_data_695 <= (fillup_transition == 1'b1) ? i_input_data[936 % IN_WIDTH] : pong_storage_data_695 ^ i_input_data[936 % IN_WIDTH];
                default: pong_storage_data_695 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_695;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_695 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_695;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_695 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_695;
            end
        end
    end
end

logic ping_storage_data_696;
logic pong_storage_data_696;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_696 <= 1'b0;
        pong_storage_data_696 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                109 / IN_WIDTH: ping_storage_data_696 <= (fillup_transition == 1'b1) ? i_input_data[109 % IN_WIDTH] : ping_storage_data_696 ^ i_input_data[109 % IN_WIDTH];
                239 / IN_WIDTH: ping_storage_data_696 <= (fillup_transition == 1'b1) ? i_input_data[239 % IN_WIDTH] : ping_storage_data_696 ^ i_input_data[239 % IN_WIDTH];
                598 / IN_WIDTH: ping_storage_data_696 <= (fillup_transition == 1'b1) ? i_input_data[598 % IN_WIDTH] : ping_storage_data_696 ^ i_input_data[598 % IN_WIDTH];
                937 / IN_WIDTH: ping_storage_data_696 <= (fillup_transition == 1'b1) ? i_input_data[937 % IN_WIDTH] : ping_storage_data_696 ^ i_input_data[937 % IN_WIDTH];
                default: ping_storage_data_696 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_696;
                endcase
            end else begin
                case (input_count)
                109 / IN_WIDTH: pong_storage_data_696 <= (fillup_transition == 1'b1) ? i_input_data[109 % IN_WIDTH] : pong_storage_data_696 ^ i_input_data[109 % IN_WIDTH];
                239 / IN_WIDTH: pong_storage_data_696 <= (fillup_transition == 1'b1) ? i_input_data[239 % IN_WIDTH] : pong_storage_data_696 ^ i_input_data[239 % IN_WIDTH];
                598 / IN_WIDTH: pong_storage_data_696 <= (fillup_transition == 1'b1) ? i_input_data[598 % IN_WIDTH] : pong_storage_data_696 ^ i_input_data[598 % IN_WIDTH];
                937 / IN_WIDTH: pong_storage_data_696 <= (fillup_transition == 1'b1) ? i_input_data[937 % IN_WIDTH] : pong_storage_data_696 ^ i_input_data[937 % IN_WIDTH];
                default: pong_storage_data_696 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_696;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_696 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_696;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_696 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_696;
            end
        end
    end
end

logic ping_storage_data_697;
logic pong_storage_data_697;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_697 <= 1'b0;
        pong_storage_data_697 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                110 / IN_WIDTH: ping_storage_data_697 <= (fillup_transition == 1'b1) ? i_input_data[110 % IN_WIDTH] : ping_storage_data_697 ^ i_input_data[110 % IN_WIDTH];
                240 / IN_WIDTH: ping_storage_data_697 <= (fillup_transition == 1'b1) ? i_input_data[240 % IN_WIDTH] : ping_storage_data_697 ^ i_input_data[240 % IN_WIDTH];
                599 / IN_WIDTH: ping_storage_data_697 <= (fillup_transition == 1'b1) ? i_input_data[599 % IN_WIDTH] : ping_storage_data_697 ^ i_input_data[599 % IN_WIDTH];
                938 / IN_WIDTH: ping_storage_data_697 <= (fillup_transition == 1'b1) ? i_input_data[938 % IN_WIDTH] : ping_storage_data_697 ^ i_input_data[938 % IN_WIDTH];
                default: ping_storage_data_697 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_697;
                endcase
            end else begin
                case (input_count)
                110 / IN_WIDTH: pong_storage_data_697 <= (fillup_transition == 1'b1) ? i_input_data[110 % IN_WIDTH] : pong_storage_data_697 ^ i_input_data[110 % IN_WIDTH];
                240 / IN_WIDTH: pong_storage_data_697 <= (fillup_transition == 1'b1) ? i_input_data[240 % IN_WIDTH] : pong_storage_data_697 ^ i_input_data[240 % IN_WIDTH];
                599 / IN_WIDTH: pong_storage_data_697 <= (fillup_transition == 1'b1) ? i_input_data[599 % IN_WIDTH] : pong_storage_data_697 ^ i_input_data[599 % IN_WIDTH];
                938 / IN_WIDTH: pong_storage_data_697 <= (fillup_transition == 1'b1) ? i_input_data[938 % IN_WIDTH] : pong_storage_data_697 ^ i_input_data[938 % IN_WIDTH];
                default: pong_storage_data_697 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_697;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_697 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_697;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_697 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_697;
            end
        end
    end
end

logic ping_storage_data_698;
logic pong_storage_data_698;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_698 <= 1'b0;
        pong_storage_data_698 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                111 / IN_WIDTH: ping_storage_data_698 <= (fillup_transition == 1'b1) ? i_input_data[111 % IN_WIDTH] : ping_storage_data_698 ^ i_input_data[111 % IN_WIDTH];
                241 / IN_WIDTH: ping_storage_data_698 <= (fillup_transition == 1'b1) ? i_input_data[241 % IN_WIDTH] : ping_storage_data_698 ^ i_input_data[241 % IN_WIDTH];
                600 / IN_WIDTH: ping_storage_data_698 <= (fillup_transition == 1'b1) ? i_input_data[600 % IN_WIDTH] : ping_storage_data_698 ^ i_input_data[600 % IN_WIDTH];
                939 / IN_WIDTH: ping_storage_data_698 <= (fillup_transition == 1'b1) ? i_input_data[939 % IN_WIDTH] : ping_storage_data_698 ^ i_input_data[939 % IN_WIDTH];
                default: ping_storage_data_698 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_698;
                endcase
            end else begin
                case (input_count)
                111 / IN_WIDTH: pong_storage_data_698 <= (fillup_transition == 1'b1) ? i_input_data[111 % IN_WIDTH] : pong_storage_data_698 ^ i_input_data[111 % IN_WIDTH];
                241 / IN_WIDTH: pong_storage_data_698 <= (fillup_transition == 1'b1) ? i_input_data[241 % IN_WIDTH] : pong_storage_data_698 ^ i_input_data[241 % IN_WIDTH];
                600 / IN_WIDTH: pong_storage_data_698 <= (fillup_transition == 1'b1) ? i_input_data[600 % IN_WIDTH] : pong_storage_data_698 ^ i_input_data[600 % IN_WIDTH];
                939 / IN_WIDTH: pong_storage_data_698 <= (fillup_transition == 1'b1) ? i_input_data[939 % IN_WIDTH] : pong_storage_data_698 ^ i_input_data[939 % IN_WIDTH];
                default: pong_storage_data_698 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_698;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_698 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_698;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_698 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_698;
            end
        end
    end
end

logic ping_storage_data_699;
logic pong_storage_data_699;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_699 <= 1'b0;
        pong_storage_data_699 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                112 / IN_WIDTH: ping_storage_data_699 <= (fillup_transition == 1'b1) ? i_input_data[112 % IN_WIDTH] : ping_storage_data_699 ^ i_input_data[112 % IN_WIDTH];
                242 / IN_WIDTH: ping_storage_data_699 <= (fillup_transition == 1'b1) ? i_input_data[242 % IN_WIDTH] : ping_storage_data_699 ^ i_input_data[242 % IN_WIDTH];
                601 / IN_WIDTH: ping_storage_data_699 <= (fillup_transition == 1'b1) ? i_input_data[601 % IN_WIDTH] : ping_storage_data_699 ^ i_input_data[601 % IN_WIDTH];
                940 / IN_WIDTH: ping_storage_data_699 <= (fillup_transition == 1'b1) ? i_input_data[940 % IN_WIDTH] : ping_storage_data_699 ^ i_input_data[940 % IN_WIDTH];
                default: ping_storage_data_699 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_699;
                endcase
            end else begin
                case (input_count)
                112 / IN_WIDTH: pong_storage_data_699 <= (fillup_transition == 1'b1) ? i_input_data[112 % IN_WIDTH] : pong_storage_data_699 ^ i_input_data[112 % IN_WIDTH];
                242 / IN_WIDTH: pong_storage_data_699 <= (fillup_transition == 1'b1) ? i_input_data[242 % IN_WIDTH] : pong_storage_data_699 ^ i_input_data[242 % IN_WIDTH];
                601 / IN_WIDTH: pong_storage_data_699 <= (fillup_transition == 1'b1) ? i_input_data[601 % IN_WIDTH] : pong_storage_data_699 ^ i_input_data[601 % IN_WIDTH];
                940 / IN_WIDTH: pong_storage_data_699 <= (fillup_transition == 1'b1) ? i_input_data[940 % IN_WIDTH] : pong_storage_data_699 ^ i_input_data[940 % IN_WIDTH];
                default: pong_storage_data_699 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_699;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_699 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_699;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_699 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_699;
            end
        end
    end
end

logic ping_storage_data_700;
logic pong_storage_data_700;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_700 <= 1'b0;
        pong_storage_data_700 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                113 / IN_WIDTH: ping_storage_data_700 <= (fillup_transition == 1'b1) ? i_input_data[113 % IN_WIDTH] : ping_storage_data_700 ^ i_input_data[113 % IN_WIDTH];
                243 / IN_WIDTH: ping_storage_data_700 <= (fillup_transition == 1'b1) ? i_input_data[243 % IN_WIDTH] : ping_storage_data_700 ^ i_input_data[243 % IN_WIDTH];
                602 / IN_WIDTH: ping_storage_data_700 <= (fillup_transition == 1'b1) ? i_input_data[602 % IN_WIDTH] : ping_storage_data_700 ^ i_input_data[602 % IN_WIDTH];
                941 / IN_WIDTH: ping_storage_data_700 <= (fillup_transition == 1'b1) ? i_input_data[941 % IN_WIDTH] : ping_storage_data_700 ^ i_input_data[941 % IN_WIDTH];
                default: ping_storage_data_700 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_700;
                endcase
            end else begin
                case (input_count)
                113 / IN_WIDTH: pong_storage_data_700 <= (fillup_transition == 1'b1) ? i_input_data[113 % IN_WIDTH] : pong_storage_data_700 ^ i_input_data[113 % IN_WIDTH];
                243 / IN_WIDTH: pong_storage_data_700 <= (fillup_transition == 1'b1) ? i_input_data[243 % IN_WIDTH] : pong_storage_data_700 ^ i_input_data[243 % IN_WIDTH];
                602 / IN_WIDTH: pong_storage_data_700 <= (fillup_transition == 1'b1) ? i_input_data[602 % IN_WIDTH] : pong_storage_data_700 ^ i_input_data[602 % IN_WIDTH];
                941 / IN_WIDTH: pong_storage_data_700 <= (fillup_transition == 1'b1) ? i_input_data[941 % IN_WIDTH] : pong_storage_data_700 ^ i_input_data[941 % IN_WIDTH];
                default: pong_storage_data_700 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_700;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_700 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_700;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_700 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_700;
            end
        end
    end
end

logic ping_storage_data_701;
logic pong_storage_data_701;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_701 <= 1'b0;
        pong_storage_data_701 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                114 / IN_WIDTH: ping_storage_data_701 <= (fillup_transition == 1'b1) ? i_input_data[114 % IN_WIDTH] : ping_storage_data_701 ^ i_input_data[114 % IN_WIDTH];
                244 / IN_WIDTH: ping_storage_data_701 <= (fillup_transition == 1'b1) ? i_input_data[244 % IN_WIDTH] : ping_storage_data_701 ^ i_input_data[244 % IN_WIDTH];
                603 / IN_WIDTH: ping_storage_data_701 <= (fillup_transition == 1'b1) ? i_input_data[603 % IN_WIDTH] : ping_storage_data_701 ^ i_input_data[603 % IN_WIDTH];
                942 / IN_WIDTH: ping_storage_data_701 <= (fillup_transition == 1'b1) ? i_input_data[942 % IN_WIDTH] : ping_storage_data_701 ^ i_input_data[942 % IN_WIDTH];
                default: ping_storage_data_701 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_701;
                endcase
            end else begin
                case (input_count)
                114 / IN_WIDTH: pong_storage_data_701 <= (fillup_transition == 1'b1) ? i_input_data[114 % IN_WIDTH] : pong_storage_data_701 ^ i_input_data[114 % IN_WIDTH];
                244 / IN_WIDTH: pong_storage_data_701 <= (fillup_transition == 1'b1) ? i_input_data[244 % IN_WIDTH] : pong_storage_data_701 ^ i_input_data[244 % IN_WIDTH];
                603 / IN_WIDTH: pong_storage_data_701 <= (fillup_transition == 1'b1) ? i_input_data[603 % IN_WIDTH] : pong_storage_data_701 ^ i_input_data[603 % IN_WIDTH];
                942 / IN_WIDTH: pong_storage_data_701 <= (fillup_transition == 1'b1) ? i_input_data[942 % IN_WIDTH] : pong_storage_data_701 ^ i_input_data[942 % IN_WIDTH];
                default: pong_storage_data_701 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_701;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_701 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_701;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_701 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_701;
            end
        end
    end
end

logic ping_storage_data_702;
logic pong_storage_data_702;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_702 <= 1'b0;
        pong_storage_data_702 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                115 / IN_WIDTH: ping_storage_data_702 <= (fillup_transition == 1'b1) ? i_input_data[115 % IN_WIDTH] : ping_storage_data_702 ^ i_input_data[115 % IN_WIDTH];
                245 / IN_WIDTH: ping_storage_data_702 <= (fillup_transition == 1'b1) ? i_input_data[245 % IN_WIDTH] : ping_storage_data_702 ^ i_input_data[245 % IN_WIDTH];
                604 / IN_WIDTH: ping_storage_data_702 <= (fillup_transition == 1'b1) ? i_input_data[604 % IN_WIDTH] : ping_storage_data_702 ^ i_input_data[604 % IN_WIDTH];
                943 / IN_WIDTH: ping_storage_data_702 <= (fillup_transition == 1'b1) ? i_input_data[943 % IN_WIDTH] : ping_storage_data_702 ^ i_input_data[943 % IN_WIDTH];
                default: ping_storage_data_702 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_702;
                endcase
            end else begin
                case (input_count)
                115 / IN_WIDTH: pong_storage_data_702 <= (fillup_transition == 1'b1) ? i_input_data[115 % IN_WIDTH] : pong_storage_data_702 ^ i_input_data[115 % IN_WIDTH];
                245 / IN_WIDTH: pong_storage_data_702 <= (fillup_transition == 1'b1) ? i_input_data[245 % IN_WIDTH] : pong_storage_data_702 ^ i_input_data[245 % IN_WIDTH];
                604 / IN_WIDTH: pong_storage_data_702 <= (fillup_transition == 1'b1) ? i_input_data[604 % IN_WIDTH] : pong_storage_data_702 ^ i_input_data[604 % IN_WIDTH];
                943 / IN_WIDTH: pong_storage_data_702 <= (fillup_transition == 1'b1) ? i_input_data[943 % IN_WIDTH] : pong_storage_data_702 ^ i_input_data[943 % IN_WIDTH];
                default: pong_storage_data_702 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_702;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_702 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_702;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_702 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_702;
            end
        end
    end
end

logic ping_storage_data_703;
logic pong_storage_data_703;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_703 <= 1'b0;
        pong_storage_data_703 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                116 / IN_WIDTH: ping_storage_data_703 <= (fillup_transition == 1'b1) ? i_input_data[116 % IN_WIDTH] : ping_storage_data_703 ^ i_input_data[116 % IN_WIDTH];
                246 / IN_WIDTH: ping_storage_data_703 <= (fillup_transition == 1'b1) ? i_input_data[246 % IN_WIDTH] : ping_storage_data_703 ^ i_input_data[246 % IN_WIDTH];
                605 / IN_WIDTH: ping_storage_data_703 <= (fillup_transition == 1'b1) ? i_input_data[605 % IN_WIDTH] : ping_storage_data_703 ^ i_input_data[605 % IN_WIDTH];
                944 / IN_WIDTH: ping_storage_data_703 <= (fillup_transition == 1'b1) ? i_input_data[944 % IN_WIDTH] : ping_storage_data_703 ^ i_input_data[944 % IN_WIDTH];
                default: ping_storage_data_703 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_703;
                endcase
            end else begin
                case (input_count)
                116 / IN_WIDTH: pong_storage_data_703 <= (fillup_transition == 1'b1) ? i_input_data[116 % IN_WIDTH] : pong_storage_data_703 ^ i_input_data[116 % IN_WIDTH];
                246 / IN_WIDTH: pong_storage_data_703 <= (fillup_transition == 1'b1) ? i_input_data[246 % IN_WIDTH] : pong_storage_data_703 ^ i_input_data[246 % IN_WIDTH];
                605 / IN_WIDTH: pong_storage_data_703 <= (fillup_transition == 1'b1) ? i_input_data[605 % IN_WIDTH] : pong_storage_data_703 ^ i_input_data[605 % IN_WIDTH];
                944 / IN_WIDTH: pong_storage_data_703 <= (fillup_transition == 1'b1) ? i_input_data[944 % IN_WIDTH] : pong_storage_data_703 ^ i_input_data[944 % IN_WIDTH];
                default: pong_storage_data_703 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_703;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_703 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_703;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_703 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_703;
            end
        end
    end
end

logic ping_storage_data_704;
logic pong_storage_data_704;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_704 <= 1'b0;
        pong_storage_data_704 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                117 / IN_WIDTH: ping_storage_data_704 <= (fillup_transition == 1'b1) ? i_input_data[117 % IN_WIDTH] : ping_storage_data_704 ^ i_input_data[117 % IN_WIDTH];
                247 / IN_WIDTH: ping_storage_data_704 <= (fillup_transition == 1'b1) ? i_input_data[247 % IN_WIDTH] : ping_storage_data_704 ^ i_input_data[247 % IN_WIDTH];
                606 / IN_WIDTH: ping_storage_data_704 <= (fillup_transition == 1'b1) ? i_input_data[606 % IN_WIDTH] : ping_storage_data_704 ^ i_input_data[606 % IN_WIDTH];
                945 / IN_WIDTH: ping_storage_data_704 <= (fillup_transition == 1'b1) ? i_input_data[945 % IN_WIDTH] : ping_storage_data_704 ^ i_input_data[945 % IN_WIDTH];
                default: ping_storage_data_704 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_704;
                endcase
            end else begin
                case (input_count)
                117 / IN_WIDTH: pong_storage_data_704 <= (fillup_transition == 1'b1) ? i_input_data[117 % IN_WIDTH] : pong_storage_data_704 ^ i_input_data[117 % IN_WIDTH];
                247 / IN_WIDTH: pong_storage_data_704 <= (fillup_transition == 1'b1) ? i_input_data[247 % IN_WIDTH] : pong_storage_data_704 ^ i_input_data[247 % IN_WIDTH];
                606 / IN_WIDTH: pong_storage_data_704 <= (fillup_transition == 1'b1) ? i_input_data[606 % IN_WIDTH] : pong_storage_data_704 ^ i_input_data[606 % IN_WIDTH];
                945 / IN_WIDTH: pong_storage_data_704 <= (fillup_transition == 1'b1) ? i_input_data[945 % IN_WIDTH] : pong_storage_data_704 ^ i_input_data[945 % IN_WIDTH];
                default: pong_storage_data_704 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_704;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_704 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_704;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_704 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_704;
            end
        end
    end
end

logic ping_storage_data_705;
logic pong_storage_data_705;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_705 <= 1'b0;
        pong_storage_data_705 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                118 / IN_WIDTH: ping_storage_data_705 <= (fillup_transition == 1'b1) ? i_input_data[118 % IN_WIDTH] : ping_storage_data_705 ^ i_input_data[118 % IN_WIDTH];
                248 / IN_WIDTH: ping_storage_data_705 <= (fillup_transition == 1'b1) ? i_input_data[248 % IN_WIDTH] : ping_storage_data_705 ^ i_input_data[248 % IN_WIDTH];
                607 / IN_WIDTH: ping_storage_data_705 <= (fillup_transition == 1'b1) ? i_input_data[607 % IN_WIDTH] : ping_storage_data_705 ^ i_input_data[607 % IN_WIDTH];
                946 / IN_WIDTH: ping_storage_data_705 <= (fillup_transition == 1'b1) ? i_input_data[946 % IN_WIDTH] : ping_storage_data_705 ^ i_input_data[946 % IN_WIDTH];
                default: ping_storage_data_705 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_705;
                endcase
            end else begin
                case (input_count)
                118 / IN_WIDTH: pong_storage_data_705 <= (fillup_transition == 1'b1) ? i_input_data[118 % IN_WIDTH] : pong_storage_data_705 ^ i_input_data[118 % IN_WIDTH];
                248 / IN_WIDTH: pong_storage_data_705 <= (fillup_transition == 1'b1) ? i_input_data[248 % IN_WIDTH] : pong_storage_data_705 ^ i_input_data[248 % IN_WIDTH];
                607 / IN_WIDTH: pong_storage_data_705 <= (fillup_transition == 1'b1) ? i_input_data[607 % IN_WIDTH] : pong_storage_data_705 ^ i_input_data[607 % IN_WIDTH];
                946 / IN_WIDTH: pong_storage_data_705 <= (fillup_transition == 1'b1) ? i_input_data[946 % IN_WIDTH] : pong_storage_data_705 ^ i_input_data[946 % IN_WIDTH];
                default: pong_storage_data_705 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_705;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_705 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_705;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_705 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_705;
            end
        end
    end
end

logic ping_storage_data_706;
logic pong_storage_data_706;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_706 <= 1'b0;
        pong_storage_data_706 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                119 / IN_WIDTH: ping_storage_data_706 <= (fillup_transition == 1'b1) ? i_input_data[119 % IN_WIDTH] : ping_storage_data_706 ^ i_input_data[119 % IN_WIDTH];
                249 / IN_WIDTH: ping_storage_data_706 <= (fillup_transition == 1'b1) ? i_input_data[249 % IN_WIDTH] : ping_storage_data_706 ^ i_input_data[249 % IN_WIDTH];
                608 / IN_WIDTH: ping_storage_data_706 <= (fillup_transition == 1'b1) ? i_input_data[608 % IN_WIDTH] : ping_storage_data_706 ^ i_input_data[608 % IN_WIDTH];
                947 / IN_WIDTH: ping_storage_data_706 <= (fillup_transition == 1'b1) ? i_input_data[947 % IN_WIDTH] : ping_storage_data_706 ^ i_input_data[947 % IN_WIDTH];
                default: ping_storage_data_706 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_706;
                endcase
            end else begin
                case (input_count)
                119 / IN_WIDTH: pong_storage_data_706 <= (fillup_transition == 1'b1) ? i_input_data[119 % IN_WIDTH] : pong_storage_data_706 ^ i_input_data[119 % IN_WIDTH];
                249 / IN_WIDTH: pong_storage_data_706 <= (fillup_transition == 1'b1) ? i_input_data[249 % IN_WIDTH] : pong_storage_data_706 ^ i_input_data[249 % IN_WIDTH];
                608 / IN_WIDTH: pong_storage_data_706 <= (fillup_transition == 1'b1) ? i_input_data[608 % IN_WIDTH] : pong_storage_data_706 ^ i_input_data[608 % IN_WIDTH];
                947 / IN_WIDTH: pong_storage_data_706 <= (fillup_transition == 1'b1) ? i_input_data[947 % IN_WIDTH] : pong_storage_data_706 ^ i_input_data[947 % IN_WIDTH];
                default: pong_storage_data_706 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_706;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_706 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_706;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_706 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_706;
            end
        end
    end
end

logic ping_storage_data_707;
logic pong_storage_data_707;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_707 <= 1'b0;
        pong_storage_data_707 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                120 / IN_WIDTH: ping_storage_data_707 <= (fillup_transition == 1'b1) ? i_input_data[120 % IN_WIDTH] : ping_storage_data_707 ^ i_input_data[120 % IN_WIDTH];
                250 / IN_WIDTH: ping_storage_data_707 <= (fillup_transition == 1'b1) ? i_input_data[250 % IN_WIDTH] : ping_storage_data_707 ^ i_input_data[250 % IN_WIDTH];
                609 / IN_WIDTH: ping_storage_data_707 <= (fillup_transition == 1'b1) ? i_input_data[609 % IN_WIDTH] : ping_storage_data_707 ^ i_input_data[609 % IN_WIDTH];
                948 / IN_WIDTH: ping_storage_data_707 <= (fillup_transition == 1'b1) ? i_input_data[948 % IN_WIDTH] : ping_storage_data_707 ^ i_input_data[948 % IN_WIDTH];
                default: ping_storage_data_707 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_707;
                endcase
            end else begin
                case (input_count)
                120 / IN_WIDTH: pong_storage_data_707 <= (fillup_transition == 1'b1) ? i_input_data[120 % IN_WIDTH] : pong_storage_data_707 ^ i_input_data[120 % IN_WIDTH];
                250 / IN_WIDTH: pong_storage_data_707 <= (fillup_transition == 1'b1) ? i_input_data[250 % IN_WIDTH] : pong_storage_data_707 ^ i_input_data[250 % IN_WIDTH];
                609 / IN_WIDTH: pong_storage_data_707 <= (fillup_transition == 1'b1) ? i_input_data[609 % IN_WIDTH] : pong_storage_data_707 ^ i_input_data[609 % IN_WIDTH];
                948 / IN_WIDTH: pong_storage_data_707 <= (fillup_transition == 1'b1) ? i_input_data[948 % IN_WIDTH] : pong_storage_data_707 ^ i_input_data[948 % IN_WIDTH];
                default: pong_storage_data_707 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_707;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_707 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_707;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_707 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_707;
            end
        end
    end
end

logic ping_storage_data_708;
logic pong_storage_data_708;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_708 <= 1'b0;
        pong_storage_data_708 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                121 / IN_WIDTH: ping_storage_data_708 <= (fillup_transition == 1'b1) ? i_input_data[121 % IN_WIDTH] : ping_storage_data_708 ^ i_input_data[121 % IN_WIDTH];
                251 / IN_WIDTH: ping_storage_data_708 <= (fillup_transition == 1'b1) ? i_input_data[251 % IN_WIDTH] : ping_storage_data_708 ^ i_input_data[251 % IN_WIDTH];
                610 / IN_WIDTH: ping_storage_data_708 <= (fillup_transition == 1'b1) ? i_input_data[610 % IN_WIDTH] : ping_storage_data_708 ^ i_input_data[610 % IN_WIDTH];
                949 / IN_WIDTH: ping_storage_data_708 <= (fillup_transition == 1'b1) ? i_input_data[949 % IN_WIDTH] : ping_storage_data_708 ^ i_input_data[949 % IN_WIDTH];
                default: ping_storage_data_708 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_708;
                endcase
            end else begin
                case (input_count)
                121 / IN_WIDTH: pong_storage_data_708 <= (fillup_transition == 1'b1) ? i_input_data[121 % IN_WIDTH] : pong_storage_data_708 ^ i_input_data[121 % IN_WIDTH];
                251 / IN_WIDTH: pong_storage_data_708 <= (fillup_transition == 1'b1) ? i_input_data[251 % IN_WIDTH] : pong_storage_data_708 ^ i_input_data[251 % IN_WIDTH];
                610 / IN_WIDTH: pong_storage_data_708 <= (fillup_transition == 1'b1) ? i_input_data[610 % IN_WIDTH] : pong_storage_data_708 ^ i_input_data[610 % IN_WIDTH];
                949 / IN_WIDTH: pong_storage_data_708 <= (fillup_transition == 1'b1) ? i_input_data[949 % IN_WIDTH] : pong_storage_data_708 ^ i_input_data[949 % IN_WIDTH];
                default: pong_storage_data_708 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_708;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_708 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_708;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_708 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_708;
            end
        end
    end
end

logic ping_storage_data_709;
logic pong_storage_data_709;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_709 <= 1'b0;
        pong_storage_data_709 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                122 / IN_WIDTH: ping_storage_data_709 <= (fillup_transition == 1'b1) ? i_input_data[122 % IN_WIDTH] : ping_storage_data_709 ^ i_input_data[122 % IN_WIDTH];
                252 / IN_WIDTH: ping_storage_data_709 <= (fillup_transition == 1'b1) ? i_input_data[252 % IN_WIDTH] : ping_storage_data_709 ^ i_input_data[252 % IN_WIDTH];
                611 / IN_WIDTH: ping_storage_data_709 <= (fillup_transition == 1'b1) ? i_input_data[611 % IN_WIDTH] : ping_storage_data_709 ^ i_input_data[611 % IN_WIDTH];
                950 / IN_WIDTH: ping_storage_data_709 <= (fillup_transition == 1'b1) ? i_input_data[950 % IN_WIDTH] : ping_storage_data_709 ^ i_input_data[950 % IN_WIDTH];
                default: ping_storage_data_709 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_709;
                endcase
            end else begin
                case (input_count)
                122 / IN_WIDTH: pong_storage_data_709 <= (fillup_transition == 1'b1) ? i_input_data[122 % IN_WIDTH] : pong_storage_data_709 ^ i_input_data[122 % IN_WIDTH];
                252 / IN_WIDTH: pong_storage_data_709 <= (fillup_transition == 1'b1) ? i_input_data[252 % IN_WIDTH] : pong_storage_data_709 ^ i_input_data[252 % IN_WIDTH];
                611 / IN_WIDTH: pong_storage_data_709 <= (fillup_transition == 1'b1) ? i_input_data[611 % IN_WIDTH] : pong_storage_data_709 ^ i_input_data[611 % IN_WIDTH];
                950 / IN_WIDTH: pong_storage_data_709 <= (fillup_transition == 1'b1) ? i_input_data[950 % IN_WIDTH] : pong_storage_data_709 ^ i_input_data[950 % IN_WIDTH];
                default: pong_storage_data_709 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_709;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_709 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_709;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_709 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_709;
            end
        end
    end
end

logic ping_storage_data_710;
logic pong_storage_data_710;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_710 <= 1'b0;
        pong_storage_data_710 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                123 / IN_WIDTH: ping_storage_data_710 <= (fillup_transition == 1'b1) ? i_input_data[123 % IN_WIDTH] : ping_storage_data_710 ^ i_input_data[123 % IN_WIDTH];
                253 / IN_WIDTH: ping_storage_data_710 <= (fillup_transition == 1'b1) ? i_input_data[253 % IN_WIDTH] : ping_storage_data_710 ^ i_input_data[253 % IN_WIDTH];
                612 / IN_WIDTH: ping_storage_data_710 <= (fillup_transition == 1'b1) ? i_input_data[612 % IN_WIDTH] : ping_storage_data_710 ^ i_input_data[612 % IN_WIDTH];
                951 / IN_WIDTH: ping_storage_data_710 <= (fillup_transition == 1'b1) ? i_input_data[951 % IN_WIDTH] : ping_storage_data_710 ^ i_input_data[951 % IN_WIDTH];
                default: ping_storage_data_710 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_710;
                endcase
            end else begin
                case (input_count)
                123 / IN_WIDTH: pong_storage_data_710 <= (fillup_transition == 1'b1) ? i_input_data[123 % IN_WIDTH] : pong_storage_data_710 ^ i_input_data[123 % IN_WIDTH];
                253 / IN_WIDTH: pong_storage_data_710 <= (fillup_transition == 1'b1) ? i_input_data[253 % IN_WIDTH] : pong_storage_data_710 ^ i_input_data[253 % IN_WIDTH];
                612 / IN_WIDTH: pong_storage_data_710 <= (fillup_transition == 1'b1) ? i_input_data[612 % IN_WIDTH] : pong_storage_data_710 ^ i_input_data[612 % IN_WIDTH];
                951 / IN_WIDTH: pong_storage_data_710 <= (fillup_transition == 1'b1) ? i_input_data[951 % IN_WIDTH] : pong_storage_data_710 ^ i_input_data[951 % IN_WIDTH];
                default: pong_storage_data_710 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_710;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_710 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_710;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_710 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_710;
            end
        end
    end
end

logic ping_storage_data_711;
logic pong_storage_data_711;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_711 <= 1'b0;
        pong_storage_data_711 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                124 / IN_WIDTH: ping_storage_data_711 <= (fillup_transition == 1'b1) ? i_input_data[124 % IN_WIDTH] : ping_storage_data_711 ^ i_input_data[124 % IN_WIDTH];
                254 / IN_WIDTH: ping_storage_data_711 <= (fillup_transition == 1'b1) ? i_input_data[254 % IN_WIDTH] : ping_storage_data_711 ^ i_input_data[254 % IN_WIDTH];
                613 / IN_WIDTH: ping_storage_data_711 <= (fillup_transition == 1'b1) ? i_input_data[613 % IN_WIDTH] : ping_storage_data_711 ^ i_input_data[613 % IN_WIDTH];
                952 / IN_WIDTH: ping_storage_data_711 <= (fillup_transition == 1'b1) ? i_input_data[952 % IN_WIDTH] : ping_storage_data_711 ^ i_input_data[952 % IN_WIDTH];
                default: ping_storage_data_711 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_711;
                endcase
            end else begin
                case (input_count)
                124 / IN_WIDTH: pong_storage_data_711 <= (fillup_transition == 1'b1) ? i_input_data[124 % IN_WIDTH] : pong_storage_data_711 ^ i_input_data[124 % IN_WIDTH];
                254 / IN_WIDTH: pong_storage_data_711 <= (fillup_transition == 1'b1) ? i_input_data[254 % IN_WIDTH] : pong_storage_data_711 ^ i_input_data[254 % IN_WIDTH];
                613 / IN_WIDTH: pong_storage_data_711 <= (fillup_transition == 1'b1) ? i_input_data[613 % IN_WIDTH] : pong_storage_data_711 ^ i_input_data[613 % IN_WIDTH];
                952 / IN_WIDTH: pong_storage_data_711 <= (fillup_transition == 1'b1) ? i_input_data[952 % IN_WIDTH] : pong_storage_data_711 ^ i_input_data[952 % IN_WIDTH];
                default: pong_storage_data_711 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_711;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_711 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_711;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_711 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_711;
            end
        end
    end
end

logic ping_storage_data_712;
logic pong_storage_data_712;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_712 <= 1'b0;
        pong_storage_data_712 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                125 / IN_WIDTH: ping_storage_data_712 <= (fillup_transition == 1'b1) ? i_input_data[125 % IN_WIDTH] : ping_storage_data_712 ^ i_input_data[125 % IN_WIDTH];
                255 / IN_WIDTH: ping_storage_data_712 <= (fillup_transition == 1'b1) ? i_input_data[255 % IN_WIDTH] : ping_storage_data_712 ^ i_input_data[255 % IN_WIDTH];
                614 / IN_WIDTH: ping_storage_data_712 <= (fillup_transition == 1'b1) ? i_input_data[614 % IN_WIDTH] : ping_storage_data_712 ^ i_input_data[614 % IN_WIDTH];
                953 / IN_WIDTH: ping_storage_data_712 <= (fillup_transition == 1'b1) ? i_input_data[953 % IN_WIDTH] : ping_storage_data_712 ^ i_input_data[953 % IN_WIDTH];
                default: ping_storage_data_712 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_712;
                endcase
            end else begin
                case (input_count)
                125 / IN_WIDTH: pong_storage_data_712 <= (fillup_transition == 1'b1) ? i_input_data[125 % IN_WIDTH] : pong_storage_data_712 ^ i_input_data[125 % IN_WIDTH];
                255 / IN_WIDTH: pong_storage_data_712 <= (fillup_transition == 1'b1) ? i_input_data[255 % IN_WIDTH] : pong_storage_data_712 ^ i_input_data[255 % IN_WIDTH];
                614 / IN_WIDTH: pong_storage_data_712 <= (fillup_transition == 1'b1) ? i_input_data[614 % IN_WIDTH] : pong_storage_data_712 ^ i_input_data[614 % IN_WIDTH];
                953 / IN_WIDTH: pong_storage_data_712 <= (fillup_transition == 1'b1) ? i_input_data[953 % IN_WIDTH] : pong_storage_data_712 ^ i_input_data[953 % IN_WIDTH];
                default: pong_storage_data_712 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_712;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_712 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_712;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_712 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_712;
            end
        end
    end
end

logic ping_storage_data_713;
logic pong_storage_data_713;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_713 <= 1'b0;
        pong_storage_data_713 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                126 / IN_WIDTH: ping_storage_data_713 <= (fillup_transition == 1'b1) ? i_input_data[126 % IN_WIDTH] : ping_storage_data_713 ^ i_input_data[126 % IN_WIDTH];
                256 / IN_WIDTH: ping_storage_data_713 <= (fillup_transition == 1'b1) ? i_input_data[256 % IN_WIDTH] : ping_storage_data_713 ^ i_input_data[256 % IN_WIDTH];
                615 / IN_WIDTH: ping_storage_data_713 <= (fillup_transition == 1'b1) ? i_input_data[615 % IN_WIDTH] : ping_storage_data_713 ^ i_input_data[615 % IN_WIDTH];
                954 / IN_WIDTH: ping_storage_data_713 <= (fillup_transition == 1'b1) ? i_input_data[954 % IN_WIDTH] : ping_storage_data_713 ^ i_input_data[954 % IN_WIDTH];
                default: ping_storage_data_713 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_713;
                endcase
            end else begin
                case (input_count)
                126 / IN_WIDTH: pong_storage_data_713 <= (fillup_transition == 1'b1) ? i_input_data[126 % IN_WIDTH] : pong_storage_data_713 ^ i_input_data[126 % IN_WIDTH];
                256 / IN_WIDTH: pong_storage_data_713 <= (fillup_transition == 1'b1) ? i_input_data[256 % IN_WIDTH] : pong_storage_data_713 ^ i_input_data[256 % IN_WIDTH];
                615 / IN_WIDTH: pong_storage_data_713 <= (fillup_transition == 1'b1) ? i_input_data[615 % IN_WIDTH] : pong_storage_data_713 ^ i_input_data[615 % IN_WIDTH];
                954 / IN_WIDTH: pong_storage_data_713 <= (fillup_transition == 1'b1) ? i_input_data[954 % IN_WIDTH] : pong_storage_data_713 ^ i_input_data[954 % IN_WIDTH];
                default: pong_storage_data_713 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_713;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_713 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_713;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_713 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_713;
            end
        end
    end
end

logic ping_storage_data_714;
logic pong_storage_data_714;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_714 <= 1'b0;
        pong_storage_data_714 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                127 / IN_WIDTH: ping_storage_data_714 <= (fillup_transition == 1'b1) ? i_input_data[127 % IN_WIDTH] : ping_storage_data_714 ^ i_input_data[127 % IN_WIDTH];
                257 / IN_WIDTH: ping_storage_data_714 <= (fillup_transition == 1'b1) ? i_input_data[257 % IN_WIDTH] : ping_storage_data_714 ^ i_input_data[257 % IN_WIDTH];
                616 / IN_WIDTH: ping_storage_data_714 <= (fillup_transition == 1'b1) ? i_input_data[616 % IN_WIDTH] : ping_storage_data_714 ^ i_input_data[616 % IN_WIDTH];
                955 / IN_WIDTH: ping_storage_data_714 <= (fillup_transition == 1'b1) ? i_input_data[955 % IN_WIDTH] : ping_storage_data_714 ^ i_input_data[955 % IN_WIDTH];
                default: ping_storage_data_714 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_714;
                endcase
            end else begin
                case (input_count)
                127 / IN_WIDTH: pong_storage_data_714 <= (fillup_transition == 1'b1) ? i_input_data[127 % IN_WIDTH] : pong_storage_data_714 ^ i_input_data[127 % IN_WIDTH];
                257 / IN_WIDTH: pong_storage_data_714 <= (fillup_transition == 1'b1) ? i_input_data[257 % IN_WIDTH] : pong_storage_data_714 ^ i_input_data[257 % IN_WIDTH];
                616 / IN_WIDTH: pong_storage_data_714 <= (fillup_transition == 1'b1) ? i_input_data[616 % IN_WIDTH] : pong_storage_data_714 ^ i_input_data[616 % IN_WIDTH];
                955 / IN_WIDTH: pong_storage_data_714 <= (fillup_transition == 1'b1) ? i_input_data[955 % IN_WIDTH] : pong_storage_data_714 ^ i_input_data[955 % IN_WIDTH];
                default: pong_storage_data_714 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_714;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_714 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_714;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_714 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_714;
            end
        end
    end
end

logic ping_storage_data_715;
logic pong_storage_data_715;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_715 <= 1'b0;
        pong_storage_data_715 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                128 / IN_WIDTH: ping_storage_data_715 <= (fillup_transition == 1'b1) ? i_input_data[128 % IN_WIDTH] : ping_storage_data_715 ^ i_input_data[128 % IN_WIDTH];
                258 / IN_WIDTH: ping_storage_data_715 <= (fillup_transition == 1'b1) ? i_input_data[258 % IN_WIDTH] : ping_storage_data_715 ^ i_input_data[258 % IN_WIDTH];
                617 / IN_WIDTH: ping_storage_data_715 <= (fillup_transition == 1'b1) ? i_input_data[617 % IN_WIDTH] : ping_storage_data_715 ^ i_input_data[617 % IN_WIDTH];
                956 / IN_WIDTH: ping_storage_data_715 <= (fillup_transition == 1'b1) ? i_input_data[956 % IN_WIDTH] : ping_storage_data_715 ^ i_input_data[956 % IN_WIDTH];
                default: ping_storage_data_715 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_715;
                endcase
            end else begin
                case (input_count)
                128 / IN_WIDTH: pong_storage_data_715 <= (fillup_transition == 1'b1) ? i_input_data[128 % IN_WIDTH] : pong_storage_data_715 ^ i_input_data[128 % IN_WIDTH];
                258 / IN_WIDTH: pong_storage_data_715 <= (fillup_transition == 1'b1) ? i_input_data[258 % IN_WIDTH] : pong_storage_data_715 ^ i_input_data[258 % IN_WIDTH];
                617 / IN_WIDTH: pong_storage_data_715 <= (fillup_transition == 1'b1) ? i_input_data[617 % IN_WIDTH] : pong_storage_data_715 ^ i_input_data[617 % IN_WIDTH];
                956 / IN_WIDTH: pong_storage_data_715 <= (fillup_transition == 1'b1) ? i_input_data[956 % IN_WIDTH] : pong_storage_data_715 ^ i_input_data[956 % IN_WIDTH];
                default: pong_storage_data_715 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_715;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_715 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_715;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_715 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_715;
            end
        end
    end
end

logic ping_storage_data_716;
logic pong_storage_data_716;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_716 <= 1'b0;
        pong_storage_data_716 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                129 / IN_WIDTH: ping_storage_data_716 <= (fillup_transition == 1'b1) ? i_input_data[129 % IN_WIDTH] : ping_storage_data_716 ^ i_input_data[129 % IN_WIDTH];
                259 / IN_WIDTH: ping_storage_data_716 <= (fillup_transition == 1'b1) ? i_input_data[259 % IN_WIDTH] : ping_storage_data_716 ^ i_input_data[259 % IN_WIDTH];
                618 / IN_WIDTH: ping_storage_data_716 <= (fillup_transition == 1'b1) ? i_input_data[618 % IN_WIDTH] : ping_storage_data_716 ^ i_input_data[618 % IN_WIDTH];
                957 / IN_WIDTH: ping_storage_data_716 <= (fillup_transition == 1'b1) ? i_input_data[957 % IN_WIDTH] : ping_storage_data_716 ^ i_input_data[957 % IN_WIDTH];
                default: ping_storage_data_716 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_716;
                endcase
            end else begin
                case (input_count)
                129 / IN_WIDTH: pong_storage_data_716 <= (fillup_transition == 1'b1) ? i_input_data[129 % IN_WIDTH] : pong_storage_data_716 ^ i_input_data[129 % IN_WIDTH];
                259 / IN_WIDTH: pong_storage_data_716 <= (fillup_transition == 1'b1) ? i_input_data[259 % IN_WIDTH] : pong_storage_data_716 ^ i_input_data[259 % IN_WIDTH];
                618 / IN_WIDTH: pong_storage_data_716 <= (fillup_transition == 1'b1) ? i_input_data[618 % IN_WIDTH] : pong_storage_data_716 ^ i_input_data[618 % IN_WIDTH];
                957 / IN_WIDTH: pong_storage_data_716 <= (fillup_transition == 1'b1) ? i_input_data[957 % IN_WIDTH] : pong_storage_data_716 ^ i_input_data[957 % IN_WIDTH];
                default: pong_storage_data_716 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_716;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_716 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_716;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_716 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_716;
            end
        end
    end
end

logic ping_storage_data_717;
logic pong_storage_data_717;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_717 <= 1'b0;
        pong_storage_data_717 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                130 / IN_WIDTH: ping_storage_data_717 <= (fillup_transition == 1'b1) ? i_input_data[130 % IN_WIDTH] : ping_storage_data_717 ^ i_input_data[130 % IN_WIDTH];
                260 / IN_WIDTH: ping_storage_data_717 <= (fillup_transition == 1'b1) ? i_input_data[260 % IN_WIDTH] : ping_storage_data_717 ^ i_input_data[260 % IN_WIDTH];
                619 / IN_WIDTH: ping_storage_data_717 <= (fillup_transition == 1'b1) ? i_input_data[619 % IN_WIDTH] : ping_storage_data_717 ^ i_input_data[619 % IN_WIDTH];
                958 / IN_WIDTH: ping_storage_data_717 <= (fillup_transition == 1'b1) ? i_input_data[958 % IN_WIDTH] : ping_storage_data_717 ^ i_input_data[958 % IN_WIDTH];
                default: ping_storage_data_717 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_717;
                endcase
            end else begin
                case (input_count)
                130 / IN_WIDTH: pong_storage_data_717 <= (fillup_transition == 1'b1) ? i_input_data[130 % IN_WIDTH] : pong_storage_data_717 ^ i_input_data[130 % IN_WIDTH];
                260 / IN_WIDTH: pong_storage_data_717 <= (fillup_transition == 1'b1) ? i_input_data[260 % IN_WIDTH] : pong_storage_data_717 ^ i_input_data[260 % IN_WIDTH];
                619 / IN_WIDTH: pong_storage_data_717 <= (fillup_transition == 1'b1) ? i_input_data[619 % IN_WIDTH] : pong_storage_data_717 ^ i_input_data[619 % IN_WIDTH];
                958 / IN_WIDTH: pong_storage_data_717 <= (fillup_transition == 1'b1) ? i_input_data[958 % IN_WIDTH] : pong_storage_data_717 ^ i_input_data[958 % IN_WIDTH];
                default: pong_storage_data_717 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_717;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_717 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_717;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_717 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_717;
            end
        end
    end
end

logic ping_storage_data_718;
logic pong_storage_data_718;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_718 <= 1'b0;
        pong_storage_data_718 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                131 / IN_WIDTH: ping_storage_data_718 <= (fillup_transition == 1'b1) ? i_input_data[131 % IN_WIDTH] : ping_storage_data_718 ^ i_input_data[131 % IN_WIDTH];
                261 / IN_WIDTH: ping_storage_data_718 <= (fillup_transition == 1'b1) ? i_input_data[261 % IN_WIDTH] : ping_storage_data_718 ^ i_input_data[261 % IN_WIDTH];
                620 / IN_WIDTH: ping_storage_data_718 <= (fillup_transition == 1'b1) ? i_input_data[620 % IN_WIDTH] : ping_storage_data_718 ^ i_input_data[620 % IN_WIDTH];
                959 / IN_WIDTH: ping_storage_data_718 <= (fillup_transition == 1'b1) ? i_input_data[959 % IN_WIDTH] : ping_storage_data_718 ^ i_input_data[959 % IN_WIDTH];
                default: ping_storage_data_718 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_718;
                endcase
            end else begin
                case (input_count)
                131 / IN_WIDTH: pong_storage_data_718 <= (fillup_transition == 1'b1) ? i_input_data[131 % IN_WIDTH] : pong_storage_data_718 ^ i_input_data[131 % IN_WIDTH];
                261 / IN_WIDTH: pong_storage_data_718 <= (fillup_transition == 1'b1) ? i_input_data[261 % IN_WIDTH] : pong_storage_data_718 ^ i_input_data[261 % IN_WIDTH];
                620 / IN_WIDTH: pong_storage_data_718 <= (fillup_transition == 1'b1) ? i_input_data[620 % IN_WIDTH] : pong_storage_data_718 ^ i_input_data[620 % IN_WIDTH];
                959 / IN_WIDTH: pong_storage_data_718 <= (fillup_transition == 1'b1) ? i_input_data[959 % IN_WIDTH] : pong_storage_data_718 ^ i_input_data[959 % IN_WIDTH];
                default: pong_storage_data_718 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_718;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_718 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_718;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_718 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_718;
            end
        end
    end
end

logic ping_storage_data_719;
logic pong_storage_data_719;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_719 <= 1'b0;
        pong_storage_data_719 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                132 / IN_WIDTH: ping_storage_data_719 <= (fillup_transition == 1'b1) ? i_input_data[132 % IN_WIDTH] : ping_storage_data_719 ^ i_input_data[132 % IN_WIDTH];
                262 / IN_WIDTH: ping_storage_data_719 <= (fillup_transition == 1'b1) ? i_input_data[262 % IN_WIDTH] : ping_storage_data_719 ^ i_input_data[262 % IN_WIDTH];
                621 / IN_WIDTH: ping_storage_data_719 <= (fillup_transition == 1'b1) ? i_input_data[621 % IN_WIDTH] : ping_storage_data_719 ^ i_input_data[621 % IN_WIDTH];
                864 / IN_WIDTH: ping_storage_data_719 <= (fillup_transition == 1'b1) ? i_input_data[864 % IN_WIDTH] : ping_storage_data_719 ^ i_input_data[864 % IN_WIDTH];
                default: ping_storage_data_719 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_719;
                endcase
            end else begin
                case (input_count)
                132 / IN_WIDTH: pong_storage_data_719 <= (fillup_transition == 1'b1) ? i_input_data[132 % IN_WIDTH] : pong_storage_data_719 ^ i_input_data[132 % IN_WIDTH];
                262 / IN_WIDTH: pong_storage_data_719 <= (fillup_transition == 1'b1) ? i_input_data[262 % IN_WIDTH] : pong_storage_data_719 ^ i_input_data[262 % IN_WIDTH];
                621 / IN_WIDTH: pong_storage_data_719 <= (fillup_transition == 1'b1) ? i_input_data[621 % IN_WIDTH] : pong_storage_data_719 ^ i_input_data[621 % IN_WIDTH];
                864 / IN_WIDTH: pong_storage_data_719 <= (fillup_transition == 1'b1) ? i_input_data[864 % IN_WIDTH] : pong_storage_data_719 ^ i_input_data[864 % IN_WIDTH];
                default: pong_storage_data_719 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_719;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_719 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_719;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_719 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_719;
            end
        end
    end
end

logic ping_storage_data_720;
logic pong_storage_data_720;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_720 <= 1'b0;
        pong_storage_data_720 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                133 / IN_WIDTH: ping_storage_data_720 <= (fillup_transition == 1'b1) ? i_input_data[133 % IN_WIDTH] : ping_storage_data_720 ^ i_input_data[133 % IN_WIDTH];
                263 / IN_WIDTH: ping_storage_data_720 <= (fillup_transition == 1'b1) ? i_input_data[263 % IN_WIDTH] : ping_storage_data_720 ^ i_input_data[263 % IN_WIDTH];
                622 / IN_WIDTH: ping_storage_data_720 <= (fillup_transition == 1'b1) ? i_input_data[622 % IN_WIDTH] : ping_storage_data_720 ^ i_input_data[622 % IN_WIDTH];
                865 / IN_WIDTH: ping_storage_data_720 <= (fillup_transition == 1'b1) ? i_input_data[865 % IN_WIDTH] : ping_storage_data_720 ^ i_input_data[865 % IN_WIDTH];
                default: ping_storage_data_720 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_720;
                endcase
            end else begin
                case (input_count)
                133 / IN_WIDTH: pong_storage_data_720 <= (fillup_transition == 1'b1) ? i_input_data[133 % IN_WIDTH] : pong_storage_data_720 ^ i_input_data[133 % IN_WIDTH];
                263 / IN_WIDTH: pong_storage_data_720 <= (fillup_transition == 1'b1) ? i_input_data[263 % IN_WIDTH] : pong_storage_data_720 ^ i_input_data[263 % IN_WIDTH];
                622 / IN_WIDTH: pong_storage_data_720 <= (fillup_transition == 1'b1) ? i_input_data[622 % IN_WIDTH] : pong_storage_data_720 ^ i_input_data[622 % IN_WIDTH];
                865 / IN_WIDTH: pong_storage_data_720 <= (fillup_transition == 1'b1) ? i_input_data[865 % IN_WIDTH] : pong_storage_data_720 ^ i_input_data[865 % IN_WIDTH];
                default: pong_storage_data_720 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_720;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_720 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_720;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_720 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_720;
            end
        end
    end
end

logic ping_storage_data_721;
logic pong_storage_data_721;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_721 <= 1'b0;
        pong_storage_data_721 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                134 / IN_WIDTH: ping_storage_data_721 <= (fillup_transition == 1'b1) ? i_input_data[134 % IN_WIDTH] : ping_storage_data_721 ^ i_input_data[134 % IN_WIDTH];
                264 / IN_WIDTH: ping_storage_data_721 <= (fillup_transition == 1'b1) ? i_input_data[264 % IN_WIDTH] : ping_storage_data_721 ^ i_input_data[264 % IN_WIDTH];
                623 / IN_WIDTH: ping_storage_data_721 <= (fillup_transition == 1'b1) ? i_input_data[623 % IN_WIDTH] : ping_storage_data_721 ^ i_input_data[623 % IN_WIDTH];
                866 / IN_WIDTH: ping_storage_data_721 <= (fillup_transition == 1'b1) ? i_input_data[866 % IN_WIDTH] : ping_storage_data_721 ^ i_input_data[866 % IN_WIDTH];
                default: ping_storage_data_721 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_721;
                endcase
            end else begin
                case (input_count)
                134 / IN_WIDTH: pong_storage_data_721 <= (fillup_transition == 1'b1) ? i_input_data[134 % IN_WIDTH] : pong_storage_data_721 ^ i_input_data[134 % IN_WIDTH];
                264 / IN_WIDTH: pong_storage_data_721 <= (fillup_transition == 1'b1) ? i_input_data[264 % IN_WIDTH] : pong_storage_data_721 ^ i_input_data[264 % IN_WIDTH];
                623 / IN_WIDTH: pong_storage_data_721 <= (fillup_transition == 1'b1) ? i_input_data[623 % IN_WIDTH] : pong_storage_data_721 ^ i_input_data[623 % IN_WIDTH];
                866 / IN_WIDTH: pong_storage_data_721 <= (fillup_transition == 1'b1) ? i_input_data[866 % IN_WIDTH] : pong_storage_data_721 ^ i_input_data[866 % IN_WIDTH];
                default: pong_storage_data_721 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_721;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_721 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_721;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_721 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_721;
            end
        end
    end
end

logic ping_storage_data_722;
logic pong_storage_data_722;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_722 <= 1'b0;
        pong_storage_data_722 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                135 / IN_WIDTH: ping_storage_data_722 <= (fillup_transition == 1'b1) ? i_input_data[135 % IN_WIDTH] : ping_storage_data_722 ^ i_input_data[135 % IN_WIDTH];
                265 / IN_WIDTH: ping_storage_data_722 <= (fillup_transition == 1'b1) ? i_input_data[265 % IN_WIDTH] : ping_storage_data_722 ^ i_input_data[265 % IN_WIDTH];
                624 / IN_WIDTH: ping_storage_data_722 <= (fillup_transition == 1'b1) ? i_input_data[624 % IN_WIDTH] : ping_storage_data_722 ^ i_input_data[624 % IN_WIDTH];
                867 / IN_WIDTH: ping_storage_data_722 <= (fillup_transition == 1'b1) ? i_input_data[867 % IN_WIDTH] : ping_storage_data_722 ^ i_input_data[867 % IN_WIDTH];
                default: ping_storage_data_722 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_722;
                endcase
            end else begin
                case (input_count)
                135 / IN_WIDTH: pong_storage_data_722 <= (fillup_transition == 1'b1) ? i_input_data[135 % IN_WIDTH] : pong_storage_data_722 ^ i_input_data[135 % IN_WIDTH];
                265 / IN_WIDTH: pong_storage_data_722 <= (fillup_transition == 1'b1) ? i_input_data[265 % IN_WIDTH] : pong_storage_data_722 ^ i_input_data[265 % IN_WIDTH];
                624 / IN_WIDTH: pong_storage_data_722 <= (fillup_transition == 1'b1) ? i_input_data[624 % IN_WIDTH] : pong_storage_data_722 ^ i_input_data[624 % IN_WIDTH];
                867 / IN_WIDTH: pong_storage_data_722 <= (fillup_transition == 1'b1) ? i_input_data[867 % IN_WIDTH] : pong_storage_data_722 ^ i_input_data[867 % IN_WIDTH];
                default: pong_storage_data_722 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_722;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_722 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_722;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_722 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_722;
            end
        end
    end
end

logic ping_storage_data_723;
logic pong_storage_data_723;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_723 <= 1'b0;
        pong_storage_data_723 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                136 / IN_WIDTH: ping_storage_data_723 <= (fillup_transition == 1'b1) ? i_input_data[136 % IN_WIDTH] : ping_storage_data_723 ^ i_input_data[136 % IN_WIDTH];
                266 / IN_WIDTH: ping_storage_data_723 <= (fillup_transition == 1'b1) ? i_input_data[266 % IN_WIDTH] : ping_storage_data_723 ^ i_input_data[266 % IN_WIDTH];
                625 / IN_WIDTH: ping_storage_data_723 <= (fillup_transition == 1'b1) ? i_input_data[625 % IN_WIDTH] : ping_storage_data_723 ^ i_input_data[625 % IN_WIDTH];
                868 / IN_WIDTH: ping_storage_data_723 <= (fillup_transition == 1'b1) ? i_input_data[868 % IN_WIDTH] : ping_storage_data_723 ^ i_input_data[868 % IN_WIDTH];
                default: ping_storage_data_723 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_723;
                endcase
            end else begin
                case (input_count)
                136 / IN_WIDTH: pong_storage_data_723 <= (fillup_transition == 1'b1) ? i_input_data[136 % IN_WIDTH] : pong_storage_data_723 ^ i_input_data[136 % IN_WIDTH];
                266 / IN_WIDTH: pong_storage_data_723 <= (fillup_transition == 1'b1) ? i_input_data[266 % IN_WIDTH] : pong_storage_data_723 ^ i_input_data[266 % IN_WIDTH];
                625 / IN_WIDTH: pong_storage_data_723 <= (fillup_transition == 1'b1) ? i_input_data[625 % IN_WIDTH] : pong_storage_data_723 ^ i_input_data[625 % IN_WIDTH];
                868 / IN_WIDTH: pong_storage_data_723 <= (fillup_transition == 1'b1) ? i_input_data[868 % IN_WIDTH] : pong_storage_data_723 ^ i_input_data[868 % IN_WIDTH];
                default: pong_storage_data_723 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_723;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_723 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_723;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_723 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_723;
            end
        end
    end
end

logic ping_storage_data_724;
logic pong_storage_data_724;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_724 <= 1'b0;
        pong_storage_data_724 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                137 / IN_WIDTH: ping_storage_data_724 <= (fillup_transition == 1'b1) ? i_input_data[137 % IN_WIDTH] : ping_storage_data_724 ^ i_input_data[137 % IN_WIDTH];
                267 / IN_WIDTH: ping_storage_data_724 <= (fillup_transition == 1'b1) ? i_input_data[267 % IN_WIDTH] : ping_storage_data_724 ^ i_input_data[267 % IN_WIDTH];
                626 / IN_WIDTH: ping_storage_data_724 <= (fillup_transition == 1'b1) ? i_input_data[626 % IN_WIDTH] : ping_storage_data_724 ^ i_input_data[626 % IN_WIDTH];
                869 / IN_WIDTH: ping_storage_data_724 <= (fillup_transition == 1'b1) ? i_input_data[869 % IN_WIDTH] : ping_storage_data_724 ^ i_input_data[869 % IN_WIDTH];
                default: ping_storage_data_724 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_724;
                endcase
            end else begin
                case (input_count)
                137 / IN_WIDTH: pong_storage_data_724 <= (fillup_transition == 1'b1) ? i_input_data[137 % IN_WIDTH] : pong_storage_data_724 ^ i_input_data[137 % IN_WIDTH];
                267 / IN_WIDTH: pong_storage_data_724 <= (fillup_transition == 1'b1) ? i_input_data[267 % IN_WIDTH] : pong_storage_data_724 ^ i_input_data[267 % IN_WIDTH];
                626 / IN_WIDTH: pong_storage_data_724 <= (fillup_transition == 1'b1) ? i_input_data[626 % IN_WIDTH] : pong_storage_data_724 ^ i_input_data[626 % IN_WIDTH];
                869 / IN_WIDTH: pong_storage_data_724 <= (fillup_transition == 1'b1) ? i_input_data[869 % IN_WIDTH] : pong_storage_data_724 ^ i_input_data[869 % IN_WIDTH];
                default: pong_storage_data_724 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_724;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_724 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_724;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_724 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_724;
            end
        end
    end
end

logic ping_storage_data_725;
logic pong_storage_data_725;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_725 <= 1'b0;
        pong_storage_data_725 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                138 / IN_WIDTH: ping_storage_data_725 <= (fillup_transition == 1'b1) ? i_input_data[138 % IN_WIDTH] : ping_storage_data_725 ^ i_input_data[138 % IN_WIDTH];
                268 / IN_WIDTH: ping_storage_data_725 <= (fillup_transition == 1'b1) ? i_input_data[268 % IN_WIDTH] : ping_storage_data_725 ^ i_input_data[268 % IN_WIDTH];
                627 / IN_WIDTH: ping_storage_data_725 <= (fillup_transition == 1'b1) ? i_input_data[627 % IN_WIDTH] : ping_storage_data_725 ^ i_input_data[627 % IN_WIDTH];
                870 / IN_WIDTH: ping_storage_data_725 <= (fillup_transition == 1'b1) ? i_input_data[870 % IN_WIDTH] : ping_storage_data_725 ^ i_input_data[870 % IN_WIDTH];
                default: ping_storage_data_725 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_725;
                endcase
            end else begin
                case (input_count)
                138 / IN_WIDTH: pong_storage_data_725 <= (fillup_transition == 1'b1) ? i_input_data[138 % IN_WIDTH] : pong_storage_data_725 ^ i_input_data[138 % IN_WIDTH];
                268 / IN_WIDTH: pong_storage_data_725 <= (fillup_transition == 1'b1) ? i_input_data[268 % IN_WIDTH] : pong_storage_data_725 ^ i_input_data[268 % IN_WIDTH];
                627 / IN_WIDTH: pong_storage_data_725 <= (fillup_transition == 1'b1) ? i_input_data[627 % IN_WIDTH] : pong_storage_data_725 ^ i_input_data[627 % IN_WIDTH];
                870 / IN_WIDTH: pong_storage_data_725 <= (fillup_transition == 1'b1) ? i_input_data[870 % IN_WIDTH] : pong_storage_data_725 ^ i_input_data[870 % IN_WIDTH];
                default: pong_storage_data_725 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_725;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_725 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_725;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_725 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_725;
            end
        end
    end
end

logic ping_storage_data_726;
logic pong_storage_data_726;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_726 <= 1'b0;
        pong_storage_data_726 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                139 / IN_WIDTH: ping_storage_data_726 <= (fillup_transition == 1'b1) ? i_input_data[139 % IN_WIDTH] : ping_storage_data_726 ^ i_input_data[139 % IN_WIDTH];
                269 / IN_WIDTH: ping_storage_data_726 <= (fillup_transition == 1'b1) ? i_input_data[269 % IN_WIDTH] : ping_storage_data_726 ^ i_input_data[269 % IN_WIDTH];
                628 / IN_WIDTH: ping_storage_data_726 <= (fillup_transition == 1'b1) ? i_input_data[628 % IN_WIDTH] : ping_storage_data_726 ^ i_input_data[628 % IN_WIDTH];
                871 / IN_WIDTH: ping_storage_data_726 <= (fillup_transition == 1'b1) ? i_input_data[871 % IN_WIDTH] : ping_storage_data_726 ^ i_input_data[871 % IN_WIDTH];
                default: ping_storage_data_726 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_726;
                endcase
            end else begin
                case (input_count)
                139 / IN_WIDTH: pong_storage_data_726 <= (fillup_transition == 1'b1) ? i_input_data[139 % IN_WIDTH] : pong_storage_data_726 ^ i_input_data[139 % IN_WIDTH];
                269 / IN_WIDTH: pong_storage_data_726 <= (fillup_transition == 1'b1) ? i_input_data[269 % IN_WIDTH] : pong_storage_data_726 ^ i_input_data[269 % IN_WIDTH];
                628 / IN_WIDTH: pong_storage_data_726 <= (fillup_transition == 1'b1) ? i_input_data[628 % IN_WIDTH] : pong_storage_data_726 ^ i_input_data[628 % IN_WIDTH];
                871 / IN_WIDTH: pong_storage_data_726 <= (fillup_transition == 1'b1) ? i_input_data[871 % IN_WIDTH] : pong_storage_data_726 ^ i_input_data[871 % IN_WIDTH];
                default: pong_storage_data_726 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_726;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_726 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_726;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_726 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_726;
            end
        end
    end
end

logic ping_storage_data_727;
logic pong_storage_data_727;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_727 <= 1'b0;
        pong_storage_data_727 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                140 / IN_WIDTH: ping_storage_data_727 <= (fillup_transition == 1'b1) ? i_input_data[140 % IN_WIDTH] : ping_storage_data_727 ^ i_input_data[140 % IN_WIDTH];
                270 / IN_WIDTH: ping_storage_data_727 <= (fillup_transition == 1'b1) ? i_input_data[270 % IN_WIDTH] : ping_storage_data_727 ^ i_input_data[270 % IN_WIDTH];
                629 / IN_WIDTH: ping_storage_data_727 <= (fillup_transition == 1'b1) ? i_input_data[629 % IN_WIDTH] : ping_storage_data_727 ^ i_input_data[629 % IN_WIDTH];
                872 / IN_WIDTH: ping_storage_data_727 <= (fillup_transition == 1'b1) ? i_input_data[872 % IN_WIDTH] : ping_storage_data_727 ^ i_input_data[872 % IN_WIDTH];
                default: ping_storage_data_727 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_727;
                endcase
            end else begin
                case (input_count)
                140 / IN_WIDTH: pong_storage_data_727 <= (fillup_transition == 1'b1) ? i_input_data[140 % IN_WIDTH] : pong_storage_data_727 ^ i_input_data[140 % IN_WIDTH];
                270 / IN_WIDTH: pong_storage_data_727 <= (fillup_transition == 1'b1) ? i_input_data[270 % IN_WIDTH] : pong_storage_data_727 ^ i_input_data[270 % IN_WIDTH];
                629 / IN_WIDTH: pong_storage_data_727 <= (fillup_transition == 1'b1) ? i_input_data[629 % IN_WIDTH] : pong_storage_data_727 ^ i_input_data[629 % IN_WIDTH];
                872 / IN_WIDTH: pong_storage_data_727 <= (fillup_transition == 1'b1) ? i_input_data[872 % IN_WIDTH] : pong_storage_data_727 ^ i_input_data[872 % IN_WIDTH];
                default: pong_storage_data_727 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_727;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_727 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_727;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_727 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_727;
            end
        end
    end
end

logic ping_storage_data_728;
logic pong_storage_data_728;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_728 <= 1'b0;
        pong_storage_data_728 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                141 / IN_WIDTH: ping_storage_data_728 <= (fillup_transition == 1'b1) ? i_input_data[141 % IN_WIDTH] : ping_storage_data_728 ^ i_input_data[141 % IN_WIDTH];
                271 / IN_WIDTH: ping_storage_data_728 <= (fillup_transition == 1'b1) ? i_input_data[271 % IN_WIDTH] : ping_storage_data_728 ^ i_input_data[271 % IN_WIDTH];
                630 / IN_WIDTH: ping_storage_data_728 <= (fillup_transition == 1'b1) ? i_input_data[630 % IN_WIDTH] : ping_storage_data_728 ^ i_input_data[630 % IN_WIDTH];
                873 / IN_WIDTH: ping_storage_data_728 <= (fillup_transition == 1'b1) ? i_input_data[873 % IN_WIDTH] : ping_storage_data_728 ^ i_input_data[873 % IN_WIDTH];
                default: ping_storage_data_728 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_728;
                endcase
            end else begin
                case (input_count)
                141 / IN_WIDTH: pong_storage_data_728 <= (fillup_transition == 1'b1) ? i_input_data[141 % IN_WIDTH] : pong_storage_data_728 ^ i_input_data[141 % IN_WIDTH];
                271 / IN_WIDTH: pong_storage_data_728 <= (fillup_transition == 1'b1) ? i_input_data[271 % IN_WIDTH] : pong_storage_data_728 ^ i_input_data[271 % IN_WIDTH];
                630 / IN_WIDTH: pong_storage_data_728 <= (fillup_transition == 1'b1) ? i_input_data[630 % IN_WIDTH] : pong_storage_data_728 ^ i_input_data[630 % IN_WIDTH];
                873 / IN_WIDTH: pong_storage_data_728 <= (fillup_transition == 1'b1) ? i_input_data[873 % IN_WIDTH] : pong_storage_data_728 ^ i_input_data[873 % IN_WIDTH];
                default: pong_storage_data_728 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_728;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_728 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_728;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_728 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_728;
            end
        end
    end
end

logic ping_storage_data_729;
logic pong_storage_data_729;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_729 <= 1'b0;
        pong_storage_data_729 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                142 / IN_WIDTH: ping_storage_data_729 <= (fillup_transition == 1'b1) ? i_input_data[142 % IN_WIDTH] : ping_storage_data_729 ^ i_input_data[142 % IN_WIDTH];
                272 / IN_WIDTH: ping_storage_data_729 <= (fillup_transition == 1'b1) ? i_input_data[272 % IN_WIDTH] : ping_storage_data_729 ^ i_input_data[272 % IN_WIDTH];
                631 / IN_WIDTH: ping_storage_data_729 <= (fillup_transition == 1'b1) ? i_input_data[631 % IN_WIDTH] : ping_storage_data_729 ^ i_input_data[631 % IN_WIDTH];
                874 / IN_WIDTH: ping_storage_data_729 <= (fillup_transition == 1'b1) ? i_input_data[874 % IN_WIDTH] : ping_storage_data_729 ^ i_input_data[874 % IN_WIDTH];
                default: ping_storage_data_729 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_729;
                endcase
            end else begin
                case (input_count)
                142 / IN_WIDTH: pong_storage_data_729 <= (fillup_transition == 1'b1) ? i_input_data[142 % IN_WIDTH] : pong_storage_data_729 ^ i_input_data[142 % IN_WIDTH];
                272 / IN_WIDTH: pong_storage_data_729 <= (fillup_transition == 1'b1) ? i_input_data[272 % IN_WIDTH] : pong_storage_data_729 ^ i_input_data[272 % IN_WIDTH];
                631 / IN_WIDTH: pong_storage_data_729 <= (fillup_transition == 1'b1) ? i_input_data[631 % IN_WIDTH] : pong_storage_data_729 ^ i_input_data[631 % IN_WIDTH];
                874 / IN_WIDTH: pong_storage_data_729 <= (fillup_transition == 1'b1) ? i_input_data[874 % IN_WIDTH] : pong_storage_data_729 ^ i_input_data[874 % IN_WIDTH];
                default: pong_storage_data_729 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_729;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_729 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_729;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_729 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_729;
            end
        end
    end
end

logic ping_storage_data_730;
logic pong_storage_data_730;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_730 <= 1'b0;
        pong_storage_data_730 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                143 / IN_WIDTH: ping_storage_data_730 <= (fillup_transition == 1'b1) ? i_input_data[143 % IN_WIDTH] : ping_storage_data_730 ^ i_input_data[143 % IN_WIDTH];
                273 / IN_WIDTH: ping_storage_data_730 <= (fillup_transition == 1'b1) ? i_input_data[273 % IN_WIDTH] : ping_storage_data_730 ^ i_input_data[273 % IN_WIDTH];
                632 / IN_WIDTH: ping_storage_data_730 <= (fillup_transition == 1'b1) ? i_input_data[632 % IN_WIDTH] : ping_storage_data_730 ^ i_input_data[632 % IN_WIDTH];
                875 / IN_WIDTH: ping_storage_data_730 <= (fillup_transition == 1'b1) ? i_input_data[875 % IN_WIDTH] : ping_storage_data_730 ^ i_input_data[875 % IN_WIDTH];
                default: ping_storage_data_730 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_730;
                endcase
            end else begin
                case (input_count)
                143 / IN_WIDTH: pong_storage_data_730 <= (fillup_transition == 1'b1) ? i_input_data[143 % IN_WIDTH] : pong_storage_data_730 ^ i_input_data[143 % IN_WIDTH];
                273 / IN_WIDTH: pong_storage_data_730 <= (fillup_transition == 1'b1) ? i_input_data[273 % IN_WIDTH] : pong_storage_data_730 ^ i_input_data[273 % IN_WIDTH];
                632 / IN_WIDTH: pong_storage_data_730 <= (fillup_transition == 1'b1) ? i_input_data[632 % IN_WIDTH] : pong_storage_data_730 ^ i_input_data[632 % IN_WIDTH];
                875 / IN_WIDTH: pong_storage_data_730 <= (fillup_transition == 1'b1) ? i_input_data[875 % IN_WIDTH] : pong_storage_data_730 ^ i_input_data[875 % IN_WIDTH];
                default: pong_storage_data_730 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_730;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_730 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_730;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_730 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_730;
            end
        end
    end
end

logic ping_storage_data_731;
logic pong_storage_data_731;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_731 <= 1'b0;
        pong_storage_data_731 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                144 / IN_WIDTH: ping_storage_data_731 <= (fillup_transition == 1'b1) ? i_input_data[144 % IN_WIDTH] : ping_storage_data_731 ^ i_input_data[144 % IN_WIDTH];
                274 / IN_WIDTH: ping_storage_data_731 <= (fillup_transition == 1'b1) ? i_input_data[274 % IN_WIDTH] : ping_storage_data_731 ^ i_input_data[274 % IN_WIDTH];
                633 / IN_WIDTH: ping_storage_data_731 <= (fillup_transition == 1'b1) ? i_input_data[633 % IN_WIDTH] : ping_storage_data_731 ^ i_input_data[633 % IN_WIDTH];
                876 / IN_WIDTH: ping_storage_data_731 <= (fillup_transition == 1'b1) ? i_input_data[876 % IN_WIDTH] : ping_storage_data_731 ^ i_input_data[876 % IN_WIDTH];
                default: ping_storage_data_731 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_731;
                endcase
            end else begin
                case (input_count)
                144 / IN_WIDTH: pong_storage_data_731 <= (fillup_transition == 1'b1) ? i_input_data[144 % IN_WIDTH] : pong_storage_data_731 ^ i_input_data[144 % IN_WIDTH];
                274 / IN_WIDTH: pong_storage_data_731 <= (fillup_transition == 1'b1) ? i_input_data[274 % IN_WIDTH] : pong_storage_data_731 ^ i_input_data[274 % IN_WIDTH];
                633 / IN_WIDTH: pong_storage_data_731 <= (fillup_transition == 1'b1) ? i_input_data[633 % IN_WIDTH] : pong_storage_data_731 ^ i_input_data[633 % IN_WIDTH];
                876 / IN_WIDTH: pong_storage_data_731 <= (fillup_transition == 1'b1) ? i_input_data[876 % IN_WIDTH] : pong_storage_data_731 ^ i_input_data[876 % IN_WIDTH];
                default: pong_storage_data_731 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_731;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_731 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_731;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_731 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_731;
            end
        end
    end
end

logic ping_storage_data_732;
logic pong_storage_data_732;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_732 <= 1'b0;
        pong_storage_data_732 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                145 / IN_WIDTH: ping_storage_data_732 <= (fillup_transition == 1'b1) ? i_input_data[145 % IN_WIDTH] : ping_storage_data_732 ^ i_input_data[145 % IN_WIDTH];
                275 / IN_WIDTH: ping_storage_data_732 <= (fillup_transition == 1'b1) ? i_input_data[275 % IN_WIDTH] : ping_storage_data_732 ^ i_input_data[275 % IN_WIDTH];
                634 / IN_WIDTH: ping_storage_data_732 <= (fillup_transition == 1'b1) ? i_input_data[634 % IN_WIDTH] : ping_storage_data_732 ^ i_input_data[634 % IN_WIDTH];
                877 / IN_WIDTH: ping_storage_data_732 <= (fillup_transition == 1'b1) ? i_input_data[877 % IN_WIDTH] : ping_storage_data_732 ^ i_input_data[877 % IN_WIDTH];
                default: ping_storage_data_732 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_732;
                endcase
            end else begin
                case (input_count)
                145 / IN_WIDTH: pong_storage_data_732 <= (fillup_transition == 1'b1) ? i_input_data[145 % IN_WIDTH] : pong_storage_data_732 ^ i_input_data[145 % IN_WIDTH];
                275 / IN_WIDTH: pong_storage_data_732 <= (fillup_transition == 1'b1) ? i_input_data[275 % IN_WIDTH] : pong_storage_data_732 ^ i_input_data[275 % IN_WIDTH];
                634 / IN_WIDTH: pong_storage_data_732 <= (fillup_transition == 1'b1) ? i_input_data[634 % IN_WIDTH] : pong_storage_data_732 ^ i_input_data[634 % IN_WIDTH];
                877 / IN_WIDTH: pong_storage_data_732 <= (fillup_transition == 1'b1) ? i_input_data[877 % IN_WIDTH] : pong_storage_data_732 ^ i_input_data[877 % IN_WIDTH];
                default: pong_storage_data_732 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_732;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_732 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_732;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_732 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_732;
            end
        end
    end
end

logic ping_storage_data_733;
logic pong_storage_data_733;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_733 <= 1'b0;
        pong_storage_data_733 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                146 / IN_WIDTH: ping_storage_data_733 <= (fillup_transition == 1'b1) ? i_input_data[146 % IN_WIDTH] : ping_storage_data_733 ^ i_input_data[146 % IN_WIDTH];
                276 / IN_WIDTH: ping_storage_data_733 <= (fillup_transition == 1'b1) ? i_input_data[276 % IN_WIDTH] : ping_storage_data_733 ^ i_input_data[276 % IN_WIDTH];
                635 / IN_WIDTH: ping_storage_data_733 <= (fillup_transition == 1'b1) ? i_input_data[635 % IN_WIDTH] : ping_storage_data_733 ^ i_input_data[635 % IN_WIDTH];
                878 / IN_WIDTH: ping_storage_data_733 <= (fillup_transition == 1'b1) ? i_input_data[878 % IN_WIDTH] : ping_storage_data_733 ^ i_input_data[878 % IN_WIDTH];
                default: ping_storage_data_733 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_733;
                endcase
            end else begin
                case (input_count)
                146 / IN_WIDTH: pong_storage_data_733 <= (fillup_transition == 1'b1) ? i_input_data[146 % IN_WIDTH] : pong_storage_data_733 ^ i_input_data[146 % IN_WIDTH];
                276 / IN_WIDTH: pong_storage_data_733 <= (fillup_transition == 1'b1) ? i_input_data[276 % IN_WIDTH] : pong_storage_data_733 ^ i_input_data[276 % IN_WIDTH];
                635 / IN_WIDTH: pong_storage_data_733 <= (fillup_transition == 1'b1) ? i_input_data[635 % IN_WIDTH] : pong_storage_data_733 ^ i_input_data[635 % IN_WIDTH];
                878 / IN_WIDTH: pong_storage_data_733 <= (fillup_transition == 1'b1) ? i_input_data[878 % IN_WIDTH] : pong_storage_data_733 ^ i_input_data[878 % IN_WIDTH];
                default: pong_storage_data_733 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_733;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_733 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_733;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_733 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_733;
            end
        end
    end
end

logic ping_storage_data_734;
logic pong_storage_data_734;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_734 <= 1'b0;
        pong_storage_data_734 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                147 / IN_WIDTH: ping_storage_data_734 <= (fillup_transition == 1'b1) ? i_input_data[147 % IN_WIDTH] : ping_storage_data_734 ^ i_input_data[147 % IN_WIDTH];
                277 / IN_WIDTH: ping_storage_data_734 <= (fillup_transition == 1'b1) ? i_input_data[277 % IN_WIDTH] : ping_storage_data_734 ^ i_input_data[277 % IN_WIDTH];
                636 / IN_WIDTH: ping_storage_data_734 <= (fillup_transition == 1'b1) ? i_input_data[636 % IN_WIDTH] : ping_storage_data_734 ^ i_input_data[636 % IN_WIDTH];
                879 / IN_WIDTH: ping_storage_data_734 <= (fillup_transition == 1'b1) ? i_input_data[879 % IN_WIDTH] : ping_storage_data_734 ^ i_input_data[879 % IN_WIDTH];
                default: ping_storage_data_734 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_734;
                endcase
            end else begin
                case (input_count)
                147 / IN_WIDTH: pong_storage_data_734 <= (fillup_transition == 1'b1) ? i_input_data[147 % IN_WIDTH] : pong_storage_data_734 ^ i_input_data[147 % IN_WIDTH];
                277 / IN_WIDTH: pong_storage_data_734 <= (fillup_transition == 1'b1) ? i_input_data[277 % IN_WIDTH] : pong_storage_data_734 ^ i_input_data[277 % IN_WIDTH];
                636 / IN_WIDTH: pong_storage_data_734 <= (fillup_transition == 1'b1) ? i_input_data[636 % IN_WIDTH] : pong_storage_data_734 ^ i_input_data[636 % IN_WIDTH];
                879 / IN_WIDTH: pong_storage_data_734 <= (fillup_transition == 1'b1) ? i_input_data[879 % IN_WIDTH] : pong_storage_data_734 ^ i_input_data[879 % IN_WIDTH];
                default: pong_storage_data_734 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_734;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_734 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_734;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_734 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_734;
            end
        end
    end
end

logic ping_storage_data_735;
logic pong_storage_data_735;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_735 <= 1'b0;
        pong_storage_data_735 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                148 / IN_WIDTH: ping_storage_data_735 <= (fillup_transition == 1'b1) ? i_input_data[148 % IN_WIDTH] : ping_storage_data_735 ^ i_input_data[148 % IN_WIDTH];
                278 / IN_WIDTH: ping_storage_data_735 <= (fillup_transition == 1'b1) ? i_input_data[278 % IN_WIDTH] : ping_storage_data_735 ^ i_input_data[278 % IN_WIDTH];
                637 / IN_WIDTH: ping_storage_data_735 <= (fillup_transition == 1'b1) ? i_input_data[637 % IN_WIDTH] : ping_storage_data_735 ^ i_input_data[637 % IN_WIDTH];
                880 / IN_WIDTH: ping_storage_data_735 <= (fillup_transition == 1'b1) ? i_input_data[880 % IN_WIDTH] : ping_storage_data_735 ^ i_input_data[880 % IN_WIDTH];
                default: ping_storage_data_735 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_735;
                endcase
            end else begin
                case (input_count)
                148 / IN_WIDTH: pong_storage_data_735 <= (fillup_transition == 1'b1) ? i_input_data[148 % IN_WIDTH] : pong_storage_data_735 ^ i_input_data[148 % IN_WIDTH];
                278 / IN_WIDTH: pong_storage_data_735 <= (fillup_transition == 1'b1) ? i_input_data[278 % IN_WIDTH] : pong_storage_data_735 ^ i_input_data[278 % IN_WIDTH];
                637 / IN_WIDTH: pong_storage_data_735 <= (fillup_transition == 1'b1) ? i_input_data[637 % IN_WIDTH] : pong_storage_data_735 ^ i_input_data[637 % IN_WIDTH];
                880 / IN_WIDTH: pong_storage_data_735 <= (fillup_transition == 1'b1) ? i_input_data[880 % IN_WIDTH] : pong_storage_data_735 ^ i_input_data[880 % IN_WIDTH];
                default: pong_storage_data_735 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_735;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_735 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_735;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_735 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_735;
            end
        end
    end
end

logic ping_storage_data_736;
logic pong_storage_data_736;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_736 <= 1'b0;
        pong_storage_data_736 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                149 / IN_WIDTH: ping_storage_data_736 <= (fillup_transition == 1'b1) ? i_input_data[149 % IN_WIDTH] : ping_storage_data_736 ^ i_input_data[149 % IN_WIDTH];
                279 / IN_WIDTH: ping_storage_data_736 <= (fillup_transition == 1'b1) ? i_input_data[279 % IN_WIDTH] : ping_storage_data_736 ^ i_input_data[279 % IN_WIDTH];
                638 / IN_WIDTH: ping_storage_data_736 <= (fillup_transition == 1'b1) ? i_input_data[638 % IN_WIDTH] : ping_storage_data_736 ^ i_input_data[638 % IN_WIDTH];
                881 / IN_WIDTH: ping_storage_data_736 <= (fillup_transition == 1'b1) ? i_input_data[881 % IN_WIDTH] : ping_storage_data_736 ^ i_input_data[881 % IN_WIDTH];
                default: ping_storage_data_736 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_736;
                endcase
            end else begin
                case (input_count)
                149 / IN_WIDTH: pong_storage_data_736 <= (fillup_transition == 1'b1) ? i_input_data[149 % IN_WIDTH] : pong_storage_data_736 ^ i_input_data[149 % IN_WIDTH];
                279 / IN_WIDTH: pong_storage_data_736 <= (fillup_transition == 1'b1) ? i_input_data[279 % IN_WIDTH] : pong_storage_data_736 ^ i_input_data[279 % IN_WIDTH];
                638 / IN_WIDTH: pong_storage_data_736 <= (fillup_transition == 1'b1) ? i_input_data[638 % IN_WIDTH] : pong_storage_data_736 ^ i_input_data[638 % IN_WIDTH];
                881 / IN_WIDTH: pong_storage_data_736 <= (fillup_transition == 1'b1) ? i_input_data[881 % IN_WIDTH] : pong_storage_data_736 ^ i_input_data[881 % IN_WIDTH];
                default: pong_storage_data_736 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_736;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_736 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_736;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_736 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_736;
            end
        end
    end
end

logic ping_storage_data_737;
logic pong_storage_data_737;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_737 <= 1'b0;
        pong_storage_data_737 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                150 / IN_WIDTH: ping_storage_data_737 <= (fillup_transition == 1'b1) ? i_input_data[150 % IN_WIDTH] : ping_storage_data_737 ^ i_input_data[150 % IN_WIDTH];
                280 / IN_WIDTH: ping_storage_data_737 <= (fillup_transition == 1'b1) ? i_input_data[280 % IN_WIDTH] : ping_storage_data_737 ^ i_input_data[280 % IN_WIDTH];
                639 / IN_WIDTH: ping_storage_data_737 <= (fillup_transition == 1'b1) ? i_input_data[639 % IN_WIDTH] : ping_storage_data_737 ^ i_input_data[639 % IN_WIDTH];
                882 / IN_WIDTH: ping_storage_data_737 <= (fillup_transition == 1'b1) ? i_input_data[882 % IN_WIDTH] : ping_storage_data_737 ^ i_input_data[882 % IN_WIDTH];
                default: ping_storage_data_737 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_737;
                endcase
            end else begin
                case (input_count)
                150 / IN_WIDTH: pong_storage_data_737 <= (fillup_transition == 1'b1) ? i_input_data[150 % IN_WIDTH] : pong_storage_data_737 ^ i_input_data[150 % IN_WIDTH];
                280 / IN_WIDTH: pong_storage_data_737 <= (fillup_transition == 1'b1) ? i_input_data[280 % IN_WIDTH] : pong_storage_data_737 ^ i_input_data[280 % IN_WIDTH];
                639 / IN_WIDTH: pong_storage_data_737 <= (fillup_transition == 1'b1) ? i_input_data[639 % IN_WIDTH] : pong_storage_data_737 ^ i_input_data[639 % IN_WIDTH];
                882 / IN_WIDTH: pong_storage_data_737 <= (fillup_transition == 1'b1) ? i_input_data[882 % IN_WIDTH] : pong_storage_data_737 ^ i_input_data[882 % IN_WIDTH];
                default: pong_storage_data_737 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_737;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_737 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_737;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_737 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_737;
            end
        end
    end
end

logic ping_storage_data_738;
logic pong_storage_data_738;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_738 <= 1'b0;
        pong_storage_data_738 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                151 / IN_WIDTH: ping_storage_data_738 <= (fillup_transition == 1'b1) ? i_input_data[151 % IN_WIDTH] : ping_storage_data_738 ^ i_input_data[151 % IN_WIDTH];
                281 / IN_WIDTH: ping_storage_data_738 <= (fillup_transition == 1'b1) ? i_input_data[281 % IN_WIDTH] : ping_storage_data_738 ^ i_input_data[281 % IN_WIDTH];
                640 / IN_WIDTH: ping_storage_data_738 <= (fillup_transition == 1'b1) ? i_input_data[640 % IN_WIDTH] : ping_storage_data_738 ^ i_input_data[640 % IN_WIDTH];
                883 / IN_WIDTH: ping_storage_data_738 <= (fillup_transition == 1'b1) ? i_input_data[883 % IN_WIDTH] : ping_storage_data_738 ^ i_input_data[883 % IN_WIDTH];
                default: ping_storage_data_738 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_738;
                endcase
            end else begin
                case (input_count)
                151 / IN_WIDTH: pong_storage_data_738 <= (fillup_transition == 1'b1) ? i_input_data[151 % IN_WIDTH] : pong_storage_data_738 ^ i_input_data[151 % IN_WIDTH];
                281 / IN_WIDTH: pong_storage_data_738 <= (fillup_transition == 1'b1) ? i_input_data[281 % IN_WIDTH] : pong_storage_data_738 ^ i_input_data[281 % IN_WIDTH];
                640 / IN_WIDTH: pong_storage_data_738 <= (fillup_transition == 1'b1) ? i_input_data[640 % IN_WIDTH] : pong_storage_data_738 ^ i_input_data[640 % IN_WIDTH];
                883 / IN_WIDTH: pong_storage_data_738 <= (fillup_transition == 1'b1) ? i_input_data[883 % IN_WIDTH] : pong_storage_data_738 ^ i_input_data[883 % IN_WIDTH];
                default: pong_storage_data_738 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_738;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_738 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_738;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_738 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_738;
            end
        end
    end
end

logic ping_storage_data_739;
logic pong_storage_data_739;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_739 <= 1'b0;
        pong_storage_data_739 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                152 / IN_WIDTH: ping_storage_data_739 <= (fillup_transition == 1'b1) ? i_input_data[152 % IN_WIDTH] : ping_storage_data_739 ^ i_input_data[152 % IN_WIDTH];
                282 / IN_WIDTH: ping_storage_data_739 <= (fillup_transition == 1'b1) ? i_input_data[282 % IN_WIDTH] : ping_storage_data_739 ^ i_input_data[282 % IN_WIDTH];
                641 / IN_WIDTH: ping_storage_data_739 <= (fillup_transition == 1'b1) ? i_input_data[641 % IN_WIDTH] : ping_storage_data_739 ^ i_input_data[641 % IN_WIDTH];
                884 / IN_WIDTH: ping_storage_data_739 <= (fillup_transition == 1'b1) ? i_input_data[884 % IN_WIDTH] : ping_storage_data_739 ^ i_input_data[884 % IN_WIDTH];
                default: ping_storage_data_739 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_739;
                endcase
            end else begin
                case (input_count)
                152 / IN_WIDTH: pong_storage_data_739 <= (fillup_transition == 1'b1) ? i_input_data[152 % IN_WIDTH] : pong_storage_data_739 ^ i_input_data[152 % IN_WIDTH];
                282 / IN_WIDTH: pong_storage_data_739 <= (fillup_transition == 1'b1) ? i_input_data[282 % IN_WIDTH] : pong_storage_data_739 ^ i_input_data[282 % IN_WIDTH];
                641 / IN_WIDTH: pong_storage_data_739 <= (fillup_transition == 1'b1) ? i_input_data[641 % IN_WIDTH] : pong_storage_data_739 ^ i_input_data[641 % IN_WIDTH];
                884 / IN_WIDTH: pong_storage_data_739 <= (fillup_transition == 1'b1) ? i_input_data[884 % IN_WIDTH] : pong_storage_data_739 ^ i_input_data[884 % IN_WIDTH];
                default: pong_storage_data_739 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_739;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_739 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_739;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_739 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_739;
            end
        end
    end
end

logic ping_storage_data_740;
logic pong_storage_data_740;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_740 <= 1'b0;
        pong_storage_data_740 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                153 / IN_WIDTH: ping_storage_data_740 <= (fillup_transition == 1'b1) ? i_input_data[153 % IN_WIDTH] : ping_storage_data_740 ^ i_input_data[153 % IN_WIDTH];
                283 / IN_WIDTH: ping_storage_data_740 <= (fillup_transition == 1'b1) ? i_input_data[283 % IN_WIDTH] : ping_storage_data_740 ^ i_input_data[283 % IN_WIDTH];
                642 / IN_WIDTH: ping_storage_data_740 <= (fillup_transition == 1'b1) ? i_input_data[642 % IN_WIDTH] : ping_storage_data_740 ^ i_input_data[642 % IN_WIDTH];
                885 / IN_WIDTH: ping_storage_data_740 <= (fillup_transition == 1'b1) ? i_input_data[885 % IN_WIDTH] : ping_storage_data_740 ^ i_input_data[885 % IN_WIDTH];
                default: ping_storage_data_740 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_740;
                endcase
            end else begin
                case (input_count)
                153 / IN_WIDTH: pong_storage_data_740 <= (fillup_transition == 1'b1) ? i_input_data[153 % IN_WIDTH] : pong_storage_data_740 ^ i_input_data[153 % IN_WIDTH];
                283 / IN_WIDTH: pong_storage_data_740 <= (fillup_transition == 1'b1) ? i_input_data[283 % IN_WIDTH] : pong_storage_data_740 ^ i_input_data[283 % IN_WIDTH];
                642 / IN_WIDTH: pong_storage_data_740 <= (fillup_transition == 1'b1) ? i_input_data[642 % IN_WIDTH] : pong_storage_data_740 ^ i_input_data[642 % IN_WIDTH];
                885 / IN_WIDTH: pong_storage_data_740 <= (fillup_transition == 1'b1) ? i_input_data[885 % IN_WIDTH] : pong_storage_data_740 ^ i_input_data[885 % IN_WIDTH];
                default: pong_storage_data_740 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_740;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_740 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_740;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_740 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_740;
            end
        end
    end
end

logic ping_storage_data_741;
logic pong_storage_data_741;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_741 <= 1'b0;
        pong_storage_data_741 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                154 / IN_WIDTH: ping_storage_data_741 <= (fillup_transition == 1'b1) ? i_input_data[154 % IN_WIDTH] : ping_storage_data_741 ^ i_input_data[154 % IN_WIDTH];
                284 / IN_WIDTH: ping_storage_data_741 <= (fillup_transition == 1'b1) ? i_input_data[284 % IN_WIDTH] : ping_storage_data_741 ^ i_input_data[284 % IN_WIDTH];
                643 / IN_WIDTH: ping_storage_data_741 <= (fillup_transition == 1'b1) ? i_input_data[643 % IN_WIDTH] : ping_storage_data_741 ^ i_input_data[643 % IN_WIDTH];
                886 / IN_WIDTH: ping_storage_data_741 <= (fillup_transition == 1'b1) ? i_input_data[886 % IN_WIDTH] : ping_storage_data_741 ^ i_input_data[886 % IN_WIDTH];
                default: ping_storage_data_741 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_741;
                endcase
            end else begin
                case (input_count)
                154 / IN_WIDTH: pong_storage_data_741 <= (fillup_transition == 1'b1) ? i_input_data[154 % IN_WIDTH] : pong_storage_data_741 ^ i_input_data[154 % IN_WIDTH];
                284 / IN_WIDTH: pong_storage_data_741 <= (fillup_transition == 1'b1) ? i_input_data[284 % IN_WIDTH] : pong_storage_data_741 ^ i_input_data[284 % IN_WIDTH];
                643 / IN_WIDTH: pong_storage_data_741 <= (fillup_transition == 1'b1) ? i_input_data[643 % IN_WIDTH] : pong_storage_data_741 ^ i_input_data[643 % IN_WIDTH];
                886 / IN_WIDTH: pong_storage_data_741 <= (fillup_transition == 1'b1) ? i_input_data[886 % IN_WIDTH] : pong_storage_data_741 ^ i_input_data[886 % IN_WIDTH];
                default: pong_storage_data_741 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_741;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_741 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_741;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_741 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_741;
            end
        end
    end
end

logic ping_storage_data_742;
logic pong_storage_data_742;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_742 <= 1'b0;
        pong_storage_data_742 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                155 / IN_WIDTH: ping_storage_data_742 <= (fillup_transition == 1'b1) ? i_input_data[155 % IN_WIDTH] : ping_storage_data_742 ^ i_input_data[155 % IN_WIDTH];
                285 / IN_WIDTH: ping_storage_data_742 <= (fillup_transition == 1'b1) ? i_input_data[285 % IN_WIDTH] : ping_storage_data_742 ^ i_input_data[285 % IN_WIDTH];
                644 / IN_WIDTH: ping_storage_data_742 <= (fillup_transition == 1'b1) ? i_input_data[644 % IN_WIDTH] : ping_storage_data_742 ^ i_input_data[644 % IN_WIDTH];
                887 / IN_WIDTH: ping_storage_data_742 <= (fillup_transition == 1'b1) ? i_input_data[887 % IN_WIDTH] : ping_storage_data_742 ^ i_input_data[887 % IN_WIDTH];
                default: ping_storage_data_742 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_742;
                endcase
            end else begin
                case (input_count)
                155 / IN_WIDTH: pong_storage_data_742 <= (fillup_transition == 1'b1) ? i_input_data[155 % IN_WIDTH] : pong_storage_data_742 ^ i_input_data[155 % IN_WIDTH];
                285 / IN_WIDTH: pong_storage_data_742 <= (fillup_transition == 1'b1) ? i_input_data[285 % IN_WIDTH] : pong_storage_data_742 ^ i_input_data[285 % IN_WIDTH];
                644 / IN_WIDTH: pong_storage_data_742 <= (fillup_transition == 1'b1) ? i_input_data[644 % IN_WIDTH] : pong_storage_data_742 ^ i_input_data[644 % IN_WIDTH];
                887 / IN_WIDTH: pong_storage_data_742 <= (fillup_transition == 1'b1) ? i_input_data[887 % IN_WIDTH] : pong_storage_data_742 ^ i_input_data[887 % IN_WIDTH];
                default: pong_storage_data_742 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_742;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_742 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_742;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_742 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_742;
            end
        end
    end
end

logic ping_storage_data_743;
logic pong_storage_data_743;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_743 <= 1'b0;
        pong_storage_data_743 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                156 / IN_WIDTH: ping_storage_data_743 <= (fillup_transition == 1'b1) ? i_input_data[156 % IN_WIDTH] : ping_storage_data_743 ^ i_input_data[156 % IN_WIDTH];
                286 / IN_WIDTH: ping_storage_data_743 <= (fillup_transition == 1'b1) ? i_input_data[286 % IN_WIDTH] : ping_storage_data_743 ^ i_input_data[286 % IN_WIDTH];
                645 / IN_WIDTH: ping_storage_data_743 <= (fillup_transition == 1'b1) ? i_input_data[645 % IN_WIDTH] : ping_storage_data_743 ^ i_input_data[645 % IN_WIDTH];
                888 / IN_WIDTH: ping_storage_data_743 <= (fillup_transition == 1'b1) ? i_input_data[888 % IN_WIDTH] : ping_storage_data_743 ^ i_input_data[888 % IN_WIDTH];
                default: ping_storage_data_743 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_743;
                endcase
            end else begin
                case (input_count)
                156 / IN_WIDTH: pong_storage_data_743 <= (fillup_transition == 1'b1) ? i_input_data[156 % IN_WIDTH] : pong_storage_data_743 ^ i_input_data[156 % IN_WIDTH];
                286 / IN_WIDTH: pong_storage_data_743 <= (fillup_transition == 1'b1) ? i_input_data[286 % IN_WIDTH] : pong_storage_data_743 ^ i_input_data[286 % IN_WIDTH];
                645 / IN_WIDTH: pong_storage_data_743 <= (fillup_transition == 1'b1) ? i_input_data[645 % IN_WIDTH] : pong_storage_data_743 ^ i_input_data[645 % IN_WIDTH];
                888 / IN_WIDTH: pong_storage_data_743 <= (fillup_transition == 1'b1) ? i_input_data[888 % IN_WIDTH] : pong_storage_data_743 ^ i_input_data[888 % IN_WIDTH];
                default: pong_storage_data_743 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_743;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_743 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_743;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_743 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_743;
            end
        end
    end
end

logic ping_storage_data_744;
logic pong_storage_data_744;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_744 <= 1'b0;
        pong_storage_data_744 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                157 / IN_WIDTH: ping_storage_data_744 <= (fillup_transition == 1'b1) ? i_input_data[157 % IN_WIDTH] : ping_storage_data_744 ^ i_input_data[157 % IN_WIDTH];
                287 / IN_WIDTH: ping_storage_data_744 <= (fillup_transition == 1'b1) ? i_input_data[287 % IN_WIDTH] : ping_storage_data_744 ^ i_input_data[287 % IN_WIDTH];
                646 / IN_WIDTH: ping_storage_data_744 <= (fillup_transition == 1'b1) ? i_input_data[646 % IN_WIDTH] : ping_storage_data_744 ^ i_input_data[646 % IN_WIDTH];
                889 / IN_WIDTH: ping_storage_data_744 <= (fillup_transition == 1'b1) ? i_input_data[889 % IN_WIDTH] : ping_storage_data_744 ^ i_input_data[889 % IN_WIDTH];
                default: ping_storage_data_744 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_744;
                endcase
            end else begin
                case (input_count)
                157 / IN_WIDTH: pong_storage_data_744 <= (fillup_transition == 1'b1) ? i_input_data[157 % IN_WIDTH] : pong_storage_data_744 ^ i_input_data[157 % IN_WIDTH];
                287 / IN_WIDTH: pong_storage_data_744 <= (fillup_transition == 1'b1) ? i_input_data[287 % IN_WIDTH] : pong_storage_data_744 ^ i_input_data[287 % IN_WIDTH];
                646 / IN_WIDTH: pong_storage_data_744 <= (fillup_transition == 1'b1) ? i_input_data[646 % IN_WIDTH] : pong_storage_data_744 ^ i_input_data[646 % IN_WIDTH];
                889 / IN_WIDTH: pong_storage_data_744 <= (fillup_transition == 1'b1) ? i_input_data[889 % IN_WIDTH] : pong_storage_data_744 ^ i_input_data[889 % IN_WIDTH];
                default: pong_storage_data_744 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_744;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_744 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_744;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_744 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_744;
            end
        end
    end
end

logic ping_storage_data_745;
logic pong_storage_data_745;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_745 <= 1'b0;
        pong_storage_data_745 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                158 / IN_WIDTH: ping_storage_data_745 <= (fillup_transition == 1'b1) ? i_input_data[158 % IN_WIDTH] : ping_storage_data_745 ^ i_input_data[158 % IN_WIDTH];
                192 / IN_WIDTH: ping_storage_data_745 <= (fillup_transition == 1'b1) ? i_input_data[192 % IN_WIDTH] : ping_storage_data_745 ^ i_input_data[192 % IN_WIDTH];
                647 / IN_WIDTH: ping_storage_data_745 <= (fillup_transition == 1'b1) ? i_input_data[647 % IN_WIDTH] : ping_storage_data_745 ^ i_input_data[647 % IN_WIDTH];
                890 / IN_WIDTH: ping_storage_data_745 <= (fillup_transition == 1'b1) ? i_input_data[890 % IN_WIDTH] : ping_storage_data_745 ^ i_input_data[890 % IN_WIDTH];
                default: ping_storage_data_745 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_745;
                endcase
            end else begin
                case (input_count)
                158 / IN_WIDTH: pong_storage_data_745 <= (fillup_transition == 1'b1) ? i_input_data[158 % IN_WIDTH] : pong_storage_data_745 ^ i_input_data[158 % IN_WIDTH];
                192 / IN_WIDTH: pong_storage_data_745 <= (fillup_transition == 1'b1) ? i_input_data[192 % IN_WIDTH] : pong_storage_data_745 ^ i_input_data[192 % IN_WIDTH];
                647 / IN_WIDTH: pong_storage_data_745 <= (fillup_transition == 1'b1) ? i_input_data[647 % IN_WIDTH] : pong_storage_data_745 ^ i_input_data[647 % IN_WIDTH];
                890 / IN_WIDTH: pong_storage_data_745 <= (fillup_transition == 1'b1) ? i_input_data[890 % IN_WIDTH] : pong_storage_data_745 ^ i_input_data[890 % IN_WIDTH];
                default: pong_storage_data_745 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_745;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_745 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_745;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_745 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_745;
            end
        end
    end
end

logic ping_storage_data_746;
logic pong_storage_data_746;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_746 <= 1'b0;
        pong_storage_data_746 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                159 / IN_WIDTH: ping_storage_data_746 <= (fillup_transition == 1'b1) ? i_input_data[159 % IN_WIDTH] : ping_storage_data_746 ^ i_input_data[159 % IN_WIDTH];
                193 / IN_WIDTH: ping_storage_data_746 <= (fillup_transition == 1'b1) ? i_input_data[193 % IN_WIDTH] : ping_storage_data_746 ^ i_input_data[193 % IN_WIDTH];
                648 / IN_WIDTH: ping_storage_data_746 <= (fillup_transition == 1'b1) ? i_input_data[648 % IN_WIDTH] : ping_storage_data_746 ^ i_input_data[648 % IN_WIDTH];
                891 / IN_WIDTH: ping_storage_data_746 <= (fillup_transition == 1'b1) ? i_input_data[891 % IN_WIDTH] : ping_storage_data_746 ^ i_input_data[891 % IN_WIDTH];
                default: ping_storage_data_746 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_746;
                endcase
            end else begin
                case (input_count)
                159 / IN_WIDTH: pong_storage_data_746 <= (fillup_transition == 1'b1) ? i_input_data[159 % IN_WIDTH] : pong_storage_data_746 ^ i_input_data[159 % IN_WIDTH];
                193 / IN_WIDTH: pong_storage_data_746 <= (fillup_transition == 1'b1) ? i_input_data[193 % IN_WIDTH] : pong_storage_data_746 ^ i_input_data[193 % IN_WIDTH];
                648 / IN_WIDTH: pong_storage_data_746 <= (fillup_transition == 1'b1) ? i_input_data[648 % IN_WIDTH] : pong_storage_data_746 ^ i_input_data[648 % IN_WIDTH];
                891 / IN_WIDTH: pong_storage_data_746 <= (fillup_transition == 1'b1) ? i_input_data[891 % IN_WIDTH] : pong_storage_data_746 ^ i_input_data[891 % IN_WIDTH];
                default: pong_storage_data_746 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_746;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_746 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_746;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_746 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_746;
            end
        end
    end
end

logic ping_storage_data_747;
logic pong_storage_data_747;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_747 <= 1'b0;
        pong_storage_data_747 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                160 / IN_WIDTH: ping_storage_data_747 <= (fillup_transition == 1'b1) ? i_input_data[160 % IN_WIDTH] : ping_storage_data_747 ^ i_input_data[160 % IN_WIDTH];
                194 / IN_WIDTH: ping_storage_data_747 <= (fillup_transition == 1'b1) ? i_input_data[194 % IN_WIDTH] : ping_storage_data_747 ^ i_input_data[194 % IN_WIDTH];
                649 / IN_WIDTH: ping_storage_data_747 <= (fillup_transition == 1'b1) ? i_input_data[649 % IN_WIDTH] : ping_storage_data_747 ^ i_input_data[649 % IN_WIDTH];
                892 / IN_WIDTH: ping_storage_data_747 <= (fillup_transition == 1'b1) ? i_input_data[892 % IN_WIDTH] : ping_storage_data_747 ^ i_input_data[892 % IN_WIDTH];
                default: ping_storage_data_747 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_747;
                endcase
            end else begin
                case (input_count)
                160 / IN_WIDTH: pong_storage_data_747 <= (fillup_transition == 1'b1) ? i_input_data[160 % IN_WIDTH] : pong_storage_data_747 ^ i_input_data[160 % IN_WIDTH];
                194 / IN_WIDTH: pong_storage_data_747 <= (fillup_transition == 1'b1) ? i_input_data[194 % IN_WIDTH] : pong_storage_data_747 ^ i_input_data[194 % IN_WIDTH];
                649 / IN_WIDTH: pong_storage_data_747 <= (fillup_transition == 1'b1) ? i_input_data[649 % IN_WIDTH] : pong_storage_data_747 ^ i_input_data[649 % IN_WIDTH];
                892 / IN_WIDTH: pong_storage_data_747 <= (fillup_transition == 1'b1) ? i_input_data[892 % IN_WIDTH] : pong_storage_data_747 ^ i_input_data[892 % IN_WIDTH];
                default: pong_storage_data_747 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_747;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_747 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_747;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_747 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_747;
            end
        end
    end
end

logic ping_storage_data_748;
logic pong_storage_data_748;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_748 <= 1'b0;
        pong_storage_data_748 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                161 / IN_WIDTH: ping_storage_data_748 <= (fillup_transition == 1'b1) ? i_input_data[161 % IN_WIDTH] : ping_storage_data_748 ^ i_input_data[161 % IN_WIDTH];
                195 / IN_WIDTH: ping_storage_data_748 <= (fillup_transition == 1'b1) ? i_input_data[195 % IN_WIDTH] : ping_storage_data_748 ^ i_input_data[195 % IN_WIDTH];
                650 / IN_WIDTH: ping_storage_data_748 <= (fillup_transition == 1'b1) ? i_input_data[650 % IN_WIDTH] : ping_storage_data_748 ^ i_input_data[650 % IN_WIDTH];
                893 / IN_WIDTH: ping_storage_data_748 <= (fillup_transition == 1'b1) ? i_input_data[893 % IN_WIDTH] : ping_storage_data_748 ^ i_input_data[893 % IN_WIDTH];
                default: ping_storage_data_748 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_748;
                endcase
            end else begin
                case (input_count)
                161 / IN_WIDTH: pong_storage_data_748 <= (fillup_transition == 1'b1) ? i_input_data[161 % IN_WIDTH] : pong_storage_data_748 ^ i_input_data[161 % IN_WIDTH];
                195 / IN_WIDTH: pong_storage_data_748 <= (fillup_transition == 1'b1) ? i_input_data[195 % IN_WIDTH] : pong_storage_data_748 ^ i_input_data[195 % IN_WIDTH];
                650 / IN_WIDTH: pong_storage_data_748 <= (fillup_transition == 1'b1) ? i_input_data[650 % IN_WIDTH] : pong_storage_data_748 ^ i_input_data[650 % IN_WIDTH];
                893 / IN_WIDTH: pong_storage_data_748 <= (fillup_transition == 1'b1) ? i_input_data[893 % IN_WIDTH] : pong_storage_data_748 ^ i_input_data[893 % IN_WIDTH];
                default: pong_storage_data_748 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_748;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_748 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_748;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_748 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_748;
            end
        end
    end
end

logic ping_storage_data_749;
logic pong_storage_data_749;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_749 <= 1'b0;
        pong_storage_data_749 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                162 / IN_WIDTH: ping_storage_data_749 <= (fillup_transition == 1'b1) ? i_input_data[162 % IN_WIDTH] : ping_storage_data_749 ^ i_input_data[162 % IN_WIDTH];
                196 / IN_WIDTH: ping_storage_data_749 <= (fillup_transition == 1'b1) ? i_input_data[196 % IN_WIDTH] : ping_storage_data_749 ^ i_input_data[196 % IN_WIDTH];
                651 / IN_WIDTH: ping_storage_data_749 <= (fillup_transition == 1'b1) ? i_input_data[651 % IN_WIDTH] : ping_storage_data_749 ^ i_input_data[651 % IN_WIDTH];
                894 / IN_WIDTH: ping_storage_data_749 <= (fillup_transition == 1'b1) ? i_input_data[894 % IN_WIDTH] : ping_storage_data_749 ^ i_input_data[894 % IN_WIDTH];
                default: ping_storage_data_749 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_749;
                endcase
            end else begin
                case (input_count)
                162 / IN_WIDTH: pong_storage_data_749 <= (fillup_transition == 1'b1) ? i_input_data[162 % IN_WIDTH] : pong_storage_data_749 ^ i_input_data[162 % IN_WIDTH];
                196 / IN_WIDTH: pong_storage_data_749 <= (fillup_transition == 1'b1) ? i_input_data[196 % IN_WIDTH] : pong_storage_data_749 ^ i_input_data[196 % IN_WIDTH];
                651 / IN_WIDTH: pong_storage_data_749 <= (fillup_transition == 1'b1) ? i_input_data[651 % IN_WIDTH] : pong_storage_data_749 ^ i_input_data[651 % IN_WIDTH];
                894 / IN_WIDTH: pong_storage_data_749 <= (fillup_transition == 1'b1) ? i_input_data[894 % IN_WIDTH] : pong_storage_data_749 ^ i_input_data[894 % IN_WIDTH];
                default: pong_storage_data_749 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_749;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_749 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_749;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_749 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_749;
            end
        end
    end
end

logic ping_storage_data_750;
logic pong_storage_data_750;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_750 <= 1'b0;
        pong_storage_data_750 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                163 / IN_WIDTH: ping_storage_data_750 <= (fillup_transition == 1'b1) ? i_input_data[163 % IN_WIDTH] : ping_storage_data_750 ^ i_input_data[163 % IN_WIDTH];
                197 / IN_WIDTH: ping_storage_data_750 <= (fillup_transition == 1'b1) ? i_input_data[197 % IN_WIDTH] : ping_storage_data_750 ^ i_input_data[197 % IN_WIDTH];
                652 / IN_WIDTH: ping_storage_data_750 <= (fillup_transition == 1'b1) ? i_input_data[652 % IN_WIDTH] : ping_storage_data_750 ^ i_input_data[652 % IN_WIDTH];
                895 / IN_WIDTH: ping_storage_data_750 <= (fillup_transition == 1'b1) ? i_input_data[895 % IN_WIDTH] : ping_storage_data_750 ^ i_input_data[895 % IN_WIDTH];
                default: ping_storage_data_750 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_750;
                endcase
            end else begin
                case (input_count)
                163 / IN_WIDTH: pong_storage_data_750 <= (fillup_transition == 1'b1) ? i_input_data[163 % IN_WIDTH] : pong_storage_data_750 ^ i_input_data[163 % IN_WIDTH];
                197 / IN_WIDTH: pong_storage_data_750 <= (fillup_transition == 1'b1) ? i_input_data[197 % IN_WIDTH] : pong_storage_data_750 ^ i_input_data[197 % IN_WIDTH];
                652 / IN_WIDTH: pong_storage_data_750 <= (fillup_transition == 1'b1) ? i_input_data[652 % IN_WIDTH] : pong_storage_data_750 ^ i_input_data[652 % IN_WIDTH];
                895 / IN_WIDTH: pong_storage_data_750 <= (fillup_transition == 1'b1) ? i_input_data[895 % IN_WIDTH] : pong_storage_data_750 ^ i_input_data[895 % IN_WIDTH];
                default: pong_storage_data_750 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_750;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_750 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_750;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_750 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_750;
            end
        end
    end
end

logic ping_storage_data_751;
logic pong_storage_data_751;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_751 <= 1'b0;
        pong_storage_data_751 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                164 / IN_WIDTH: ping_storage_data_751 <= (fillup_transition == 1'b1) ? i_input_data[164 % IN_WIDTH] : ping_storage_data_751 ^ i_input_data[164 % IN_WIDTH];
                198 / IN_WIDTH: ping_storage_data_751 <= (fillup_transition == 1'b1) ? i_input_data[198 % IN_WIDTH] : ping_storage_data_751 ^ i_input_data[198 % IN_WIDTH];
                653 / IN_WIDTH: ping_storage_data_751 <= (fillup_transition == 1'b1) ? i_input_data[653 % IN_WIDTH] : ping_storage_data_751 ^ i_input_data[653 % IN_WIDTH];
                896 / IN_WIDTH: ping_storage_data_751 <= (fillup_transition == 1'b1) ? i_input_data[896 % IN_WIDTH] : ping_storage_data_751 ^ i_input_data[896 % IN_WIDTH];
                default: ping_storage_data_751 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_751;
                endcase
            end else begin
                case (input_count)
                164 / IN_WIDTH: pong_storage_data_751 <= (fillup_transition == 1'b1) ? i_input_data[164 % IN_WIDTH] : pong_storage_data_751 ^ i_input_data[164 % IN_WIDTH];
                198 / IN_WIDTH: pong_storage_data_751 <= (fillup_transition == 1'b1) ? i_input_data[198 % IN_WIDTH] : pong_storage_data_751 ^ i_input_data[198 % IN_WIDTH];
                653 / IN_WIDTH: pong_storage_data_751 <= (fillup_transition == 1'b1) ? i_input_data[653 % IN_WIDTH] : pong_storage_data_751 ^ i_input_data[653 % IN_WIDTH];
                896 / IN_WIDTH: pong_storage_data_751 <= (fillup_transition == 1'b1) ? i_input_data[896 % IN_WIDTH] : pong_storage_data_751 ^ i_input_data[896 % IN_WIDTH];
                default: pong_storage_data_751 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_751;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_751 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_751;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_751 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_751;
            end
        end
    end
end

logic ping_storage_data_752;
logic pong_storage_data_752;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_752 <= 1'b0;
        pong_storage_data_752 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                165 / IN_WIDTH: ping_storage_data_752 <= (fillup_transition == 1'b1) ? i_input_data[165 % IN_WIDTH] : ping_storage_data_752 ^ i_input_data[165 % IN_WIDTH];
                199 / IN_WIDTH: ping_storage_data_752 <= (fillup_transition == 1'b1) ? i_input_data[199 % IN_WIDTH] : ping_storage_data_752 ^ i_input_data[199 % IN_WIDTH];
                654 / IN_WIDTH: ping_storage_data_752 <= (fillup_transition == 1'b1) ? i_input_data[654 % IN_WIDTH] : ping_storage_data_752 ^ i_input_data[654 % IN_WIDTH];
                897 / IN_WIDTH: ping_storage_data_752 <= (fillup_transition == 1'b1) ? i_input_data[897 % IN_WIDTH] : ping_storage_data_752 ^ i_input_data[897 % IN_WIDTH];
                default: ping_storage_data_752 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_752;
                endcase
            end else begin
                case (input_count)
                165 / IN_WIDTH: pong_storage_data_752 <= (fillup_transition == 1'b1) ? i_input_data[165 % IN_WIDTH] : pong_storage_data_752 ^ i_input_data[165 % IN_WIDTH];
                199 / IN_WIDTH: pong_storage_data_752 <= (fillup_transition == 1'b1) ? i_input_data[199 % IN_WIDTH] : pong_storage_data_752 ^ i_input_data[199 % IN_WIDTH];
                654 / IN_WIDTH: pong_storage_data_752 <= (fillup_transition == 1'b1) ? i_input_data[654 % IN_WIDTH] : pong_storage_data_752 ^ i_input_data[654 % IN_WIDTH];
                897 / IN_WIDTH: pong_storage_data_752 <= (fillup_transition == 1'b1) ? i_input_data[897 % IN_WIDTH] : pong_storage_data_752 ^ i_input_data[897 % IN_WIDTH];
                default: pong_storage_data_752 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_752;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_752 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_752;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_752 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_752;
            end
        end
    end
end

logic ping_storage_data_753;
logic pong_storage_data_753;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_753 <= 1'b0;
        pong_storage_data_753 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                166 / IN_WIDTH: ping_storage_data_753 <= (fillup_transition == 1'b1) ? i_input_data[166 % IN_WIDTH] : ping_storage_data_753 ^ i_input_data[166 % IN_WIDTH];
                200 / IN_WIDTH: ping_storage_data_753 <= (fillup_transition == 1'b1) ? i_input_data[200 % IN_WIDTH] : ping_storage_data_753 ^ i_input_data[200 % IN_WIDTH];
                655 / IN_WIDTH: ping_storage_data_753 <= (fillup_transition == 1'b1) ? i_input_data[655 % IN_WIDTH] : ping_storage_data_753 ^ i_input_data[655 % IN_WIDTH];
                898 / IN_WIDTH: ping_storage_data_753 <= (fillup_transition == 1'b1) ? i_input_data[898 % IN_WIDTH] : ping_storage_data_753 ^ i_input_data[898 % IN_WIDTH];
                default: ping_storage_data_753 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_753;
                endcase
            end else begin
                case (input_count)
                166 / IN_WIDTH: pong_storage_data_753 <= (fillup_transition == 1'b1) ? i_input_data[166 % IN_WIDTH] : pong_storage_data_753 ^ i_input_data[166 % IN_WIDTH];
                200 / IN_WIDTH: pong_storage_data_753 <= (fillup_transition == 1'b1) ? i_input_data[200 % IN_WIDTH] : pong_storage_data_753 ^ i_input_data[200 % IN_WIDTH];
                655 / IN_WIDTH: pong_storage_data_753 <= (fillup_transition == 1'b1) ? i_input_data[655 % IN_WIDTH] : pong_storage_data_753 ^ i_input_data[655 % IN_WIDTH];
                898 / IN_WIDTH: pong_storage_data_753 <= (fillup_transition == 1'b1) ? i_input_data[898 % IN_WIDTH] : pong_storage_data_753 ^ i_input_data[898 % IN_WIDTH];
                default: pong_storage_data_753 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_753;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_753 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_753;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_753 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_753;
            end
        end
    end
end

logic ping_storage_data_754;
logic pong_storage_data_754;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_754 <= 1'b0;
        pong_storage_data_754 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                167 / IN_WIDTH: ping_storage_data_754 <= (fillup_transition == 1'b1) ? i_input_data[167 % IN_WIDTH] : ping_storage_data_754 ^ i_input_data[167 % IN_WIDTH];
                201 / IN_WIDTH: ping_storage_data_754 <= (fillup_transition == 1'b1) ? i_input_data[201 % IN_WIDTH] : ping_storage_data_754 ^ i_input_data[201 % IN_WIDTH];
                656 / IN_WIDTH: ping_storage_data_754 <= (fillup_transition == 1'b1) ? i_input_data[656 % IN_WIDTH] : ping_storage_data_754 ^ i_input_data[656 % IN_WIDTH];
                899 / IN_WIDTH: ping_storage_data_754 <= (fillup_transition == 1'b1) ? i_input_data[899 % IN_WIDTH] : ping_storage_data_754 ^ i_input_data[899 % IN_WIDTH];
                default: ping_storage_data_754 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_754;
                endcase
            end else begin
                case (input_count)
                167 / IN_WIDTH: pong_storage_data_754 <= (fillup_transition == 1'b1) ? i_input_data[167 % IN_WIDTH] : pong_storage_data_754 ^ i_input_data[167 % IN_WIDTH];
                201 / IN_WIDTH: pong_storage_data_754 <= (fillup_transition == 1'b1) ? i_input_data[201 % IN_WIDTH] : pong_storage_data_754 ^ i_input_data[201 % IN_WIDTH];
                656 / IN_WIDTH: pong_storage_data_754 <= (fillup_transition == 1'b1) ? i_input_data[656 % IN_WIDTH] : pong_storage_data_754 ^ i_input_data[656 % IN_WIDTH];
                899 / IN_WIDTH: pong_storage_data_754 <= (fillup_transition == 1'b1) ? i_input_data[899 % IN_WIDTH] : pong_storage_data_754 ^ i_input_data[899 % IN_WIDTH];
                default: pong_storage_data_754 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_754;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_754 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_754;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_754 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_754;
            end
        end
    end
end

logic ping_storage_data_755;
logic pong_storage_data_755;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_755 <= 1'b0;
        pong_storage_data_755 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                168 / IN_WIDTH: ping_storage_data_755 <= (fillup_transition == 1'b1) ? i_input_data[168 % IN_WIDTH] : ping_storage_data_755 ^ i_input_data[168 % IN_WIDTH];
                202 / IN_WIDTH: ping_storage_data_755 <= (fillup_transition == 1'b1) ? i_input_data[202 % IN_WIDTH] : ping_storage_data_755 ^ i_input_data[202 % IN_WIDTH];
                657 / IN_WIDTH: ping_storage_data_755 <= (fillup_transition == 1'b1) ? i_input_data[657 % IN_WIDTH] : ping_storage_data_755 ^ i_input_data[657 % IN_WIDTH];
                900 / IN_WIDTH: ping_storage_data_755 <= (fillup_transition == 1'b1) ? i_input_data[900 % IN_WIDTH] : ping_storage_data_755 ^ i_input_data[900 % IN_WIDTH];
                default: ping_storage_data_755 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_755;
                endcase
            end else begin
                case (input_count)
                168 / IN_WIDTH: pong_storage_data_755 <= (fillup_transition == 1'b1) ? i_input_data[168 % IN_WIDTH] : pong_storage_data_755 ^ i_input_data[168 % IN_WIDTH];
                202 / IN_WIDTH: pong_storage_data_755 <= (fillup_transition == 1'b1) ? i_input_data[202 % IN_WIDTH] : pong_storage_data_755 ^ i_input_data[202 % IN_WIDTH];
                657 / IN_WIDTH: pong_storage_data_755 <= (fillup_transition == 1'b1) ? i_input_data[657 % IN_WIDTH] : pong_storage_data_755 ^ i_input_data[657 % IN_WIDTH];
                900 / IN_WIDTH: pong_storage_data_755 <= (fillup_transition == 1'b1) ? i_input_data[900 % IN_WIDTH] : pong_storage_data_755 ^ i_input_data[900 % IN_WIDTH];
                default: pong_storage_data_755 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_755;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_755 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_755;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_755 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_755;
            end
        end
    end
end

logic ping_storage_data_756;
logic pong_storage_data_756;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_756 <= 1'b0;
        pong_storage_data_756 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                169 / IN_WIDTH: ping_storage_data_756 <= (fillup_transition == 1'b1) ? i_input_data[169 % IN_WIDTH] : ping_storage_data_756 ^ i_input_data[169 % IN_WIDTH];
                203 / IN_WIDTH: ping_storage_data_756 <= (fillup_transition == 1'b1) ? i_input_data[203 % IN_WIDTH] : ping_storage_data_756 ^ i_input_data[203 % IN_WIDTH];
                658 / IN_WIDTH: ping_storage_data_756 <= (fillup_transition == 1'b1) ? i_input_data[658 % IN_WIDTH] : ping_storage_data_756 ^ i_input_data[658 % IN_WIDTH];
                901 / IN_WIDTH: ping_storage_data_756 <= (fillup_transition == 1'b1) ? i_input_data[901 % IN_WIDTH] : ping_storage_data_756 ^ i_input_data[901 % IN_WIDTH];
                default: ping_storage_data_756 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_756;
                endcase
            end else begin
                case (input_count)
                169 / IN_WIDTH: pong_storage_data_756 <= (fillup_transition == 1'b1) ? i_input_data[169 % IN_WIDTH] : pong_storage_data_756 ^ i_input_data[169 % IN_WIDTH];
                203 / IN_WIDTH: pong_storage_data_756 <= (fillup_transition == 1'b1) ? i_input_data[203 % IN_WIDTH] : pong_storage_data_756 ^ i_input_data[203 % IN_WIDTH];
                658 / IN_WIDTH: pong_storage_data_756 <= (fillup_transition == 1'b1) ? i_input_data[658 % IN_WIDTH] : pong_storage_data_756 ^ i_input_data[658 % IN_WIDTH];
                901 / IN_WIDTH: pong_storage_data_756 <= (fillup_transition == 1'b1) ? i_input_data[901 % IN_WIDTH] : pong_storage_data_756 ^ i_input_data[901 % IN_WIDTH];
                default: pong_storage_data_756 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_756;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_756 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_756;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_756 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_756;
            end
        end
    end
end

logic ping_storage_data_757;
logic pong_storage_data_757;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_757 <= 1'b0;
        pong_storage_data_757 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                170 / IN_WIDTH: ping_storage_data_757 <= (fillup_transition == 1'b1) ? i_input_data[170 % IN_WIDTH] : ping_storage_data_757 ^ i_input_data[170 % IN_WIDTH];
                204 / IN_WIDTH: ping_storage_data_757 <= (fillup_transition == 1'b1) ? i_input_data[204 % IN_WIDTH] : ping_storage_data_757 ^ i_input_data[204 % IN_WIDTH];
                659 / IN_WIDTH: ping_storage_data_757 <= (fillup_transition == 1'b1) ? i_input_data[659 % IN_WIDTH] : ping_storage_data_757 ^ i_input_data[659 % IN_WIDTH];
                902 / IN_WIDTH: ping_storage_data_757 <= (fillup_transition == 1'b1) ? i_input_data[902 % IN_WIDTH] : ping_storage_data_757 ^ i_input_data[902 % IN_WIDTH];
                default: ping_storage_data_757 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_757;
                endcase
            end else begin
                case (input_count)
                170 / IN_WIDTH: pong_storage_data_757 <= (fillup_transition == 1'b1) ? i_input_data[170 % IN_WIDTH] : pong_storage_data_757 ^ i_input_data[170 % IN_WIDTH];
                204 / IN_WIDTH: pong_storage_data_757 <= (fillup_transition == 1'b1) ? i_input_data[204 % IN_WIDTH] : pong_storage_data_757 ^ i_input_data[204 % IN_WIDTH];
                659 / IN_WIDTH: pong_storage_data_757 <= (fillup_transition == 1'b1) ? i_input_data[659 % IN_WIDTH] : pong_storage_data_757 ^ i_input_data[659 % IN_WIDTH];
                902 / IN_WIDTH: pong_storage_data_757 <= (fillup_transition == 1'b1) ? i_input_data[902 % IN_WIDTH] : pong_storage_data_757 ^ i_input_data[902 % IN_WIDTH];
                default: pong_storage_data_757 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_757;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_757 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_757;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_757 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_757;
            end
        end
    end
end

logic ping_storage_data_758;
logic pong_storage_data_758;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_758 <= 1'b0;
        pong_storage_data_758 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                171 / IN_WIDTH: ping_storage_data_758 <= (fillup_transition == 1'b1) ? i_input_data[171 % IN_WIDTH] : ping_storage_data_758 ^ i_input_data[171 % IN_WIDTH];
                205 / IN_WIDTH: ping_storage_data_758 <= (fillup_transition == 1'b1) ? i_input_data[205 % IN_WIDTH] : ping_storage_data_758 ^ i_input_data[205 % IN_WIDTH];
                660 / IN_WIDTH: ping_storage_data_758 <= (fillup_transition == 1'b1) ? i_input_data[660 % IN_WIDTH] : ping_storage_data_758 ^ i_input_data[660 % IN_WIDTH];
                903 / IN_WIDTH: ping_storage_data_758 <= (fillup_transition == 1'b1) ? i_input_data[903 % IN_WIDTH] : ping_storage_data_758 ^ i_input_data[903 % IN_WIDTH];
                default: ping_storage_data_758 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_758;
                endcase
            end else begin
                case (input_count)
                171 / IN_WIDTH: pong_storage_data_758 <= (fillup_transition == 1'b1) ? i_input_data[171 % IN_WIDTH] : pong_storage_data_758 ^ i_input_data[171 % IN_WIDTH];
                205 / IN_WIDTH: pong_storage_data_758 <= (fillup_transition == 1'b1) ? i_input_data[205 % IN_WIDTH] : pong_storage_data_758 ^ i_input_data[205 % IN_WIDTH];
                660 / IN_WIDTH: pong_storage_data_758 <= (fillup_transition == 1'b1) ? i_input_data[660 % IN_WIDTH] : pong_storage_data_758 ^ i_input_data[660 % IN_WIDTH];
                903 / IN_WIDTH: pong_storage_data_758 <= (fillup_transition == 1'b1) ? i_input_data[903 % IN_WIDTH] : pong_storage_data_758 ^ i_input_data[903 % IN_WIDTH];
                default: pong_storage_data_758 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_758;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_758 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_758;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_758 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_758;
            end
        end
    end
end

logic ping_storage_data_759;
logic pong_storage_data_759;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_759 <= 1'b0;
        pong_storage_data_759 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                172 / IN_WIDTH: ping_storage_data_759 <= (fillup_transition == 1'b1) ? i_input_data[172 % IN_WIDTH] : ping_storage_data_759 ^ i_input_data[172 % IN_WIDTH];
                206 / IN_WIDTH: ping_storage_data_759 <= (fillup_transition == 1'b1) ? i_input_data[206 % IN_WIDTH] : ping_storage_data_759 ^ i_input_data[206 % IN_WIDTH];
                661 / IN_WIDTH: ping_storage_data_759 <= (fillup_transition == 1'b1) ? i_input_data[661 % IN_WIDTH] : ping_storage_data_759 ^ i_input_data[661 % IN_WIDTH];
                904 / IN_WIDTH: ping_storage_data_759 <= (fillup_transition == 1'b1) ? i_input_data[904 % IN_WIDTH] : ping_storage_data_759 ^ i_input_data[904 % IN_WIDTH];
                default: ping_storage_data_759 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_759;
                endcase
            end else begin
                case (input_count)
                172 / IN_WIDTH: pong_storage_data_759 <= (fillup_transition == 1'b1) ? i_input_data[172 % IN_WIDTH] : pong_storage_data_759 ^ i_input_data[172 % IN_WIDTH];
                206 / IN_WIDTH: pong_storage_data_759 <= (fillup_transition == 1'b1) ? i_input_data[206 % IN_WIDTH] : pong_storage_data_759 ^ i_input_data[206 % IN_WIDTH];
                661 / IN_WIDTH: pong_storage_data_759 <= (fillup_transition == 1'b1) ? i_input_data[661 % IN_WIDTH] : pong_storage_data_759 ^ i_input_data[661 % IN_WIDTH];
                904 / IN_WIDTH: pong_storage_data_759 <= (fillup_transition == 1'b1) ? i_input_data[904 % IN_WIDTH] : pong_storage_data_759 ^ i_input_data[904 % IN_WIDTH];
                default: pong_storage_data_759 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_759;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_759 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_759;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_759 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_759;
            end
        end
    end
end

logic ping_storage_data_760;
logic pong_storage_data_760;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_760 <= 1'b0;
        pong_storage_data_760 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                173 / IN_WIDTH: ping_storage_data_760 <= (fillup_transition == 1'b1) ? i_input_data[173 % IN_WIDTH] : ping_storage_data_760 ^ i_input_data[173 % IN_WIDTH];
                207 / IN_WIDTH: ping_storage_data_760 <= (fillup_transition == 1'b1) ? i_input_data[207 % IN_WIDTH] : ping_storage_data_760 ^ i_input_data[207 % IN_WIDTH];
                662 / IN_WIDTH: ping_storage_data_760 <= (fillup_transition == 1'b1) ? i_input_data[662 % IN_WIDTH] : ping_storage_data_760 ^ i_input_data[662 % IN_WIDTH];
                905 / IN_WIDTH: ping_storage_data_760 <= (fillup_transition == 1'b1) ? i_input_data[905 % IN_WIDTH] : ping_storage_data_760 ^ i_input_data[905 % IN_WIDTH];
                default: ping_storage_data_760 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_760;
                endcase
            end else begin
                case (input_count)
                173 / IN_WIDTH: pong_storage_data_760 <= (fillup_transition == 1'b1) ? i_input_data[173 % IN_WIDTH] : pong_storage_data_760 ^ i_input_data[173 % IN_WIDTH];
                207 / IN_WIDTH: pong_storage_data_760 <= (fillup_transition == 1'b1) ? i_input_data[207 % IN_WIDTH] : pong_storage_data_760 ^ i_input_data[207 % IN_WIDTH];
                662 / IN_WIDTH: pong_storage_data_760 <= (fillup_transition == 1'b1) ? i_input_data[662 % IN_WIDTH] : pong_storage_data_760 ^ i_input_data[662 % IN_WIDTH];
                905 / IN_WIDTH: pong_storage_data_760 <= (fillup_transition == 1'b1) ? i_input_data[905 % IN_WIDTH] : pong_storage_data_760 ^ i_input_data[905 % IN_WIDTH];
                default: pong_storage_data_760 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_760;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_760 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_760;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_760 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_760;
            end
        end
    end
end

logic ping_storage_data_761;
logic pong_storage_data_761;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_761 <= 1'b0;
        pong_storage_data_761 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                174 / IN_WIDTH: ping_storage_data_761 <= (fillup_transition == 1'b1) ? i_input_data[174 % IN_WIDTH] : ping_storage_data_761 ^ i_input_data[174 % IN_WIDTH];
                208 / IN_WIDTH: ping_storage_data_761 <= (fillup_transition == 1'b1) ? i_input_data[208 % IN_WIDTH] : ping_storage_data_761 ^ i_input_data[208 % IN_WIDTH];
                663 / IN_WIDTH: ping_storage_data_761 <= (fillup_transition == 1'b1) ? i_input_data[663 % IN_WIDTH] : ping_storage_data_761 ^ i_input_data[663 % IN_WIDTH];
                906 / IN_WIDTH: ping_storage_data_761 <= (fillup_transition == 1'b1) ? i_input_data[906 % IN_WIDTH] : ping_storage_data_761 ^ i_input_data[906 % IN_WIDTH];
                default: ping_storage_data_761 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_761;
                endcase
            end else begin
                case (input_count)
                174 / IN_WIDTH: pong_storage_data_761 <= (fillup_transition == 1'b1) ? i_input_data[174 % IN_WIDTH] : pong_storage_data_761 ^ i_input_data[174 % IN_WIDTH];
                208 / IN_WIDTH: pong_storage_data_761 <= (fillup_transition == 1'b1) ? i_input_data[208 % IN_WIDTH] : pong_storage_data_761 ^ i_input_data[208 % IN_WIDTH];
                663 / IN_WIDTH: pong_storage_data_761 <= (fillup_transition == 1'b1) ? i_input_data[663 % IN_WIDTH] : pong_storage_data_761 ^ i_input_data[663 % IN_WIDTH];
                906 / IN_WIDTH: pong_storage_data_761 <= (fillup_transition == 1'b1) ? i_input_data[906 % IN_WIDTH] : pong_storage_data_761 ^ i_input_data[906 % IN_WIDTH];
                default: pong_storage_data_761 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_761;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_761 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_761;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_761 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_761;
            end
        end
    end
end

logic ping_storage_data_762;
logic pong_storage_data_762;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_762 <= 1'b0;
        pong_storage_data_762 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                175 / IN_WIDTH: ping_storage_data_762 <= (fillup_transition == 1'b1) ? i_input_data[175 % IN_WIDTH] : ping_storage_data_762 ^ i_input_data[175 % IN_WIDTH];
                209 / IN_WIDTH: ping_storage_data_762 <= (fillup_transition == 1'b1) ? i_input_data[209 % IN_WIDTH] : ping_storage_data_762 ^ i_input_data[209 % IN_WIDTH];
                664 / IN_WIDTH: ping_storage_data_762 <= (fillup_transition == 1'b1) ? i_input_data[664 % IN_WIDTH] : ping_storage_data_762 ^ i_input_data[664 % IN_WIDTH];
                907 / IN_WIDTH: ping_storage_data_762 <= (fillup_transition == 1'b1) ? i_input_data[907 % IN_WIDTH] : ping_storage_data_762 ^ i_input_data[907 % IN_WIDTH];
                default: ping_storage_data_762 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_762;
                endcase
            end else begin
                case (input_count)
                175 / IN_WIDTH: pong_storage_data_762 <= (fillup_transition == 1'b1) ? i_input_data[175 % IN_WIDTH] : pong_storage_data_762 ^ i_input_data[175 % IN_WIDTH];
                209 / IN_WIDTH: pong_storage_data_762 <= (fillup_transition == 1'b1) ? i_input_data[209 % IN_WIDTH] : pong_storage_data_762 ^ i_input_data[209 % IN_WIDTH];
                664 / IN_WIDTH: pong_storage_data_762 <= (fillup_transition == 1'b1) ? i_input_data[664 % IN_WIDTH] : pong_storage_data_762 ^ i_input_data[664 % IN_WIDTH];
                907 / IN_WIDTH: pong_storage_data_762 <= (fillup_transition == 1'b1) ? i_input_data[907 % IN_WIDTH] : pong_storage_data_762 ^ i_input_data[907 % IN_WIDTH];
                default: pong_storage_data_762 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_762;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_762 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_762;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_762 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_762;
            end
        end
    end
end

logic ping_storage_data_763;
logic pong_storage_data_763;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_763 <= 1'b0;
        pong_storage_data_763 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                176 / IN_WIDTH: ping_storage_data_763 <= (fillup_transition == 1'b1) ? i_input_data[176 % IN_WIDTH] : ping_storage_data_763 ^ i_input_data[176 % IN_WIDTH];
                210 / IN_WIDTH: ping_storage_data_763 <= (fillup_transition == 1'b1) ? i_input_data[210 % IN_WIDTH] : ping_storage_data_763 ^ i_input_data[210 % IN_WIDTH];
                665 / IN_WIDTH: ping_storage_data_763 <= (fillup_transition == 1'b1) ? i_input_data[665 % IN_WIDTH] : ping_storage_data_763 ^ i_input_data[665 % IN_WIDTH];
                908 / IN_WIDTH: ping_storage_data_763 <= (fillup_transition == 1'b1) ? i_input_data[908 % IN_WIDTH] : ping_storage_data_763 ^ i_input_data[908 % IN_WIDTH];
                default: ping_storage_data_763 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_763;
                endcase
            end else begin
                case (input_count)
                176 / IN_WIDTH: pong_storage_data_763 <= (fillup_transition == 1'b1) ? i_input_data[176 % IN_WIDTH] : pong_storage_data_763 ^ i_input_data[176 % IN_WIDTH];
                210 / IN_WIDTH: pong_storage_data_763 <= (fillup_transition == 1'b1) ? i_input_data[210 % IN_WIDTH] : pong_storage_data_763 ^ i_input_data[210 % IN_WIDTH];
                665 / IN_WIDTH: pong_storage_data_763 <= (fillup_transition == 1'b1) ? i_input_data[665 % IN_WIDTH] : pong_storage_data_763 ^ i_input_data[665 % IN_WIDTH];
                908 / IN_WIDTH: pong_storage_data_763 <= (fillup_transition == 1'b1) ? i_input_data[908 % IN_WIDTH] : pong_storage_data_763 ^ i_input_data[908 % IN_WIDTH];
                default: pong_storage_data_763 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_763;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_763 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_763;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_763 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_763;
            end
        end
    end
end

logic ping_storage_data_764;
logic pong_storage_data_764;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_764 <= 1'b0;
        pong_storage_data_764 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                177 / IN_WIDTH: ping_storage_data_764 <= (fillup_transition == 1'b1) ? i_input_data[177 % IN_WIDTH] : ping_storage_data_764 ^ i_input_data[177 % IN_WIDTH];
                211 / IN_WIDTH: ping_storage_data_764 <= (fillup_transition == 1'b1) ? i_input_data[211 % IN_WIDTH] : ping_storage_data_764 ^ i_input_data[211 % IN_WIDTH];
                666 / IN_WIDTH: ping_storage_data_764 <= (fillup_transition == 1'b1) ? i_input_data[666 % IN_WIDTH] : ping_storage_data_764 ^ i_input_data[666 % IN_WIDTH];
                909 / IN_WIDTH: ping_storage_data_764 <= (fillup_transition == 1'b1) ? i_input_data[909 % IN_WIDTH] : ping_storage_data_764 ^ i_input_data[909 % IN_WIDTH];
                default: ping_storage_data_764 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_764;
                endcase
            end else begin
                case (input_count)
                177 / IN_WIDTH: pong_storage_data_764 <= (fillup_transition == 1'b1) ? i_input_data[177 % IN_WIDTH] : pong_storage_data_764 ^ i_input_data[177 % IN_WIDTH];
                211 / IN_WIDTH: pong_storage_data_764 <= (fillup_transition == 1'b1) ? i_input_data[211 % IN_WIDTH] : pong_storage_data_764 ^ i_input_data[211 % IN_WIDTH];
                666 / IN_WIDTH: pong_storage_data_764 <= (fillup_transition == 1'b1) ? i_input_data[666 % IN_WIDTH] : pong_storage_data_764 ^ i_input_data[666 % IN_WIDTH];
                909 / IN_WIDTH: pong_storage_data_764 <= (fillup_transition == 1'b1) ? i_input_data[909 % IN_WIDTH] : pong_storage_data_764 ^ i_input_data[909 % IN_WIDTH];
                default: pong_storage_data_764 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_764;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_764 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_764;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_764 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_764;
            end
        end
    end
end

logic ping_storage_data_765;
logic pong_storage_data_765;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_765 <= 1'b0;
        pong_storage_data_765 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                178 / IN_WIDTH: ping_storage_data_765 <= (fillup_transition == 1'b1) ? i_input_data[178 % IN_WIDTH] : ping_storage_data_765 ^ i_input_data[178 % IN_WIDTH];
                212 / IN_WIDTH: ping_storage_data_765 <= (fillup_transition == 1'b1) ? i_input_data[212 % IN_WIDTH] : ping_storage_data_765 ^ i_input_data[212 % IN_WIDTH];
                667 / IN_WIDTH: ping_storage_data_765 <= (fillup_transition == 1'b1) ? i_input_data[667 % IN_WIDTH] : ping_storage_data_765 ^ i_input_data[667 % IN_WIDTH];
                910 / IN_WIDTH: ping_storage_data_765 <= (fillup_transition == 1'b1) ? i_input_data[910 % IN_WIDTH] : ping_storage_data_765 ^ i_input_data[910 % IN_WIDTH];
                default: ping_storage_data_765 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_765;
                endcase
            end else begin
                case (input_count)
                178 / IN_WIDTH: pong_storage_data_765 <= (fillup_transition == 1'b1) ? i_input_data[178 % IN_WIDTH] : pong_storage_data_765 ^ i_input_data[178 % IN_WIDTH];
                212 / IN_WIDTH: pong_storage_data_765 <= (fillup_transition == 1'b1) ? i_input_data[212 % IN_WIDTH] : pong_storage_data_765 ^ i_input_data[212 % IN_WIDTH];
                667 / IN_WIDTH: pong_storage_data_765 <= (fillup_transition == 1'b1) ? i_input_data[667 % IN_WIDTH] : pong_storage_data_765 ^ i_input_data[667 % IN_WIDTH];
                910 / IN_WIDTH: pong_storage_data_765 <= (fillup_transition == 1'b1) ? i_input_data[910 % IN_WIDTH] : pong_storage_data_765 ^ i_input_data[910 % IN_WIDTH];
                default: pong_storage_data_765 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_765;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_765 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_765;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_765 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_765;
            end
        end
    end
end

logic ping_storage_data_766;
logic pong_storage_data_766;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_766 <= 1'b0;
        pong_storage_data_766 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                179 / IN_WIDTH: ping_storage_data_766 <= (fillup_transition == 1'b1) ? i_input_data[179 % IN_WIDTH] : ping_storage_data_766 ^ i_input_data[179 % IN_WIDTH];
                213 / IN_WIDTH: ping_storage_data_766 <= (fillup_transition == 1'b1) ? i_input_data[213 % IN_WIDTH] : ping_storage_data_766 ^ i_input_data[213 % IN_WIDTH];
                668 / IN_WIDTH: ping_storage_data_766 <= (fillup_transition == 1'b1) ? i_input_data[668 % IN_WIDTH] : ping_storage_data_766 ^ i_input_data[668 % IN_WIDTH];
                911 / IN_WIDTH: ping_storage_data_766 <= (fillup_transition == 1'b1) ? i_input_data[911 % IN_WIDTH] : ping_storage_data_766 ^ i_input_data[911 % IN_WIDTH];
                default: ping_storage_data_766 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_766;
                endcase
            end else begin
                case (input_count)
                179 / IN_WIDTH: pong_storage_data_766 <= (fillup_transition == 1'b1) ? i_input_data[179 % IN_WIDTH] : pong_storage_data_766 ^ i_input_data[179 % IN_WIDTH];
                213 / IN_WIDTH: pong_storage_data_766 <= (fillup_transition == 1'b1) ? i_input_data[213 % IN_WIDTH] : pong_storage_data_766 ^ i_input_data[213 % IN_WIDTH];
                668 / IN_WIDTH: pong_storage_data_766 <= (fillup_transition == 1'b1) ? i_input_data[668 % IN_WIDTH] : pong_storage_data_766 ^ i_input_data[668 % IN_WIDTH];
                911 / IN_WIDTH: pong_storage_data_766 <= (fillup_transition == 1'b1) ? i_input_data[911 % IN_WIDTH] : pong_storage_data_766 ^ i_input_data[911 % IN_WIDTH];
                default: pong_storage_data_766 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_766;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_766 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_766;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_766 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_766;
            end
        end
    end
end

logic ping_storage_data_767;
logic pong_storage_data_767;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_767 <= 1'b0;
        pong_storage_data_767 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                180 / IN_WIDTH: ping_storage_data_767 <= (fillup_transition == 1'b1) ? i_input_data[180 % IN_WIDTH] : ping_storage_data_767 ^ i_input_data[180 % IN_WIDTH];
                214 / IN_WIDTH: ping_storage_data_767 <= (fillup_transition == 1'b1) ? i_input_data[214 % IN_WIDTH] : ping_storage_data_767 ^ i_input_data[214 % IN_WIDTH];
                669 / IN_WIDTH: ping_storage_data_767 <= (fillup_transition == 1'b1) ? i_input_data[669 % IN_WIDTH] : ping_storage_data_767 ^ i_input_data[669 % IN_WIDTH];
                912 / IN_WIDTH: ping_storage_data_767 <= (fillup_transition == 1'b1) ? i_input_data[912 % IN_WIDTH] : ping_storage_data_767 ^ i_input_data[912 % IN_WIDTH];
                default: ping_storage_data_767 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_767;
                endcase
            end else begin
                case (input_count)
                180 / IN_WIDTH: pong_storage_data_767 <= (fillup_transition == 1'b1) ? i_input_data[180 % IN_WIDTH] : pong_storage_data_767 ^ i_input_data[180 % IN_WIDTH];
                214 / IN_WIDTH: pong_storage_data_767 <= (fillup_transition == 1'b1) ? i_input_data[214 % IN_WIDTH] : pong_storage_data_767 ^ i_input_data[214 % IN_WIDTH];
                669 / IN_WIDTH: pong_storage_data_767 <= (fillup_transition == 1'b1) ? i_input_data[669 % IN_WIDTH] : pong_storage_data_767 ^ i_input_data[669 % IN_WIDTH];
                912 / IN_WIDTH: pong_storage_data_767 <= (fillup_transition == 1'b1) ? i_input_data[912 % IN_WIDTH] : pong_storage_data_767 ^ i_input_data[912 % IN_WIDTH];
                default: pong_storage_data_767 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_767;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_767 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_767;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_767 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_767;
            end
        end
    end
end

logic ping_storage_data_768;
logic pong_storage_data_768;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_768 <= 1'b0;
        pong_storage_data_768 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                84 / IN_WIDTH: ping_storage_data_768 <= (fillup_transition == 1'b1) ? i_input_data[84 % IN_WIDTH] : ping_storage_data_768 ^ i_input_data[84 % IN_WIDTH];
                397 / IN_WIDTH: ping_storage_data_768 <= (fillup_transition == 1'b1) ? i_input_data[397 % IN_WIDTH] : ping_storage_data_768 ^ i_input_data[397 % IN_WIDTH];
                552 / IN_WIDTH: ping_storage_data_768 <= (fillup_transition == 1'b1) ? i_input_data[552 % IN_WIDTH] : ping_storage_data_768 ^ i_input_data[552 % IN_WIDTH];
                725 / IN_WIDTH: ping_storage_data_768 <= (fillup_transition == 1'b1) ? i_input_data[725 % IN_WIDTH] : ping_storage_data_768 ^ i_input_data[725 % IN_WIDTH];
                1101 / IN_WIDTH: ping_storage_data_768 <= (fillup_transition == 1'b1) ? i_input_data[1101 % IN_WIDTH] : ping_storage_data_768 ^ i_input_data[1101 % IN_WIDTH];
                default: ping_storage_data_768 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_768;
                endcase
            end else begin
                case (input_count)
                84 / IN_WIDTH: pong_storage_data_768 <= (fillup_transition == 1'b1) ? i_input_data[84 % IN_WIDTH] : pong_storage_data_768 ^ i_input_data[84 % IN_WIDTH];
                397 / IN_WIDTH: pong_storage_data_768 <= (fillup_transition == 1'b1) ? i_input_data[397 % IN_WIDTH] : pong_storage_data_768 ^ i_input_data[397 % IN_WIDTH];
                552 / IN_WIDTH: pong_storage_data_768 <= (fillup_transition == 1'b1) ? i_input_data[552 % IN_WIDTH] : pong_storage_data_768 ^ i_input_data[552 % IN_WIDTH];
                725 / IN_WIDTH: pong_storage_data_768 <= (fillup_transition == 1'b1) ? i_input_data[725 % IN_WIDTH] : pong_storage_data_768 ^ i_input_data[725 % IN_WIDTH];
                1101 / IN_WIDTH: pong_storage_data_768 <= (fillup_transition == 1'b1) ? i_input_data[1101 % IN_WIDTH] : pong_storage_data_768 ^ i_input_data[1101 % IN_WIDTH];
                default: pong_storage_data_768 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_768;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_768 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_768;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_768 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_768;
            end
        end
    end
end

logic ping_storage_data_769;
logic pong_storage_data_769;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_769 <= 1'b0;
        pong_storage_data_769 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                85 / IN_WIDTH: ping_storage_data_769 <= (fillup_transition == 1'b1) ? i_input_data[85 % IN_WIDTH] : ping_storage_data_769 ^ i_input_data[85 % IN_WIDTH];
                398 / IN_WIDTH: ping_storage_data_769 <= (fillup_transition == 1'b1) ? i_input_data[398 % IN_WIDTH] : ping_storage_data_769 ^ i_input_data[398 % IN_WIDTH];
                553 / IN_WIDTH: ping_storage_data_769 <= (fillup_transition == 1'b1) ? i_input_data[553 % IN_WIDTH] : ping_storage_data_769 ^ i_input_data[553 % IN_WIDTH];
                726 / IN_WIDTH: ping_storage_data_769 <= (fillup_transition == 1'b1) ? i_input_data[726 % IN_WIDTH] : ping_storage_data_769 ^ i_input_data[726 % IN_WIDTH];
                1102 / IN_WIDTH: ping_storage_data_769 <= (fillup_transition == 1'b1) ? i_input_data[1102 % IN_WIDTH] : ping_storage_data_769 ^ i_input_data[1102 % IN_WIDTH];
                default: ping_storage_data_769 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_769;
                endcase
            end else begin
                case (input_count)
                85 / IN_WIDTH: pong_storage_data_769 <= (fillup_transition == 1'b1) ? i_input_data[85 % IN_WIDTH] : pong_storage_data_769 ^ i_input_data[85 % IN_WIDTH];
                398 / IN_WIDTH: pong_storage_data_769 <= (fillup_transition == 1'b1) ? i_input_data[398 % IN_WIDTH] : pong_storage_data_769 ^ i_input_data[398 % IN_WIDTH];
                553 / IN_WIDTH: pong_storage_data_769 <= (fillup_transition == 1'b1) ? i_input_data[553 % IN_WIDTH] : pong_storage_data_769 ^ i_input_data[553 % IN_WIDTH];
                726 / IN_WIDTH: pong_storage_data_769 <= (fillup_transition == 1'b1) ? i_input_data[726 % IN_WIDTH] : pong_storage_data_769 ^ i_input_data[726 % IN_WIDTH];
                1102 / IN_WIDTH: pong_storage_data_769 <= (fillup_transition == 1'b1) ? i_input_data[1102 % IN_WIDTH] : pong_storage_data_769 ^ i_input_data[1102 % IN_WIDTH];
                default: pong_storage_data_769 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_769;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_769 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_769;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_769 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_769;
            end
        end
    end
end

logic ping_storage_data_770;
logic pong_storage_data_770;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_770 <= 1'b0;
        pong_storage_data_770 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                86 / IN_WIDTH: ping_storage_data_770 <= (fillup_transition == 1'b1) ? i_input_data[86 % IN_WIDTH] : ping_storage_data_770 ^ i_input_data[86 % IN_WIDTH];
                399 / IN_WIDTH: ping_storage_data_770 <= (fillup_transition == 1'b1) ? i_input_data[399 % IN_WIDTH] : ping_storage_data_770 ^ i_input_data[399 % IN_WIDTH];
                554 / IN_WIDTH: ping_storage_data_770 <= (fillup_transition == 1'b1) ? i_input_data[554 % IN_WIDTH] : ping_storage_data_770 ^ i_input_data[554 % IN_WIDTH];
                727 / IN_WIDTH: ping_storage_data_770 <= (fillup_transition == 1'b1) ? i_input_data[727 % IN_WIDTH] : ping_storage_data_770 ^ i_input_data[727 % IN_WIDTH];
                1103 / IN_WIDTH: ping_storage_data_770 <= (fillup_transition == 1'b1) ? i_input_data[1103 % IN_WIDTH] : ping_storage_data_770 ^ i_input_data[1103 % IN_WIDTH];
                default: ping_storage_data_770 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_770;
                endcase
            end else begin
                case (input_count)
                86 / IN_WIDTH: pong_storage_data_770 <= (fillup_transition == 1'b1) ? i_input_data[86 % IN_WIDTH] : pong_storage_data_770 ^ i_input_data[86 % IN_WIDTH];
                399 / IN_WIDTH: pong_storage_data_770 <= (fillup_transition == 1'b1) ? i_input_data[399 % IN_WIDTH] : pong_storage_data_770 ^ i_input_data[399 % IN_WIDTH];
                554 / IN_WIDTH: pong_storage_data_770 <= (fillup_transition == 1'b1) ? i_input_data[554 % IN_WIDTH] : pong_storage_data_770 ^ i_input_data[554 % IN_WIDTH];
                727 / IN_WIDTH: pong_storage_data_770 <= (fillup_transition == 1'b1) ? i_input_data[727 % IN_WIDTH] : pong_storage_data_770 ^ i_input_data[727 % IN_WIDTH];
                1103 / IN_WIDTH: pong_storage_data_770 <= (fillup_transition == 1'b1) ? i_input_data[1103 % IN_WIDTH] : pong_storage_data_770 ^ i_input_data[1103 % IN_WIDTH];
                default: pong_storage_data_770 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_770;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_770 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_770;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_770 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_770;
            end
        end
    end
end

logic ping_storage_data_771;
logic pong_storage_data_771;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_771 <= 1'b0;
        pong_storage_data_771 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                87 / IN_WIDTH: ping_storage_data_771 <= (fillup_transition == 1'b1) ? i_input_data[87 % IN_WIDTH] : ping_storage_data_771 ^ i_input_data[87 % IN_WIDTH];
                400 / IN_WIDTH: ping_storage_data_771 <= (fillup_transition == 1'b1) ? i_input_data[400 % IN_WIDTH] : ping_storage_data_771 ^ i_input_data[400 % IN_WIDTH];
                555 / IN_WIDTH: ping_storage_data_771 <= (fillup_transition == 1'b1) ? i_input_data[555 % IN_WIDTH] : ping_storage_data_771 ^ i_input_data[555 % IN_WIDTH];
                728 / IN_WIDTH: ping_storage_data_771 <= (fillup_transition == 1'b1) ? i_input_data[728 % IN_WIDTH] : ping_storage_data_771 ^ i_input_data[728 % IN_WIDTH];
                1104 / IN_WIDTH: ping_storage_data_771 <= (fillup_transition == 1'b1) ? i_input_data[1104 % IN_WIDTH] : ping_storage_data_771 ^ i_input_data[1104 % IN_WIDTH];
                default: ping_storage_data_771 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_771;
                endcase
            end else begin
                case (input_count)
                87 / IN_WIDTH: pong_storage_data_771 <= (fillup_transition == 1'b1) ? i_input_data[87 % IN_WIDTH] : pong_storage_data_771 ^ i_input_data[87 % IN_WIDTH];
                400 / IN_WIDTH: pong_storage_data_771 <= (fillup_transition == 1'b1) ? i_input_data[400 % IN_WIDTH] : pong_storage_data_771 ^ i_input_data[400 % IN_WIDTH];
                555 / IN_WIDTH: pong_storage_data_771 <= (fillup_transition == 1'b1) ? i_input_data[555 % IN_WIDTH] : pong_storage_data_771 ^ i_input_data[555 % IN_WIDTH];
                728 / IN_WIDTH: pong_storage_data_771 <= (fillup_transition == 1'b1) ? i_input_data[728 % IN_WIDTH] : pong_storage_data_771 ^ i_input_data[728 % IN_WIDTH];
                1104 / IN_WIDTH: pong_storage_data_771 <= (fillup_transition == 1'b1) ? i_input_data[1104 % IN_WIDTH] : pong_storage_data_771 ^ i_input_data[1104 % IN_WIDTH];
                default: pong_storage_data_771 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_771;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_771 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_771;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_771 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_771;
            end
        end
    end
end

logic ping_storage_data_772;
logic pong_storage_data_772;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_772 <= 1'b0;
        pong_storage_data_772 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                88 / IN_WIDTH: ping_storage_data_772 <= (fillup_transition == 1'b1) ? i_input_data[88 % IN_WIDTH] : ping_storage_data_772 ^ i_input_data[88 % IN_WIDTH];
                401 / IN_WIDTH: ping_storage_data_772 <= (fillup_transition == 1'b1) ? i_input_data[401 % IN_WIDTH] : ping_storage_data_772 ^ i_input_data[401 % IN_WIDTH];
                556 / IN_WIDTH: ping_storage_data_772 <= (fillup_transition == 1'b1) ? i_input_data[556 % IN_WIDTH] : ping_storage_data_772 ^ i_input_data[556 % IN_WIDTH];
                729 / IN_WIDTH: ping_storage_data_772 <= (fillup_transition == 1'b1) ? i_input_data[729 % IN_WIDTH] : ping_storage_data_772 ^ i_input_data[729 % IN_WIDTH];
                1105 / IN_WIDTH: ping_storage_data_772 <= (fillup_transition == 1'b1) ? i_input_data[1105 % IN_WIDTH] : ping_storage_data_772 ^ i_input_data[1105 % IN_WIDTH];
                default: ping_storage_data_772 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_772;
                endcase
            end else begin
                case (input_count)
                88 / IN_WIDTH: pong_storage_data_772 <= (fillup_transition == 1'b1) ? i_input_data[88 % IN_WIDTH] : pong_storage_data_772 ^ i_input_data[88 % IN_WIDTH];
                401 / IN_WIDTH: pong_storage_data_772 <= (fillup_transition == 1'b1) ? i_input_data[401 % IN_WIDTH] : pong_storage_data_772 ^ i_input_data[401 % IN_WIDTH];
                556 / IN_WIDTH: pong_storage_data_772 <= (fillup_transition == 1'b1) ? i_input_data[556 % IN_WIDTH] : pong_storage_data_772 ^ i_input_data[556 % IN_WIDTH];
                729 / IN_WIDTH: pong_storage_data_772 <= (fillup_transition == 1'b1) ? i_input_data[729 % IN_WIDTH] : pong_storage_data_772 ^ i_input_data[729 % IN_WIDTH];
                1105 / IN_WIDTH: pong_storage_data_772 <= (fillup_transition == 1'b1) ? i_input_data[1105 % IN_WIDTH] : pong_storage_data_772 ^ i_input_data[1105 % IN_WIDTH];
                default: pong_storage_data_772 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_772;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_772 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_772;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_772 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_772;
            end
        end
    end
end

logic ping_storage_data_773;
logic pong_storage_data_773;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_773 <= 1'b0;
        pong_storage_data_773 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                89 / IN_WIDTH: ping_storage_data_773 <= (fillup_transition == 1'b1) ? i_input_data[89 % IN_WIDTH] : ping_storage_data_773 ^ i_input_data[89 % IN_WIDTH];
                402 / IN_WIDTH: ping_storage_data_773 <= (fillup_transition == 1'b1) ? i_input_data[402 % IN_WIDTH] : ping_storage_data_773 ^ i_input_data[402 % IN_WIDTH];
                557 / IN_WIDTH: ping_storage_data_773 <= (fillup_transition == 1'b1) ? i_input_data[557 % IN_WIDTH] : ping_storage_data_773 ^ i_input_data[557 % IN_WIDTH];
                730 / IN_WIDTH: ping_storage_data_773 <= (fillup_transition == 1'b1) ? i_input_data[730 % IN_WIDTH] : ping_storage_data_773 ^ i_input_data[730 % IN_WIDTH];
                1106 / IN_WIDTH: ping_storage_data_773 <= (fillup_transition == 1'b1) ? i_input_data[1106 % IN_WIDTH] : ping_storage_data_773 ^ i_input_data[1106 % IN_WIDTH];
                default: ping_storage_data_773 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_773;
                endcase
            end else begin
                case (input_count)
                89 / IN_WIDTH: pong_storage_data_773 <= (fillup_transition == 1'b1) ? i_input_data[89 % IN_WIDTH] : pong_storage_data_773 ^ i_input_data[89 % IN_WIDTH];
                402 / IN_WIDTH: pong_storage_data_773 <= (fillup_transition == 1'b1) ? i_input_data[402 % IN_WIDTH] : pong_storage_data_773 ^ i_input_data[402 % IN_WIDTH];
                557 / IN_WIDTH: pong_storage_data_773 <= (fillup_transition == 1'b1) ? i_input_data[557 % IN_WIDTH] : pong_storage_data_773 ^ i_input_data[557 % IN_WIDTH];
                730 / IN_WIDTH: pong_storage_data_773 <= (fillup_transition == 1'b1) ? i_input_data[730 % IN_WIDTH] : pong_storage_data_773 ^ i_input_data[730 % IN_WIDTH];
                1106 / IN_WIDTH: pong_storage_data_773 <= (fillup_transition == 1'b1) ? i_input_data[1106 % IN_WIDTH] : pong_storage_data_773 ^ i_input_data[1106 % IN_WIDTH];
                default: pong_storage_data_773 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_773;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_773 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_773;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_773 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_773;
            end
        end
    end
end

logic ping_storage_data_774;
logic pong_storage_data_774;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_774 <= 1'b0;
        pong_storage_data_774 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                90 / IN_WIDTH: ping_storage_data_774 <= (fillup_transition == 1'b1) ? i_input_data[90 % IN_WIDTH] : ping_storage_data_774 ^ i_input_data[90 % IN_WIDTH];
                403 / IN_WIDTH: ping_storage_data_774 <= (fillup_transition == 1'b1) ? i_input_data[403 % IN_WIDTH] : ping_storage_data_774 ^ i_input_data[403 % IN_WIDTH];
                558 / IN_WIDTH: ping_storage_data_774 <= (fillup_transition == 1'b1) ? i_input_data[558 % IN_WIDTH] : ping_storage_data_774 ^ i_input_data[558 % IN_WIDTH];
                731 / IN_WIDTH: ping_storage_data_774 <= (fillup_transition == 1'b1) ? i_input_data[731 % IN_WIDTH] : ping_storage_data_774 ^ i_input_data[731 % IN_WIDTH];
                1107 / IN_WIDTH: ping_storage_data_774 <= (fillup_transition == 1'b1) ? i_input_data[1107 % IN_WIDTH] : ping_storage_data_774 ^ i_input_data[1107 % IN_WIDTH];
                default: ping_storage_data_774 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_774;
                endcase
            end else begin
                case (input_count)
                90 / IN_WIDTH: pong_storage_data_774 <= (fillup_transition == 1'b1) ? i_input_data[90 % IN_WIDTH] : pong_storage_data_774 ^ i_input_data[90 % IN_WIDTH];
                403 / IN_WIDTH: pong_storage_data_774 <= (fillup_transition == 1'b1) ? i_input_data[403 % IN_WIDTH] : pong_storage_data_774 ^ i_input_data[403 % IN_WIDTH];
                558 / IN_WIDTH: pong_storage_data_774 <= (fillup_transition == 1'b1) ? i_input_data[558 % IN_WIDTH] : pong_storage_data_774 ^ i_input_data[558 % IN_WIDTH];
                731 / IN_WIDTH: pong_storage_data_774 <= (fillup_transition == 1'b1) ? i_input_data[731 % IN_WIDTH] : pong_storage_data_774 ^ i_input_data[731 % IN_WIDTH];
                1107 / IN_WIDTH: pong_storage_data_774 <= (fillup_transition == 1'b1) ? i_input_data[1107 % IN_WIDTH] : pong_storage_data_774 ^ i_input_data[1107 % IN_WIDTH];
                default: pong_storage_data_774 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_774;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_774 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_774;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_774 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_774;
            end
        end
    end
end

logic ping_storage_data_775;
logic pong_storage_data_775;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_775 <= 1'b0;
        pong_storage_data_775 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                91 / IN_WIDTH: ping_storage_data_775 <= (fillup_transition == 1'b1) ? i_input_data[91 % IN_WIDTH] : ping_storage_data_775 ^ i_input_data[91 % IN_WIDTH];
                404 / IN_WIDTH: ping_storage_data_775 <= (fillup_transition == 1'b1) ? i_input_data[404 % IN_WIDTH] : ping_storage_data_775 ^ i_input_data[404 % IN_WIDTH];
                559 / IN_WIDTH: ping_storage_data_775 <= (fillup_transition == 1'b1) ? i_input_data[559 % IN_WIDTH] : ping_storage_data_775 ^ i_input_data[559 % IN_WIDTH];
                732 / IN_WIDTH: ping_storage_data_775 <= (fillup_transition == 1'b1) ? i_input_data[732 % IN_WIDTH] : ping_storage_data_775 ^ i_input_data[732 % IN_WIDTH];
                1108 / IN_WIDTH: ping_storage_data_775 <= (fillup_transition == 1'b1) ? i_input_data[1108 % IN_WIDTH] : ping_storage_data_775 ^ i_input_data[1108 % IN_WIDTH];
                default: ping_storage_data_775 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_775;
                endcase
            end else begin
                case (input_count)
                91 / IN_WIDTH: pong_storage_data_775 <= (fillup_transition == 1'b1) ? i_input_data[91 % IN_WIDTH] : pong_storage_data_775 ^ i_input_data[91 % IN_WIDTH];
                404 / IN_WIDTH: pong_storage_data_775 <= (fillup_transition == 1'b1) ? i_input_data[404 % IN_WIDTH] : pong_storage_data_775 ^ i_input_data[404 % IN_WIDTH];
                559 / IN_WIDTH: pong_storage_data_775 <= (fillup_transition == 1'b1) ? i_input_data[559 % IN_WIDTH] : pong_storage_data_775 ^ i_input_data[559 % IN_WIDTH];
                732 / IN_WIDTH: pong_storage_data_775 <= (fillup_transition == 1'b1) ? i_input_data[732 % IN_WIDTH] : pong_storage_data_775 ^ i_input_data[732 % IN_WIDTH];
                1108 / IN_WIDTH: pong_storage_data_775 <= (fillup_transition == 1'b1) ? i_input_data[1108 % IN_WIDTH] : pong_storage_data_775 ^ i_input_data[1108 % IN_WIDTH];
                default: pong_storage_data_775 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_775;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_775 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_775;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_775 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_775;
            end
        end
    end
end

logic ping_storage_data_776;
logic pong_storage_data_776;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_776 <= 1'b0;
        pong_storage_data_776 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                92 / IN_WIDTH: ping_storage_data_776 <= (fillup_transition == 1'b1) ? i_input_data[92 % IN_WIDTH] : ping_storage_data_776 ^ i_input_data[92 % IN_WIDTH];
                405 / IN_WIDTH: ping_storage_data_776 <= (fillup_transition == 1'b1) ? i_input_data[405 % IN_WIDTH] : ping_storage_data_776 ^ i_input_data[405 % IN_WIDTH];
                560 / IN_WIDTH: ping_storage_data_776 <= (fillup_transition == 1'b1) ? i_input_data[560 % IN_WIDTH] : ping_storage_data_776 ^ i_input_data[560 % IN_WIDTH];
                733 / IN_WIDTH: ping_storage_data_776 <= (fillup_transition == 1'b1) ? i_input_data[733 % IN_WIDTH] : ping_storage_data_776 ^ i_input_data[733 % IN_WIDTH];
                1109 / IN_WIDTH: ping_storage_data_776 <= (fillup_transition == 1'b1) ? i_input_data[1109 % IN_WIDTH] : ping_storage_data_776 ^ i_input_data[1109 % IN_WIDTH];
                default: ping_storage_data_776 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_776;
                endcase
            end else begin
                case (input_count)
                92 / IN_WIDTH: pong_storage_data_776 <= (fillup_transition == 1'b1) ? i_input_data[92 % IN_WIDTH] : pong_storage_data_776 ^ i_input_data[92 % IN_WIDTH];
                405 / IN_WIDTH: pong_storage_data_776 <= (fillup_transition == 1'b1) ? i_input_data[405 % IN_WIDTH] : pong_storage_data_776 ^ i_input_data[405 % IN_WIDTH];
                560 / IN_WIDTH: pong_storage_data_776 <= (fillup_transition == 1'b1) ? i_input_data[560 % IN_WIDTH] : pong_storage_data_776 ^ i_input_data[560 % IN_WIDTH];
                733 / IN_WIDTH: pong_storage_data_776 <= (fillup_transition == 1'b1) ? i_input_data[733 % IN_WIDTH] : pong_storage_data_776 ^ i_input_data[733 % IN_WIDTH];
                1109 / IN_WIDTH: pong_storage_data_776 <= (fillup_transition == 1'b1) ? i_input_data[1109 % IN_WIDTH] : pong_storage_data_776 ^ i_input_data[1109 % IN_WIDTH];
                default: pong_storage_data_776 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_776;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_776 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_776;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_776 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_776;
            end
        end
    end
end

logic ping_storage_data_777;
logic pong_storage_data_777;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_777 <= 1'b0;
        pong_storage_data_777 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                93 / IN_WIDTH: ping_storage_data_777 <= (fillup_transition == 1'b1) ? i_input_data[93 % IN_WIDTH] : ping_storage_data_777 ^ i_input_data[93 % IN_WIDTH];
                406 / IN_WIDTH: ping_storage_data_777 <= (fillup_transition == 1'b1) ? i_input_data[406 % IN_WIDTH] : ping_storage_data_777 ^ i_input_data[406 % IN_WIDTH];
                561 / IN_WIDTH: ping_storage_data_777 <= (fillup_transition == 1'b1) ? i_input_data[561 % IN_WIDTH] : ping_storage_data_777 ^ i_input_data[561 % IN_WIDTH];
                734 / IN_WIDTH: ping_storage_data_777 <= (fillup_transition == 1'b1) ? i_input_data[734 % IN_WIDTH] : ping_storage_data_777 ^ i_input_data[734 % IN_WIDTH];
                1110 / IN_WIDTH: ping_storage_data_777 <= (fillup_transition == 1'b1) ? i_input_data[1110 % IN_WIDTH] : ping_storage_data_777 ^ i_input_data[1110 % IN_WIDTH];
                default: ping_storage_data_777 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_777;
                endcase
            end else begin
                case (input_count)
                93 / IN_WIDTH: pong_storage_data_777 <= (fillup_transition == 1'b1) ? i_input_data[93 % IN_WIDTH] : pong_storage_data_777 ^ i_input_data[93 % IN_WIDTH];
                406 / IN_WIDTH: pong_storage_data_777 <= (fillup_transition == 1'b1) ? i_input_data[406 % IN_WIDTH] : pong_storage_data_777 ^ i_input_data[406 % IN_WIDTH];
                561 / IN_WIDTH: pong_storage_data_777 <= (fillup_transition == 1'b1) ? i_input_data[561 % IN_WIDTH] : pong_storage_data_777 ^ i_input_data[561 % IN_WIDTH];
                734 / IN_WIDTH: pong_storage_data_777 <= (fillup_transition == 1'b1) ? i_input_data[734 % IN_WIDTH] : pong_storage_data_777 ^ i_input_data[734 % IN_WIDTH];
                1110 / IN_WIDTH: pong_storage_data_777 <= (fillup_transition == 1'b1) ? i_input_data[1110 % IN_WIDTH] : pong_storage_data_777 ^ i_input_data[1110 % IN_WIDTH];
                default: pong_storage_data_777 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_777;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_777 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_777;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_777 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_777;
            end
        end
    end
end

logic ping_storage_data_778;
logic pong_storage_data_778;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_778 <= 1'b0;
        pong_storage_data_778 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                94 / IN_WIDTH: ping_storage_data_778 <= (fillup_transition == 1'b1) ? i_input_data[94 % IN_WIDTH] : ping_storage_data_778 ^ i_input_data[94 % IN_WIDTH];
                407 / IN_WIDTH: ping_storage_data_778 <= (fillup_transition == 1'b1) ? i_input_data[407 % IN_WIDTH] : ping_storage_data_778 ^ i_input_data[407 % IN_WIDTH];
                562 / IN_WIDTH: ping_storage_data_778 <= (fillup_transition == 1'b1) ? i_input_data[562 % IN_WIDTH] : ping_storage_data_778 ^ i_input_data[562 % IN_WIDTH];
                735 / IN_WIDTH: ping_storage_data_778 <= (fillup_transition == 1'b1) ? i_input_data[735 % IN_WIDTH] : ping_storage_data_778 ^ i_input_data[735 % IN_WIDTH];
                1111 / IN_WIDTH: ping_storage_data_778 <= (fillup_transition == 1'b1) ? i_input_data[1111 % IN_WIDTH] : ping_storage_data_778 ^ i_input_data[1111 % IN_WIDTH];
                default: ping_storage_data_778 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_778;
                endcase
            end else begin
                case (input_count)
                94 / IN_WIDTH: pong_storage_data_778 <= (fillup_transition == 1'b1) ? i_input_data[94 % IN_WIDTH] : pong_storage_data_778 ^ i_input_data[94 % IN_WIDTH];
                407 / IN_WIDTH: pong_storage_data_778 <= (fillup_transition == 1'b1) ? i_input_data[407 % IN_WIDTH] : pong_storage_data_778 ^ i_input_data[407 % IN_WIDTH];
                562 / IN_WIDTH: pong_storage_data_778 <= (fillup_transition == 1'b1) ? i_input_data[562 % IN_WIDTH] : pong_storage_data_778 ^ i_input_data[562 % IN_WIDTH];
                735 / IN_WIDTH: pong_storage_data_778 <= (fillup_transition == 1'b1) ? i_input_data[735 % IN_WIDTH] : pong_storage_data_778 ^ i_input_data[735 % IN_WIDTH];
                1111 / IN_WIDTH: pong_storage_data_778 <= (fillup_transition == 1'b1) ? i_input_data[1111 % IN_WIDTH] : pong_storage_data_778 ^ i_input_data[1111 % IN_WIDTH];
                default: pong_storage_data_778 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_778;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_778 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_778;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_778 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_778;
            end
        end
    end
end

logic ping_storage_data_779;
logic pong_storage_data_779;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_779 <= 1'b0;
        pong_storage_data_779 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                95 / IN_WIDTH: ping_storage_data_779 <= (fillup_transition == 1'b1) ? i_input_data[95 % IN_WIDTH] : ping_storage_data_779 ^ i_input_data[95 % IN_WIDTH];
                408 / IN_WIDTH: ping_storage_data_779 <= (fillup_transition == 1'b1) ? i_input_data[408 % IN_WIDTH] : ping_storage_data_779 ^ i_input_data[408 % IN_WIDTH];
                563 / IN_WIDTH: ping_storage_data_779 <= (fillup_transition == 1'b1) ? i_input_data[563 % IN_WIDTH] : ping_storage_data_779 ^ i_input_data[563 % IN_WIDTH];
                736 / IN_WIDTH: ping_storage_data_779 <= (fillup_transition == 1'b1) ? i_input_data[736 % IN_WIDTH] : ping_storage_data_779 ^ i_input_data[736 % IN_WIDTH];
                1112 / IN_WIDTH: ping_storage_data_779 <= (fillup_transition == 1'b1) ? i_input_data[1112 % IN_WIDTH] : ping_storage_data_779 ^ i_input_data[1112 % IN_WIDTH];
                default: ping_storage_data_779 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_779;
                endcase
            end else begin
                case (input_count)
                95 / IN_WIDTH: pong_storage_data_779 <= (fillup_transition == 1'b1) ? i_input_data[95 % IN_WIDTH] : pong_storage_data_779 ^ i_input_data[95 % IN_WIDTH];
                408 / IN_WIDTH: pong_storage_data_779 <= (fillup_transition == 1'b1) ? i_input_data[408 % IN_WIDTH] : pong_storage_data_779 ^ i_input_data[408 % IN_WIDTH];
                563 / IN_WIDTH: pong_storage_data_779 <= (fillup_transition == 1'b1) ? i_input_data[563 % IN_WIDTH] : pong_storage_data_779 ^ i_input_data[563 % IN_WIDTH];
                736 / IN_WIDTH: pong_storage_data_779 <= (fillup_transition == 1'b1) ? i_input_data[736 % IN_WIDTH] : pong_storage_data_779 ^ i_input_data[736 % IN_WIDTH];
                1112 / IN_WIDTH: pong_storage_data_779 <= (fillup_transition == 1'b1) ? i_input_data[1112 % IN_WIDTH] : pong_storage_data_779 ^ i_input_data[1112 % IN_WIDTH];
                default: pong_storage_data_779 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_779;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_779 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_779;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_779 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_779;
            end
        end
    end
end

logic ping_storage_data_780;
logic pong_storage_data_780;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_780 <= 1'b0;
        pong_storage_data_780 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                0 / IN_WIDTH: ping_storage_data_780 <= (fillup_transition == 1'b1) ? i_input_data[0 % IN_WIDTH] : ping_storage_data_780 ^ i_input_data[0 % IN_WIDTH];
                409 / IN_WIDTH: ping_storage_data_780 <= (fillup_transition == 1'b1) ? i_input_data[409 % IN_WIDTH] : ping_storage_data_780 ^ i_input_data[409 % IN_WIDTH];
                564 / IN_WIDTH: ping_storage_data_780 <= (fillup_transition == 1'b1) ? i_input_data[564 % IN_WIDTH] : ping_storage_data_780 ^ i_input_data[564 % IN_WIDTH];
                737 / IN_WIDTH: ping_storage_data_780 <= (fillup_transition == 1'b1) ? i_input_data[737 % IN_WIDTH] : ping_storage_data_780 ^ i_input_data[737 % IN_WIDTH];
                1113 / IN_WIDTH: ping_storage_data_780 <= (fillup_transition == 1'b1) ? i_input_data[1113 % IN_WIDTH] : ping_storage_data_780 ^ i_input_data[1113 % IN_WIDTH];
                default: ping_storage_data_780 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_780;
                endcase
            end else begin
                case (input_count)
                0 / IN_WIDTH: pong_storage_data_780 <= (fillup_transition == 1'b1) ? i_input_data[0 % IN_WIDTH] : pong_storage_data_780 ^ i_input_data[0 % IN_WIDTH];
                409 / IN_WIDTH: pong_storage_data_780 <= (fillup_transition == 1'b1) ? i_input_data[409 % IN_WIDTH] : pong_storage_data_780 ^ i_input_data[409 % IN_WIDTH];
                564 / IN_WIDTH: pong_storage_data_780 <= (fillup_transition == 1'b1) ? i_input_data[564 % IN_WIDTH] : pong_storage_data_780 ^ i_input_data[564 % IN_WIDTH];
                737 / IN_WIDTH: pong_storage_data_780 <= (fillup_transition == 1'b1) ? i_input_data[737 % IN_WIDTH] : pong_storage_data_780 ^ i_input_data[737 % IN_WIDTH];
                1113 / IN_WIDTH: pong_storage_data_780 <= (fillup_transition == 1'b1) ? i_input_data[1113 % IN_WIDTH] : pong_storage_data_780 ^ i_input_data[1113 % IN_WIDTH];
                default: pong_storage_data_780 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_780;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_780 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_780;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_780 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_780;
            end
        end
    end
end

logic ping_storage_data_781;
logic pong_storage_data_781;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_781 <= 1'b0;
        pong_storage_data_781 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                1 / IN_WIDTH: ping_storage_data_781 <= (fillup_transition == 1'b1) ? i_input_data[1 % IN_WIDTH] : ping_storage_data_781 ^ i_input_data[1 % IN_WIDTH];
                410 / IN_WIDTH: ping_storage_data_781 <= (fillup_transition == 1'b1) ? i_input_data[410 % IN_WIDTH] : ping_storage_data_781 ^ i_input_data[410 % IN_WIDTH];
                565 / IN_WIDTH: ping_storage_data_781 <= (fillup_transition == 1'b1) ? i_input_data[565 % IN_WIDTH] : ping_storage_data_781 ^ i_input_data[565 % IN_WIDTH];
                738 / IN_WIDTH: ping_storage_data_781 <= (fillup_transition == 1'b1) ? i_input_data[738 % IN_WIDTH] : ping_storage_data_781 ^ i_input_data[738 % IN_WIDTH];
                1114 / IN_WIDTH: ping_storage_data_781 <= (fillup_transition == 1'b1) ? i_input_data[1114 % IN_WIDTH] : ping_storage_data_781 ^ i_input_data[1114 % IN_WIDTH];
                default: ping_storage_data_781 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_781;
                endcase
            end else begin
                case (input_count)
                1 / IN_WIDTH: pong_storage_data_781 <= (fillup_transition == 1'b1) ? i_input_data[1 % IN_WIDTH] : pong_storage_data_781 ^ i_input_data[1 % IN_WIDTH];
                410 / IN_WIDTH: pong_storage_data_781 <= (fillup_transition == 1'b1) ? i_input_data[410 % IN_WIDTH] : pong_storage_data_781 ^ i_input_data[410 % IN_WIDTH];
                565 / IN_WIDTH: pong_storage_data_781 <= (fillup_transition == 1'b1) ? i_input_data[565 % IN_WIDTH] : pong_storage_data_781 ^ i_input_data[565 % IN_WIDTH];
                738 / IN_WIDTH: pong_storage_data_781 <= (fillup_transition == 1'b1) ? i_input_data[738 % IN_WIDTH] : pong_storage_data_781 ^ i_input_data[738 % IN_WIDTH];
                1114 / IN_WIDTH: pong_storage_data_781 <= (fillup_transition == 1'b1) ? i_input_data[1114 % IN_WIDTH] : pong_storage_data_781 ^ i_input_data[1114 % IN_WIDTH];
                default: pong_storage_data_781 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_781;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_781 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_781;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_781 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_781;
            end
        end
    end
end

logic ping_storage_data_782;
logic pong_storage_data_782;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_782 <= 1'b0;
        pong_storage_data_782 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                2 / IN_WIDTH: ping_storage_data_782 <= (fillup_transition == 1'b1) ? i_input_data[2 % IN_WIDTH] : ping_storage_data_782 ^ i_input_data[2 % IN_WIDTH];
                411 / IN_WIDTH: ping_storage_data_782 <= (fillup_transition == 1'b1) ? i_input_data[411 % IN_WIDTH] : ping_storage_data_782 ^ i_input_data[411 % IN_WIDTH];
                566 / IN_WIDTH: ping_storage_data_782 <= (fillup_transition == 1'b1) ? i_input_data[566 % IN_WIDTH] : ping_storage_data_782 ^ i_input_data[566 % IN_WIDTH];
                739 / IN_WIDTH: ping_storage_data_782 <= (fillup_transition == 1'b1) ? i_input_data[739 % IN_WIDTH] : ping_storage_data_782 ^ i_input_data[739 % IN_WIDTH];
                1115 / IN_WIDTH: ping_storage_data_782 <= (fillup_transition == 1'b1) ? i_input_data[1115 % IN_WIDTH] : ping_storage_data_782 ^ i_input_data[1115 % IN_WIDTH];
                default: ping_storage_data_782 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_782;
                endcase
            end else begin
                case (input_count)
                2 / IN_WIDTH: pong_storage_data_782 <= (fillup_transition == 1'b1) ? i_input_data[2 % IN_WIDTH] : pong_storage_data_782 ^ i_input_data[2 % IN_WIDTH];
                411 / IN_WIDTH: pong_storage_data_782 <= (fillup_transition == 1'b1) ? i_input_data[411 % IN_WIDTH] : pong_storage_data_782 ^ i_input_data[411 % IN_WIDTH];
                566 / IN_WIDTH: pong_storage_data_782 <= (fillup_transition == 1'b1) ? i_input_data[566 % IN_WIDTH] : pong_storage_data_782 ^ i_input_data[566 % IN_WIDTH];
                739 / IN_WIDTH: pong_storage_data_782 <= (fillup_transition == 1'b1) ? i_input_data[739 % IN_WIDTH] : pong_storage_data_782 ^ i_input_data[739 % IN_WIDTH];
                1115 / IN_WIDTH: pong_storage_data_782 <= (fillup_transition == 1'b1) ? i_input_data[1115 % IN_WIDTH] : pong_storage_data_782 ^ i_input_data[1115 % IN_WIDTH];
                default: pong_storage_data_782 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_782;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_782 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_782;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_782 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_782;
            end
        end
    end
end

logic ping_storage_data_783;
logic pong_storage_data_783;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_783 <= 1'b0;
        pong_storage_data_783 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                3 / IN_WIDTH: ping_storage_data_783 <= (fillup_transition == 1'b1) ? i_input_data[3 % IN_WIDTH] : ping_storage_data_783 ^ i_input_data[3 % IN_WIDTH];
                412 / IN_WIDTH: ping_storage_data_783 <= (fillup_transition == 1'b1) ? i_input_data[412 % IN_WIDTH] : ping_storage_data_783 ^ i_input_data[412 % IN_WIDTH];
                567 / IN_WIDTH: ping_storage_data_783 <= (fillup_transition == 1'b1) ? i_input_data[567 % IN_WIDTH] : ping_storage_data_783 ^ i_input_data[567 % IN_WIDTH];
                740 / IN_WIDTH: ping_storage_data_783 <= (fillup_transition == 1'b1) ? i_input_data[740 % IN_WIDTH] : ping_storage_data_783 ^ i_input_data[740 % IN_WIDTH];
                1116 / IN_WIDTH: ping_storage_data_783 <= (fillup_transition == 1'b1) ? i_input_data[1116 % IN_WIDTH] : ping_storage_data_783 ^ i_input_data[1116 % IN_WIDTH];
                default: ping_storage_data_783 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_783;
                endcase
            end else begin
                case (input_count)
                3 / IN_WIDTH: pong_storage_data_783 <= (fillup_transition == 1'b1) ? i_input_data[3 % IN_WIDTH] : pong_storage_data_783 ^ i_input_data[3 % IN_WIDTH];
                412 / IN_WIDTH: pong_storage_data_783 <= (fillup_transition == 1'b1) ? i_input_data[412 % IN_WIDTH] : pong_storage_data_783 ^ i_input_data[412 % IN_WIDTH];
                567 / IN_WIDTH: pong_storage_data_783 <= (fillup_transition == 1'b1) ? i_input_data[567 % IN_WIDTH] : pong_storage_data_783 ^ i_input_data[567 % IN_WIDTH];
                740 / IN_WIDTH: pong_storage_data_783 <= (fillup_transition == 1'b1) ? i_input_data[740 % IN_WIDTH] : pong_storage_data_783 ^ i_input_data[740 % IN_WIDTH];
                1116 / IN_WIDTH: pong_storage_data_783 <= (fillup_transition == 1'b1) ? i_input_data[1116 % IN_WIDTH] : pong_storage_data_783 ^ i_input_data[1116 % IN_WIDTH];
                default: pong_storage_data_783 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_783;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_783 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_783;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_783 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_783;
            end
        end
    end
end

logic ping_storage_data_784;
logic pong_storage_data_784;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_784 <= 1'b0;
        pong_storage_data_784 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                4 / IN_WIDTH: ping_storage_data_784 <= (fillup_transition == 1'b1) ? i_input_data[4 % IN_WIDTH] : ping_storage_data_784 ^ i_input_data[4 % IN_WIDTH];
                413 / IN_WIDTH: ping_storage_data_784 <= (fillup_transition == 1'b1) ? i_input_data[413 % IN_WIDTH] : ping_storage_data_784 ^ i_input_data[413 % IN_WIDTH];
                568 / IN_WIDTH: ping_storage_data_784 <= (fillup_transition == 1'b1) ? i_input_data[568 % IN_WIDTH] : ping_storage_data_784 ^ i_input_data[568 % IN_WIDTH];
                741 / IN_WIDTH: ping_storage_data_784 <= (fillup_transition == 1'b1) ? i_input_data[741 % IN_WIDTH] : ping_storage_data_784 ^ i_input_data[741 % IN_WIDTH];
                1117 / IN_WIDTH: ping_storage_data_784 <= (fillup_transition == 1'b1) ? i_input_data[1117 % IN_WIDTH] : ping_storage_data_784 ^ i_input_data[1117 % IN_WIDTH];
                default: ping_storage_data_784 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_784;
                endcase
            end else begin
                case (input_count)
                4 / IN_WIDTH: pong_storage_data_784 <= (fillup_transition == 1'b1) ? i_input_data[4 % IN_WIDTH] : pong_storage_data_784 ^ i_input_data[4 % IN_WIDTH];
                413 / IN_WIDTH: pong_storage_data_784 <= (fillup_transition == 1'b1) ? i_input_data[413 % IN_WIDTH] : pong_storage_data_784 ^ i_input_data[413 % IN_WIDTH];
                568 / IN_WIDTH: pong_storage_data_784 <= (fillup_transition == 1'b1) ? i_input_data[568 % IN_WIDTH] : pong_storage_data_784 ^ i_input_data[568 % IN_WIDTH];
                741 / IN_WIDTH: pong_storage_data_784 <= (fillup_transition == 1'b1) ? i_input_data[741 % IN_WIDTH] : pong_storage_data_784 ^ i_input_data[741 % IN_WIDTH];
                1117 / IN_WIDTH: pong_storage_data_784 <= (fillup_transition == 1'b1) ? i_input_data[1117 % IN_WIDTH] : pong_storage_data_784 ^ i_input_data[1117 % IN_WIDTH];
                default: pong_storage_data_784 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_784;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_784 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_784;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_784 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_784;
            end
        end
    end
end

logic ping_storage_data_785;
logic pong_storage_data_785;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_785 <= 1'b0;
        pong_storage_data_785 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                5 / IN_WIDTH: ping_storage_data_785 <= (fillup_transition == 1'b1) ? i_input_data[5 % IN_WIDTH] : ping_storage_data_785 ^ i_input_data[5 % IN_WIDTH];
                414 / IN_WIDTH: ping_storage_data_785 <= (fillup_transition == 1'b1) ? i_input_data[414 % IN_WIDTH] : ping_storage_data_785 ^ i_input_data[414 % IN_WIDTH];
                569 / IN_WIDTH: ping_storage_data_785 <= (fillup_transition == 1'b1) ? i_input_data[569 % IN_WIDTH] : ping_storage_data_785 ^ i_input_data[569 % IN_WIDTH];
                742 / IN_WIDTH: ping_storage_data_785 <= (fillup_transition == 1'b1) ? i_input_data[742 % IN_WIDTH] : ping_storage_data_785 ^ i_input_data[742 % IN_WIDTH];
                1118 / IN_WIDTH: ping_storage_data_785 <= (fillup_transition == 1'b1) ? i_input_data[1118 % IN_WIDTH] : ping_storage_data_785 ^ i_input_data[1118 % IN_WIDTH];
                default: ping_storage_data_785 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_785;
                endcase
            end else begin
                case (input_count)
                5 / IN_WIDTH: pong_storage_data_785 <= (fillup_transition == 1'b1) ? i_input_data[5 % IN_WIDTH] : pong_storage_data_785 ^ i_input_data[5 % IN_WIDTH];
                414 / IN_WIDTH: pong_storage_data_785 <= (fillup_transition == 1'b1) ? i_input_data[414 % IN_WIDTH] : pong_storage_data_785 ^ i_input_data[414 % IN_WIDTH];
                569 / IN_WIDTH: pong_storage_data_785 <= (fillup_transition == 1'b1) ? i_input_data[569 % IN_WIDTH] : pong_storage_data_785 ^ i_input_data[569 % IN_WIDTH];
                742 / IN_WIDTH: pong_storage_data_785 <= (fillup_transition == 1'b1) ? i_input_data[742 % IN_WIDTH] : pong_storage_data_785 ^ i_input_data[742 % IN_WIDTH];
                1118 / IN_WIDTH: pong_storage_data_785 <= (fillup_transition == 1'b1) ? i_input_data[1118 % IN_WIDTH] : pong_storage_data_785 ^ i_input_data[1118 % IN_WIDTH];
                default: pong_storage_data_785 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_785;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_785 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_785;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_785 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_785;
            end
        end
    end
end

logic ping_storage_data_786;
logic pong_storage_data_786;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_786 <= 1'b0;
        pong_storage_data_786 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                6 / IN_WIDTH: ping_storage_data_786 <= (fillup_transition == 1'b1) ? i_input_data[6 % IN_WIDTH] : ping_storage_data_786 ^ i_input_data[6 % IN_WIDTH];
                415 / IN_WIDTH: ping_storage_data_786 <= (fillup_transition == 1'b1) ? i_input_data[415 % IN_WIDTH] : ping_storage_data_786 ^ i_input_data[415 % IN_WIDTH];
                570 / IN_WIDTH: ping_storage_data_786 <= (fillup_transition == 1'b1) ? i_input_data[570 % IN_WIDTH] : ping_storage_data_786 ^ i_input_data[570 % IN_WIDTH];
                743 / IN_WIDTH: ping_storage_data_786 <= (fillup_transition == 1'b1) ? i_input_data[743 % IN_WIDTH] : ping_storage_data_786 ^ i_input_data[743 % IN_WIDTH];
                1119 / IN_WIDTH: ping_storage_data_786 <= (fillup_transition == 1'b1) ? i_input_data[1119 % IN_WIDTH] : ping_storage_data_786 ^ i_input_data[1119 % IN_WIDTH];
                default: ping_storage_data_786 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_786;
                endcase
            end else begin
                case (input_count)
                6 / IN_WIDTH: pong_storage_data_786 <= (fillup_transition == 1'b1) ? i_input_data[6 % IN_WIDTH] : pong_storage_data_786 ^ i_input_data[6 % IN_WIDTH];
                415 / IN_WIDTH: pong_storage_data_786 <= (fillup_transition == 1'b1) ? i_input_data[415 % IN_WIDTH] : pong_storage_data_786 ^ i_input_data[415 % IN_WIDTH];
                570 / IN_WIDTH: pong_storage_data_786 <= (fillup_transition == 1'b1) ? i_input_data[570 % IN_WIDTH] : pong_storage_data_786 ^ i_input_data[570 % IN_WIDTH];
                743 / IN_WIDTH: pong_storage_data_786 <= (fillup_transition == 1'b1) ? i_input_data[743 % IN_WIDTH] : pong_storage_data_786 ^ i_input_data[743 % IN_WIDTH];
                1119 / IN_WIDTH: pong_storage_data_786 <= (fillup_transition == 1'b1) ? i_input_data[1119 % IN_WIDTH] : pong_storage_data_786 ^ i_input_data[1119 % IN_WIDTH];
                default: pong_storage_data_786 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_786;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_786 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_786;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_786 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_786;
            end
        end
    end
end

logic ping_storage_data_787;
logic pong_storage_data_787;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_787 <= 1'b0;
        pong_storage_data_787 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                7 / IN_WIDTH: ping_storage_data_787 <= (fillup_transition == 1'b1) ? i_input_data[7 % IN_WIDTH] : ping_storage_data_787 ^ i_input_data[7 % IN_WIDTH];
                416 / IN_WIDTH: ping_storage_data_787 <= (fillup_transition == 1'b1) ? i_input_data[416 % IN_WIDTH] : ping_storage_data_787 ^ i_input_data[416 % IN_WIDTH];
                571 / IN_WIDTH: ping_storage_data_787 <= (fillup_transition == 1'b1) ? i_input_data[571 % IN_WIDTH] : ping_storage_data_787 ^ i_input_data[571 % IN_WIDTH];
                744 / IN_WIDTH: ping_storage_data_787 <= (fillup_transition == 1'b1) ? i_input_data[744 % IN_WIDTH] : ping_storage_data_787 ^ i_input_data[744 % IN_WIDTH];
                1120 / IN_WIDTH: ping_storage_data_787 <= (fillup_transition == 1'b1) ? i_input_data[1120 % IN_WIDTH] : ping_storage_data_787 ^ i_input_data[1120 % IN_WIDTH];
                default: ping_storage_data_787 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_787;
                endcase
            end else begin
                case (input_count)
                7 / IN_WIDTH: pong_storage_data_787 <= (fillup_transition == 1'b1) ? i_input_data[7 % IN_WIDTH] : pong_storage_data_787 ^ i_input_data[7 % IN_WIDTH];
                416 / IN_WIDTH: pong_storage_data_787 <= (fillup_transition == 1'b1) ? i_input_data[416 % IN_WIDTH] : pong_storage_data_787 ^ i_input_data[416 % IN_WIDTH];
                571 / IN_WIDTH: pong_storage_data_787 <= (fillup_transition == 1'b1) ? i_input_data[571 % IN_WIDTH] : pong_storage_data_787 ^ i_input_data[571 % IN_WIDTH];
                744 / IN_WIDTH: pong_storage_data_787 <= (fillup_transition == 1'b1) ? i_input_data[744 % IN_WIDTH] : pong_storage_data_787 ^ i_input_data[744 % IN_WIDTH];
                1120 / IN_WIDTH: pong_storage_data_787 <= (fillup_transition == 1'b1) ? i_input_data[1120 % IN_WIDTH] : pong_storage_data_787 ^ i_input_data[1120 % IN_WIDTH];
                default: pong_storage_data_787 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_787;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_787 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_787;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_787 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_787;
            end
        end
    end
end

logic ping_storage_data_788;
logic pong_storage_data_788;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_788 <= 1'b0;
        pong_storage_data_788 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                8 / IN_WIDTH: ping_storage_data_788 <= (fillup_transition == 1'b1) ? i_input_data[8 % IN_WIDTH] : ping_storage_data_788 ^ i_input_data[8 % IN_WIDTH];
                417 / IN_WIDTH: ping_storage_data_788 <= (fillup_transition == 1'b1) ? i_input_data[417 % IN_WIDTH] : ping_storage_data_788 ^ i_input_data[417 % IN_WIDTH];
                572 / IN_WIDTH: ping_storage_data_788 <= (fillup_transition == 1'b1) ? i_input_data[572 % IN_WIDTH] : ping_storage_data_788 ^ i_input_data[572 % IN_WIDTH];
                745 / IN_WIDTH: ping_storage_data_788 <= (fillup_transition == 1'b1) ? i_input_data[745 % IN_WIDTH] : ping_storage_data_788 ^ i_input_data[745 % IN_WIDTH];
                1121 / IN_WIDTH: ping_storage_data_788 <= (fillup_transition == 1'b1) ? i_input_data[1121 % IN_WIDTH] : ping_storage_data_788 ^ i_input_data[1121 % IN_WIDTH];
                default: ping_storage_data_788 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_788;
                endcase
            end else begin
                case (input_count)
                8 / IN_WIDTH: pong_storage_data_788 <= (fillup_transition == 1'b1) ? i_input_data[8 % IN_WIDTH] : pong_storage_data_788 ^ i_input_data[8 % IN_WIDTH];
                417 / IN_WIDTH: pong_storage_data_788 <= (fillup_transition == 1'b1) ? i_input_data[417 % IN_WIDTH] : pong_storage_data_788 ^ i_input_data[417 % IN_WIDTH];
                572 / IN_WIDTH: pong_storage_data_788 <= (fillup_transition == 1'b1) ? i_input_data[572 % IN_WIDTH] : pong_storage_data_788 ^ i_input_data[572 % IN_WIDTH];
                745 / IN_WIDTH: pong_storage_data_788 <= (fillup_transition == 1'b1) ? i_input_data[745 % IN_WIDTH] : pong_storage_data_788 ^ i_input_data[745 % IN_WIDTH];
                1121 / IN_WIDTH: pong_storage_data_788 <= (fillup_transition == 1'b1) ? i_input_data[1121 % IN_WIDTH] : pong_storage_data_788 ^ i_input_data[1121 % IN_WIDTH];
                default: pong_storage_data_788 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_788;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_788 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_788;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_788 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_788;
            end
        end
    end
end

logic ping_storage_data_789;
logic pong_storage_data_789;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_789 <= 1'b0;
        pong_storage_data_789 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                9 / IN_WIDTH: ping_storage_data_789 <= (fillup_transition == 1'b1) ? i_input_data[9 % IN_WIDTH] : ping_storage_data_789 ^ i_input_data[9 % IN_WIDTH];
                418 / IN_WIDTH: ping_storage_data_789 <= (fillup_transition == 1'b1) ? i_input_data[418 % IN_WIDTH] : ping_storage_data_789 ^ i_input_data[418 % IN_WIDTH];
                573 / IN_WIDTH: ping_storage_data_789 <= (fillup_transition == 1'b1) ? i_input_data[573 % IN_WIDTH] : ping_storage_data_789 ^ i_input_data[573 % IN_WIDTH];
                746 / IN_WIDTH: ping_storage_data_789 <= (fillup_transition == 1'b1) ? i_input_data[746 % IN_WIDTH] : ping_storage_data_789 ^ i_input_data[746 % IN_WIDTH];
                1122 / IN_WIDTH: ping_storage_data_789 <= (fillup_transition == 1'b1) ? i_input_data[1122 % IN_WIDTH] : ping_storage_data_789 ^ i_input_data[1122 % IN_WIDTH];
                default: ping_storage_data_789 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_789;
                endcase
            end else begin
                case (input_count)
                9 / IN_WIDTH: pong_storage_data_789 <= (fillup_transition == 1'b1) ? i_input_data[9 % IN_WIDTH] : pong_storage_data_789 ^ i_input_data[9 % IN_WIDTH];
                418 / IN_WIDTH: pong_storage_data_789 <= (fillup_transition == 1'b1) ? i_input_data[418 % IN_WIDTH] : pong_storage_data_789 ^ i_input_data[418 % IN_WIDTH];
                573 / IN_WIDTH: pong_storage_data_789 <= (fillup_transition == 1'b1) ? i_input_data[573 % IN_WIDTH] : pong_storage_data_789 ^ i_input_data[573 % IN_WIDTH];
                746 / IN_WIDTH: pong_storage_data_789 <= (fillup_transition == 1'b1) ? i_input_data[746 % IN_WIDTH] : pong_storage_data_789 ^ i_input_data[746 % IN_WIDTH];
                1122 / IN_WIDTH: pong_storage_data_789 <= (fillup_transition == 1'b1) ? i_input_data[1122 % IN_WIDTH] : pong_storage_data_789 ^ i_input_data[1122 % IN_WIDTH];
                default: pong_storage_data_789 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_789;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_789 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_789;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_789 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_789;
            end
        end
    end
end

logic ping_storage_data_790;
logic pong_storage_data_790;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_790 <= 1'b0;
        pong_storage_data_790 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                10 / IN_WIDTH: ping_storage_data_790 <= (fillup_transition == 1'b1) ? i_input_data[10 % IN_WIDTH] : ping_storage_data_790 ^ i_input_data[10 % IN_WIDTH];
                419 / IN_WIDTH: ping_storage_data_790 <= (fillup_transition == 1'b1) ? i_input_data[419 % IN_WIDTH] : ping_storage_data_790 ^ i_input_data[419 % IN_WIDTH];
                574 / IN_WIDTH: ping_storage_data_790 <= (fillup_transition == 1'b1) ? i_input_data[574 % IN_WIDTH] : ping_storage_data_790 ^ i_input_data[574 % IN_WIDTH];
                747 / IN_WIDTH: ping_storage_data_790 <= (fillup_transition == 1'b1) ? i_input_data[747 % IN_WIDTH] : ping_storage_data_790 ^ i_input_data[747 % IN_WIDTH];
                1123 / IN_WIDTH: ping_storage_data_790 <= (fillup_transition == 1'b1) ? i_input_data[1123 % IN_WIDTH] : ping_storage_data_790 ^ i_input_data[1123 % IN_WIDTH];
                default: ping_storage_data_790 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_790;
                endcase
            end else begin
                case (input_count)
                10 / IN_WIDTH: pong_storage_data_790 <= (fillup_transition == 1'b1) ? i_input_data[10 % IN_WIDTH] : pong_storage_data_790 ^ i_input_data[10 % IN_WIDTH];
                419 / IN_WIDTH: pong_storage_data_790 <= (fillup_transition == 1'b1) ? i_input_data[419 % IN_WIDTH] : pong_storage_data_790 ^ i_input_data[419 % IN_WIDTH];
                574 / IN_WIDTH: pong_storage_data_790 <= (fillup_transition == 1'b1) ? i_input_data[574 % IN_WIDTH] : pong_storage_data_790 ^ i_input_data[574 % IN_WIDTH];
                747 / IN_WIDTH: pong_storage_data_790 <= (fillup_transition == 1'b1) ? i_input_data[747 % IN_WIDTH] : pong_storage_data_790 ^ i_input_data[747 % IN_WIDTH];
                1123 / IN_WIDTH: pong_storage_data_790 <= (fillup_transition == 1'b1) ? i_input_data[1123 % IN_WIDTH] : pong_storage_data_790 ^ i_input_data[1123 % IN_WIDTH];
                default: pong_storage_data_790 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_790;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_790 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_790;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_790 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_790;
            end
        end
    end
end

logic ping_storage_data_791;
logic pong_storage_data_791;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_791 <= 1'b0;
        pong_storage_data_791 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                11 / IN_WIDTH: ping_storage_data_791 <= (fillup_transition == 1'b1) ? i_input_data[11 % IN_WIDTH] : ping_storage_data_791 ^ i_input_data[11 % IN_WIDTH];
                420 / IN_WIDTH: ping_storage_data_791 <= (fillup_transition == 1'b1) ? i_input_data[420 % IN_WIDTH] : ping_storage_data_791 ^ i_input_data[420 % IN_WIDTH];
                575 / IN_WIDTH: ping_storage_data_791 <= (fillup_transition == 1'b1) ? i_input_data[575 % IN_WIDTH] : ping_storage_data_791 ^ i_input_data[575 % IN_WIDTH];
                748 / IN_WIDTH: ping_storage_data_791 <= (fillup_transition == 1'b1) ? i_input_data[748 % IN_WIDTH] : ping_storage_data_791 ^ i_input_data[748 % IN_WIDTH];
                1124 / IN_WIDTH: ping_storage_data_791 <= (fillup_transition == 1'b1) ? i_input_data[1124 % IN_WIDTH] : ping_storage_data_791 ^ i_input_data[1124 % IN_WIDTH];
                default: ping_storage_data_791 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_791;
                endcase
            end else begin
                case (input_count)
                11 / IN_WIDTH: pong_storage_data_791 <= (fillup_transition == 1'b1) ? i_input_data[11 % IN_WIDTH] : pong_storage_data_791 ^ i_input_data[11 % IN_WIDTH];
                420 / IN_WIDTH: pong_storage_data_791 <= (fillup_transition == 1'b1) ? i_input_data[420 % IN_WIDTH] : pong_storage_data_791 ^ i_input_data[420 % IN_WIDTH];
                575 / IN_WIDTH: pong_storage_data_791 <= (fillup_transition == 1'b1) ? i_input_data[575 % IN_WIDTH] : pong_storage_data_791 ^ i_input_data[575 % IN_WIDTH];
                748 / IN_WIDTH: pong_storage_data_791 <= (fillup_transition == 1'b1) ? i_input_data[748 % IN_WIDTH] : pong_storage_data_791 ^ i_input_data[748 % IN_WIDTH];
                1124 / IN_WIDTH: pong_storage_data_791 <= (fillup_transition == 1'b1) ? i_input_data[1124 % IN_WIDTH] : pong_storage_data_791 ^ i_input_data[1124 % IN_WIDTH];
                default: pong_storage_data_791 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_791;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_791 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_791;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_791 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_791;
            end
        end
    end
end

logic ping_storage_data_792;
logic pong_storage_data_792;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_792 <= 1'b0;
        pong_storage_data_792 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                12 / IN_WIDTH: ping_storage_data_792 <= (fillup_transition == 1'b1) ? i_input_data[12 % IN_WIDTH] : ping_storage_data_792 ^ i_input_data[12 % IN_WIDTH];
                421 / IN_WIDTH: ping_storage_data_792 <= (fillup_transition == 1'b1) ? i_input_data[421 % IN_WIDTH] : ping_storage_data_792 ^ i_input_data[421 % IN_WIDTH];
                480 / IN_WIDTH: ping_storage_data_792 <= (fillup_transition == 1'b1) ? i_input_data[480 % IN_WIDTH] : ping_storage_data_792 ^ i_input_data[480 % IN_WIDTH];
                749 / IN_WIDTH: ping_storage_data_792 <= (fillup_transition == 1'b1) ? i_input_data[749 % IN_WIDTH] : ping_storage_data_792 ^ i_input_data[749 % IN_WIDTH];
                1125 / IN_WIDTH: ping_storage_data_792 <= (fillup_transition == 1'b1) ? i_input_data[1125 % IN_WIDTH] : ping_storage_data_792 ^ i_input_data[1125 % IN_WIDTH];
                default: ping_storage_data_792 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_792;
                endcase
            end else begin
                case (input_count)
                12 / IN_WIDTH: pong_storage_data_792 <= (fillup_transition == 1'b1) ? i_input_data[12 % IN_WIDTH] : pong_storage_data_792 ^ i_input_data[12 % IN_WIDTH];
                421 / IN_WIDTH: pong_storage_data_792 <= (fillup_transition == 1'b1) ? i_input_data[421 % IN_WIDTH] : pong_storage_data_792 ^ i_input_data[421 % IN_WIDTH];
                480 / IN_WIDTH: pong_storage_data_792 <= (fillup_transition == 1'b1) ? i_input_data[480 % IN_WIDTH] : pong_storage_data_792 ^ i_input_data[480 % IN_WIDTH];
                749 / IN_WIDTH: pong_storage_data_792 <= (fillup_transition == 1'b1) ? i_input_data[749 % IN_WIDTH] : pong_storage_data_792 ^ i_input_data[749 % IN_WIDTH];
                1125 / IN_WIDTH: pong_storage_data_792 <= (fillup_transition == 1'b1) ? i_input_data[1125 % IN_WIDTH] : pong_storage_data_792 ^ i_input_data[1125 % IN_WIDTH];
                default: pong_storage_data_792 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_792;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_792 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_792;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_792 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_792;
            end
        end
    end
end

logic ping_storage_data_793;
logic pong_storage_data_793;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_793 <= 1'b0;
        pong_storage_data_793 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                13 / IN_WIDTH: ping_storage_data_793 <= (fillup_transition == 1'b1) ? i_input_data[13 % IN_WIDTH] : ping_storage_data_793 ^ i_input_data[13 % IN_WIDTH];
                422 / IN_WIDTH: ping_storage_data_793 <= (fillup_transition == 1'b1) ? i_input_data[422 % IN_WIDTH] : ping_storage_data_793 ^ i_input_data[422 % IN_WIDTH];
                481 / IN_WIDTH: ping_storage_data_793 <= (fillup_transition == 1'b1) ? i_input_data[481 % IN_WIDTH] : ping_storage_data_793 ^ i_input_data[481 % IN_WIDTH];
                750 / IN_WIDTH: ping_storage_data_793 <= (fillup_transition == 1'b1) ? i_input_data[750 % IN_WIDTH] : ping_storage_data_793 ^ i_input_data[750 % IN_WIDTH];
                1126 / IN_WIDTH: ping_storage_data_793 <= (fillup_transition == 1'b1) ? i_input_data[1126 % IN_WIDTH] : ping_storage_data_793 ^ i_input_data[1126 % IN_WIDTH];
                default: ping_storage_data_793 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_793;
                endcase
            end else begin
                case (input_count)
                13 / IN_WIDTH: pong_storage_data_793 <= (fillup_transition == 1'b1) ? i_input_data[13 % IN_WIDTH] : pong_storage_data_793 ^ i_input_data[13 % IN_WIDTH];
                422 / IN_WIDTH: pong_storage_data_793 <= (fillup_transition == 1'b1) ? i_input_data[422 % IN_WIDTH] : pong_storage_data_793 ^ i_input_data[422 % IN_WIDTH];
                481 / IN_WIDTH: pong_storage_data_793 <= (fillup_transition == 1'b1) ? i_input_data[481 % IN_WIDTH] : pong_storage_data_793 ^ i_input_data[481 % IN_WIDTH];
                750 / IN_WIDTH: pong_storage_data_793 <= (fillup_transition == 1'b1) ? i_input_data[750 % IN_WIDTH] : pong_storage_data_793 ^ i_input_data[750 % IN_WIDTH];
                1126 / IN_WIDTH: pong_storage_data_793 <= (fillup_transition == 1'b1) ? i_input_data[1126 % IN_WIDTH] : pong_storage_data_793 ^ i_input_data[1126 % IN_WIDTH];
                default: pong_storage_data_793 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_793;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_793 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_793;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_793 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_793;
            end
        end
    end
end

logic ping_storage_data_794;
logic pong_storage_data_794;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_794 <= 1'b0;
        pong_storage_data_794 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                14 / IN_WIDTH: ping_storage_data_794 <= (fillup_transition == 1'b1) ? i_input_data[14 % IN_WIDTH] : ping_storage_data_794 ^ i_input_data[14 % IN_WIDTH];
                423 / IN_WIDTH: ping_storage_data_794 <= (fillup_transition == 1'b1) ? i_input_data[423 % IN_WIDTH] : ping_storage_data_794 ^ i_input_data[423 % IN_WIDTH];
                482 / IN_WIDTH: ping_storage_data_794 <= (fillup_transition == 1'b1) ? i_input_data[482 % IN_WIDTH] : ping_storage_data_794 ^ i_input_data[482 % IN_WIDTH];
                751 / IN_WIDTH: ping_storage_data_794 <= (fillup_transition == 1'b1) ? i_input_data[751 % IN_WIDTH] : ping_storage_data_794 ^ i_input_data[751 % IN_WIDTH];
                1127 / IN_WIDTH: ping_storage_data_794 <= (fillup_transition == 1'b1) ? i_input_data[1127 % IN_WIDTH] : ping_storage_data_794 ^ i_input_data[1127 % IN_WIDTH];
                default: ping_storage_data_794 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_794;
                endcase
            end else begin
                case (input_count)
                14 / IN_WIDTH: pong_storage_data_794 <= (fillup_transition == 1'b1) ? i_input_data[14 % IN_WIDTH] : pong_storage_data_794 ^ i_input_data[14 % IN_WIDTH];
                423 / IN_WIDTH: pong_storage_data_794 <= (fillup_transition == 1'b1) ? i_input_data[423 % IN_WIDTH] : pong_storage_data_794 ^ i_input_data[423 % IN_WIDTH];
                482 / IN_WIDTH: pong_storage_data_794 <= (fillup_transition == 1'b1) ? i_input_data[482 % IN_WIDTH] : pong_storage_data_794 ^ i_input_data[482 % IN_WIDTH];
                751 / IN_WIDTH: pong_storage_data_794 <= (fillup_transition == 1'b1) ? i_input_data[751 % IN_WIDTH] : pong_storage_data_794 ^ i_input_data[751 % IN_WIDTH];
                1127 / IN_WIDTH: pong_storage_data_794 <= (fillup_transition == 1'b1) ? i_input_data[1127 % IN_WIDTH] : pong_storage_data_794 ^ i_input_data[1127 % IN_WIDTH];
                default: pong_storage_data_794 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_794;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_794 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_794;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_794 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_794;
            end
        end
    end
end

logic ping_storage_data_795;
logic pong_storage_data_795;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_795 <= 1'b0;
        pong_storage_data_795 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                15 / IN_WIDTH: ping_storage_data_795 <= (fillup_transition == 1'b1) ? i_input_data[15 % IN_WIDTH] : ping_storage_data_795 ^ i_input_data[15 % IN_WIDTH];
                424 / IN_WIDTH: ping_storage_data_795 <= (fillup_transition == 1'b1) ? i_input_data[424 % IN_WIDTH] : ping_storage_data_795 ^ i_input_data[424 % IN_WIDTH];
                483 / IN_WIDTH: ping_storage_data_795 <= (fillup_transition == 1'b1) ? i_input_data[483 % IN_WIDTH] : ping_storage_data_795 ^ i_input_data[483 % IN_WIDTH];
                752 / IN_WIDTH: ping_storage_data_795 <= (fillup_transition == 1'b1) ? i_input_data[752 % IN_WIDTH] : ping_storage_data_795 ^ i_input_data[752 % IN_WIDTH];
                1128 / IN_WIDTH: ping_storage_data_795 <= (fillup_transition == 1'b1) ? i_input_data[1128 % IN_WIDTH] : ping_storage_data_795 ^ i_input_data[1128 % IN_WIDTH];
                default: ping_storage_data_795 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_795;
                endcase
            end else begin
                case (input_count)
                15 / IN_WIDTH: pong_storage_data_795 <= (fillup_transition == 1'b1) ? i_input_data[15 % IN_WIDTH] : pong_storage_data_795 ^ i_input_data[15 % IN_WIDTH];
                424 / IN_WIDTH: pong_storage_data_795 <= (fillup_transition == 1'b1) ? i_input_data[424 % IN_WIDTH] : pong_storage_data_795 ^ i_input_data[424 % IN_WIDTH];
                483 / IN_WIDTH: pong_storage_data_795 <= (fillup_transition == 1'b1) ? i_input_data[483 % IN_WIDTH] : pong_storage_data_795 ^ i_input_data[483 % IN_WIDTH];
                752 / IN_WIDTH: pong_storage_data_795 <= (fillup_transition == 1'b1) ? i_input_data[752 % IN_WIDTH] : pong_storage_data_795 ^ i_input_data[752 % IN_WIDTH];
                1128 / IN_WIDTH: pong_storage_data_795 <= (fillup_transition == 1'b1) ? i_input_data[1128 % IN_WIDTH] : pong_storage_data_795 ^ i_input_data[1128 % IN_WIDTH];
                default: pong_storage_data_795 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_795;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_795 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_795;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_795 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_795;
            end
        end
    end
end

logic ping_storage_data_796;
logic pong_storage_data_796;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_796 <= 1'b0;
        pong_storage_data_796 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                16 / IN_WIDTH: ping_storage_data_796 <= (fillup_transition == 1'b1) ? i_input_data[16 % IN_WIDTH] : ping_storage_data_796 ^ i_input_data[16 % IN_WIDTH];
                425 / IN_WIDTH: ping_storage_data_796 <= (fillup_transition == 1'b1) ? i_input_data[425 % IN_WIDTH] : ping_storage_data_796 ^ i_input_data[425 % IN_WIDTH];
                484 / IN_WIDTH: ping_storage_data_796 <= (fillup_transition == 1'b1) ? i_input_data[484 % IN_WIDTH] : ping_storage_data_796 ^ i_input_data[484 % IN_WIDTH];
                753 / IN_WIDTH: ping_storage_data_796 <= (fillup_transition == 1'b1) ? i_input_data[753 % IN_WIDTH] : ping_storage_data_796 ^ i_input_data[753 % IN_WIDTH];
                1129 / IN_WIDTH: ping_storage_data_796 <= (fillup_transition == 1'b1) ? i_input_data[1129 % IN_WIDTH] : ping_storage_data_796 ^ i_input_data[1129 % IN_WIDTH];
                default: ping_storage_data_796 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_796;
                endcase
            end else begin
                case (input_count)
                16 / IN_WIDTH: pong_storage_data_796 <= (fillup_transition == 1'b1) ? i_input_data[16 % IN_WIDTH] : pong_storage_data_796 ^ i_input_data[16 % IN_WIDTH];
                425 / IN_WIDTH: pong_storage_data_796 <= (fillup_transition == 1'b1) ? i_input_data[425 % IN_WIDTH] : pong_storage_data_796 ^ i_input_data[425 % IN_WIDTH];
                484 / IN_WIDTH: pong_storage_data_796 <= (fillup_transition == 1'b1) ? i_input_data[484 % IN_WIDTH] : pong_storage_data_796 ^ i_input_data[484 % IN_WIDTH];
                753 / IN_WIDTH: pong_storage_data_796 <= (fillup_transition == 1'b1) ? i_input_data[753 % IN_WIDTH] : pong_storage_data_796 ^ i_input_data[753 % IN_WIDTH];
                1129 / IN_WIDTH: pong_storage_data_796 <= (fillup_transition == 1'b1) ? i_input_data[1129 % IN_WIDTH] : pong_storage_data_796 ^ i_input_data[1129 % IN_WIDTH];
                default: pong_storage_data_796 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_796;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_796 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_796;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_796 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_796;
            end
        end
    end
end

logic ping_storage_data_797;
logic pong_storage_data_797;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_797 <= 1'b0;
        pong_storage_data_797 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                17 / IN_WIDTH: ping_storage_data_797 <= (fillup_transition == 1'b1) ? i_input_data[17 % IN_WIDTH] : ping_storage_data_797 ^ i_input_data[17 % IN_WIDTH];
                426 / IN_WIDTH: ping_storage_data_797 <= (fillup_transition == 1'b1) ? i_input_data[426 % IN_WIDTH] : ping_storage_data_797 ^ i_input_data[426 % IN_WIDTH];
                485 / IN_WIDTH: ping_storage_data_797 <= (fillup_transition == 1'b1) ? i_input_data[485 % IN_WIDTH] : ping_storage_data_797 ^ i_input_data[485 % IN_WIDTH];
                754 / IN_WIDTH: ping_storage_data_797 <= (fillup_transition == 1'b1) ? i_input_data[754 % IN_WIDTH] : ping_storage_data_797 ^ i_input_data[754 % IN_WIDTH];
                1130 / IN_WIDTH: ping_storage_data_797 <= (fillup_transition == 1'b1) ? i_input_data[1130 % IN_WIDTH] : ping_storage_data_797 ^ i_input_data[1130 % IN_WIDTH];
                default: ping_storage_data_797 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_797;
                endcase
            end else begin
                case (input_count)
                17 / IN_WIDTH: pong_storage_data_797 <= (fillup_transition == 1'b1) ? i_input_data[17 % IN_WIDTH] : pong_storage_data_797 ^ i_input_data[17 % IN_WIDTH];
                426 / IN_WIDTH: pong_storage_data_797 <= (fillup_transition == 1'b1) ? i_input_data[426 % IN_WIDTH] : pong_storage_data_797 ^ i_input_data[426 % IN_WIDTH];
                485 / IN_WIDTH: pong_storage_data_797 <= (fillup_transition == 1'b1) ? i_input_data[485 % IN_WIDTH] : pong_storage_data_797 ^ i_input_data[485 % IN_WIDTH];
                754 / IN_WIDTH: pong_storage_data_797 <= (fillup_transition == 1'b1) ? i_input_data[754 % IN_WIDTH] : pong_storage_data_797 ^ i_input_data[754 % IN_WIDTH];
                1130 / IN_WIDTH: pong_storage_data_797 <= (fillup_transition == 1'b1) ? i_input_data[1130 % IN_WIDTH] : pong_storage_data_797 ^ i_input_data[1130 % IN_WIDTH];
                default: pong_storage_data_797 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_797;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_797 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_797;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_797 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_797;
            end
        end
    end
end

logic ping_storage_data_798;
logic pong_storage_data_798;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_798 <= 1'b0;
        pong_storage_data_798 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                18 / IN_WIDTH: ping_storage_data_798 <= (fillup_transition == 1'b1) ? i_input_data[18 % IN_WIDTH] : ping_storage_data_798 ^ i_input_data[18 % IN_WIDTH];
                427 / IN_WIDTH: ping_storage_data_798 <= (fillup_transition == 1'b1) ? i_input_data[427 % IN_WIDTH] : ping_storage_data_798 ^ i_input_data[427 % IN_WIDTH];
                486 / IN_WIDTH: ping_storage_data_798 <= (fillup_transition == 1'b1) ? i_input_data[486 % IN_WIDTH] : ping_storage_data_798 ^ i_input_data[486 % IN_WIDTH];
                755 / IN_WIDTH: ping_storage_data_798 <= (fillup_transition == 1'b1) ? i_input_data[755 % IN_WIDTH] : ping_storage_data_798 ^ i_input_data[755 % IN_WIDTH];
                1131 / IN_WIDTH: ping_storage_data_798 <= (fillup_transition == 1'b1) ? i_input_data[1131 % IN_WIDTH] : ping_storage_data_798 ^ i_input_data[1131 % IN_WIDTH];
                default: ping_storage_data_798 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_798;
                endcase
            end else begin
                case (input_count)
                18 / IN_WIDTH: pong_storage_data_798 <= (fillup_transition == 1'b1) ? i_input_data[18 % IN_WIDTH] : pong_storage_data_798 ^ i_input_data[18 % IN_WIDTH];
                427 / IN_WIDTH: pong_storage_data_798 <= (fillup_transition == 1'b1) ? i_input_data[427 % IN_WIDTH] : pong_storage_data_798 ^ i_input_data[427 % IN_WIDTH];
                486 / IN_WIDTH: pong_storage_data_798 <= (fillup_transition == 1'b1) ? i_input_data[486 % IN_WIDTH] : pong_storage_data_798 ^ i_input_data[486 % IN_WIDTH];
                755 / IN_WIDTH: pong_storage_data_798 <= (fillup_transition == 1'b1) ? i_input_data[755 % IN_WIDTH] : pong_storage_data_798 ^ i_input_data[755 % IN_WIDTH];
                1131 / IN_WIDTH: pong_storage_data_798 <= (fillup_transition == 1'b1) ? i_input_data[1131 % IN_WIDTH] : pong_storage_data_798 ^ i_input_data[1131 % IN_WIDTH];
                default: pong_storage_data_798 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_798;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_798 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_798;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_798 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_798;
            end
        end
    end
end

logic ping_storage_data_799;
logic pong_storage_data_799;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_799 <= 1'b0;
        pong_storage_data_799 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                19 / IN_WIDTH: ping_storage_data_799 <= (fillup_transition == 1'b1) ? i_input_data[19 % IN_WIDTH] : ping_storage_data_799 ^ i_input_data[19 % IN_WIDTH];
                428 / IN_WIDTH: ping_storage_data_799 <= (fillup_transition == 1'b1) ? i_input_data[428 % IN_WIDTH] : ping_storage_data_799 ^ i_input_data[428 % IN_WIDTH];
                487 / IN_WIDTH: ping_storage_data_799 <= (fillup_transition == 1'b1) ? i_input_data[487 % IN_WIDTH] : ping_storage_data_799 ^ i_input_data[487 % IN_WIDTH];
                756 / IN_WIDTH: ping_storage_data_799 <= (fillup_transition == 1'b1) ? i_input_data[756 % IN_WIDTH] : ping_storage_data_799 ^ i_input_data[756 % IN_WIDTH];
                1132 / IN_WIDTH: ping_storage_data_799 <= (fillup_transition == 1'b1) ? i_input_data[1132 % IN_WIDTH] : ping_storage_data_799 ^ i_input_data[1132 % IN_WIDTH];
                default: ping_storage_data_799 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_799;
                endcase
            end else begin
                case (input_count)
                19 / IN_WIDTH: pong_storage_data_799 <= (fillup_transition == 1'b1) ? i_input_data[19 % IN_WIDTH] : pong_storage_data_799 ^ i_input_data[19 % IN_WIDTH];
                428 / IN_WIDTH: pong_storage_data_799 <= (fillup_transition == 1'b1) ? i_input_data[428 % IN_WIDTH] : pong_storage_data_799 ^ i_input_data[428 % IN_WIDTH];
                487 / IN_WIDTH: pong_storage_data_799 <= (fillup_transition == 1'b1) ? i_input_data[487 % IN_WIDTH] : pong_storage_data_799 ^ i_input_data[487 % IN_WIDTH];
                756 / IN_WIDTH: pong_storage_data_799 <= (fillup_transition == 1'b1) ? i_input_data[756 % IN_WIDTH] : pong_storage_data_799 ^ i_input_data[756 % IN_WIDTH];
                1132 / IN_WIDTH: pong_storage_data_799 <= (fillup_transition == 1'b1) ? i_input_data[1132 % IN_WIDTH] : pong_storage_data_799 ^ i_input_data[1132 % IN_WIDTH];
                default: pong_storage_data_799 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_799;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_799 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_799;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_799 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_799;
            end
        end
    end
end

logic ping_storage_data_800;
logic pong_storage_data_800;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_800 <= 1'b0;
        pong_storage_data_800 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                20 / IN_WIDTH: ping_storage_data_800 <= (fillup_transition == 1'b1) ? i_input_data[20 % IN_WIDTH] : ping_storage_data_800 ^ i_input_data[20 % IN_WIDTH];
                429 / IN_WIDTH: ping_storage_data_800 <= (fillup_transition == 1'b1) ? i_input_data[429 % IN_WIDTH] : ping_storage_data_800 ^ i_input_data[429 % IN_WIDTH];
                488 / IN_WIDTH: ping_storage_data_800 <= (fillup_transition == 1'b1) ? i_input_data[488 % IN_WIDTH] : ping_storage_data_800 ^ i_input_data[488 % IN_WIDTH];
                757 / IN_WIDTH: ping_storage_data_800 <= (fillup_transition == 1'b1) ? i_input_data[757 % IN_WIDTH] : ping_storage_data_800 ^ i_input_data[757 % IN_WIDTH];
                1133 / IN_WIDTH: ping_storage_data_800 <= (fillup_transition == 1'b1) ? i_input_data[1133 % IN_WIDTH] : ping_storage_data_800 ^ i_input_data[1133 % IN_WIDTH];
                default: ping_storage_data_800 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_800;
                endcase
            end else begin
                case (input_count)
                20 / IN_WIDTH: pong_storage_data_800 <= (fillup_transition == 1'b1) ? i_input_data[20 % IN_WIDTH] : pong_storage_data_800 ^ i_input_data[20 % IN_WIDTH];
                429 / IN_WIDTH: pong_storage_data_800 <= (fillup_transition == 1'b1) ? i_input_data[429 % IN_WIDTH] : pong_storage_data_800 ^ i_input_data[429 % IN_WIDTH];
                488 / IN_WIDTH: pong_storage_data_800 <= (fillup_transition == 1'b1) ? i_input_data[488 % IN_WIDTH] : pong_storage_data_800 ^ i_input_data[488 % IN_WIDTH];
                757 / IN_WIDTH: pong_storage_data_800 <= (fillup_transition == 1'b1) ? i_input_data[757 % IN_WIDTH] : pong_storage_data_800 ^ i_input_data[757 % IN_WIDTH];
                1133 / IN_WIDTH: pong_storage_data_800 <= (fillup_transition == 1'b1) ? i_input_data[1133 % IN_WIDTH] : pong_storage_data_800 ^ i_input_data[1133 % IN_WIDTH];
                default: pong_storage_data_800 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_800;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_800 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_800;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_800 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_800;
            end
        end
    end
end

logic ping_storage_data_801;
logic pong_storage_data_801;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_801 <= 1'b0;
        pong_storage_data_801 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                21 / IN_WIDTH: ping_storage_data_801 <= (fillup_transition == 1'b1) ? i_input_data[21 % IN_WIDTH] : ping_storage_data_801 ^ i_input_data[21 % IN_WIDTH];
                430 / IN_WIDTH: ping_storage_data_801 <= (fillup_transition == 1'b1) ? i_input_data[430 % IN_WIDTH] : ping_storage_data_801 ^ i_input_data[430 % IN_WIDTH];
                489 / IN_WIDTH: ping_storage_data_801 <= (fillup_transition == 1'b1) ? i_input_data[489 % IN_WIDTH] : ping_storage_data_801 ^ i_input_data[489 % IN_WIDTH];
                758 / IN_WIDTH: ping_storage_data_801 <= (fillup_transition == 1'b1) ? i_input_data[758 % IN_WIDTH] : ping_storage_data_801 ^ i_input_data[758 % IN_WIDTH];
                1134 / IN_WIDTH: ping_storage_data_801 <= (fillup_transition == 1'b1) ? i_input_data[1134 % IN_WIDTH] : ping_storage_data_801 ^ i_input_data[1134 % IN_WIDTH];
                default: ping_storage_data_801 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_801;
                endcase
            end else begin
                case (input_count)
                21 / IN_WIDTH: pong_storage_data_801 <= (fillup_transition == 1'b1) ? i_input_data[21 % IN_WIDTH] : pong_storage_data_801 ^ i_input_data[21 % IN_WIDTH];
                430 / IN_WIDTH: pong_storage_data_801 <= (fillup_transition == 1'b1) ? i_input_data[430 % IN_WIDTH] : pong_storage_data_801 ^ i_input_data[430 % IN_WIDTH];
                489 / IN_WIDTH: pong_storage_data_801 <= (fillup_transition == 1'b1) ? i_input_data[489 % IN_WIDTH] : pong_storage_data_801 ^ i_input_data[489 % IN_WIDTH];
                758 / IN_WIDTH: pong_storage_data_801 <= (fillup_transition == 1'b1) ? i_input_data[758 % IN_WIDTH] : pong_storage_data_801 ^ i_input_data[758 % IN_WIDTH];
                1134 / IN_WIDTH: pong_storage_data_801 <= (fillup_transition == 1'b1) ? i_input_data[1134 % IN_WIDTH] : pong_storage_data_801 ^ i_input_data[1134 % IN_WIDTH];
                default: pong_storage_data_801 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_801;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_801 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_801;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_801 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_801;
            end
        end
    end
end

logic ping_storage_data_802;
logic pong_storage_data_802;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_802 <= 1'b0;
        pong_storage_data_802 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                22 / IN_WIDTH: ping_storage_data_802 <= (fillup_transition == 1'b1) ? i_input_data[22 % IN_WIDTH] : ping_storage_data_802 ^ i_input_data[22 % IN_WIDTH];
                431 / IN_WIDTH: ping_storage_data_802 <= (fillup_transition == 1'b1) ? i_input_data[431 % IN_WIDTH] : ping_storage_data_802 ^ i_input_data[431 % IN_WIDTH];
                490 / IN_WIDTH: ping_storage_data_802 <= (fillup_transition == 1'b1) ? i_input_data[490 % IN_WIDTH] : ping_storage_data_802 ^ i_input_data[490 % IN_WIDTH];
                759 / IN_WIDTH: ping_storage_data_802 <= (fillup_transition == 1'b1) ? i_input_data[759 % IN_WIDTH] : ping_storage_data_802 ^ i_input_data[759 % IN_WIDTH];
                1135 / IN_WIDTH: ping_storage_data_802 <= (fillup_transition == 1'b1) ? i_input_data[1135 % IN_WIDTH] : ping_storage_data_802 ^ i_input_data[1135 % IN_WIDTH];
                default: ping_storage_data_802 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_802;
                endcase
            end else begin
                case (input_count)
                22 / IN_WIDTH: pong_storage_data_802 <= (fillup_transition == 1'b1) ? i_input_data[22 % IN_WIDTH] : pong_storage_data_802 ^ i_input_data[22 % IN_WIDTH];
                431 / IN_WIDTH: pong_storage_data_802 <= (fillup_transition == 1'b1) ? i_input_data[431 % IN_WIDTH] : pong_storage_data_802 ^ i_input_data[431 % IN_WIDTH];
                490 / IN_WIDTH: pong_storage_data_802 <= (fillup_transition == 1'b1) ? i_input_data[490 % IN_WIDTH] : pong_storage_data_802 ^ i_input_data[490 % IN_WIDTH];
                759 / IN_WIDTH: pong_storage_data_802 <= (fillup_transition == 1'b1) ? i_input_data[759 % IN_WIDTH] : pong_storage_data_802 ^ i_input_data[759 % IN_WIDTH];
                1135 / IN_WIDTH: pong_storage_data_802 <= (fillup_transition == 1'b1) ? i_input_data[1135 % IN_WIDTH] : pong_storage_data_802 ^ i_input_data[1135 % IN_WIDTH];
                default: pong_storage_data_802 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_802;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_802 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_802;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_802 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_802;
            end
        end
    end
end

logic ping_storage_data_803;
logic pong_storage_data_803;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_803 <= 1'b0;
        pong_storage_data_803 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                23 / IN_WIDTH: ping_storage_data_803 <= (fillup_transition == 1'b1) ? i_input_data[23 % IN_WIDTH] : ping_storage_data_803 ^ i_input_data[23 % IN_WIDTH];
                432 / IN_WIDTH: ping_storage_data_803 <= (fillup_transition == 1'b1) ? i_input_data[432 % IN_WIDTH] : ping_storage_data_803 ^ i_input_data[432 % IN_WIDTH];
                491 / IN_WIDTH: ping_storage_data_803 <= (fillup_transition == 1'b1) ? i_input_data[491 % IN_WIDTH] : ping_storage_data_803 ^ i_input_data[491 % IN_WIDTH];
                760 / IN_WIDTH: ping_storage_data_803 <= (fillup_transition == 1'b1) ? i_input_data[760 % IN_WIDTH] : ping_storage_data_803 ^ i_input_data[760 % IN_WIDTH];
                1136 / IN_WIDTH: ping_storage_data_803 <= (fillup_transition == 1'b1) ? i_input_data[1136 % IN_WIDTH] : ping_storage_data_803 ^ i_input_data[1136 % IN_WIDTH];
                default: ping_storage_data_803 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_803;
                endcase
            end else begin
                case (input_count)
                23 / IN_WIDTH: pong_storage_data_803 <= (fillup_transition == 1'b1) ? i_input_data[23 % IN_WIDTH] : pong_storage_data_803 ^ i_input_data[23 % IN_WIDTH];
                432 / IN_WIDTH: pong_storage_data_803 <= (fillup_transition == 1'b1) ? i_input_data[432 % IN_WIDTH] : pong_storage_data_803 ^ i_input_data[432 % IN_WIDTH];
                491 / IN_WIDTH: pong_storage_data_803 <= (fillup_transition == 1'b1) ? i_input_data[491 % IN_WIDTH] : pong_storage_data_803 ^ i_input_data[491 % IN_WIDTH];
                760 / IN_WIDTH: pong_storage_data_803 <= (fillup_transition == 1'b1) ? i_input_data[760 % IN_WIDTH] : pong_storage_data_803 ^ i_input_data[760 % IN_WIDTH];
                1136 / IN_WIDTH: pong_storage_data_803 <= (fillup_transition == 1'b1) ? i_input_data[1136 % IN_WIDTH] : pong_storage_data_803 ^ i_input_data[1136 % IN_WIDTH];
                default: pong_storage_data_803 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_803;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_803 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_803;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_803 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_803;
            end
        end
    end
end

logic ping_storage_data_804;
logic pong_storage_data_804;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_804 <= 1'b0;
        pong_storage_data_804 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                24 / IN_WIDTH: ping_storage_data_804 <= (fillup_transition == 1'b1) ? i_input_data[24 % IN_WIDTH] : ping_storage_data_804 ^ i_input_data[24 % IN_WIDTH];
                433 / IN_WIDTH: ping_storage_data_804 <= (fillup_transition == 1'b1) ? i_input_data[433 % IN_WIDTH] : ping_storage_data_804 ^ i_input_data[433 % IN_WIDTH];
                492 / IN_WIDTH: ping_storage_data_804 <= (fillup_transition == 1'b1) ? i_input_data[492 % IN_WIDTH] : ping_storage_data_804 ^ i_input_data[492 % IN_WIDTH];
                761 / IN_WIDTH: ping_storage_data_804 <= (fillup_transition == 1'b1) ? i_input_data[761 % IN_WIDTH] : ping_storage_data_804 ^ i_input_data[761 % IN_WIDTH];
                1137 / IN_WIDTH: ping_storage_data_804 <= (fillup_transition == 1'b1) ? i_input_data[1137 % IN_WIDTH] : ping_storage_data_804 ^ i_input_data[1137 % IN_WIDTH];
                default: ping_storage_data_804 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_804;
                endcase
            end else begin
                case (input_count)
                24 / IN_WIDTH: pong_storage_data_804 <= (fillup_transition == 1'b1) ? i_input_data[24 % IN_WIDTH] : pong_storage_data_804 ^ i_input_data[24 % IN_WIDTH];
                433 / IN_WIDTH: pong_storage_data_804 <= (fillup_transition == 1'b1) ? i_input_data[433 % IN_WIDTH] : pong_storage_data_804 ^ i_input_data[433 % IN_WIDTH];
                492 / IN_WIDTH: pong_storage_data_804 <= (fillup_transition == 1'b1) ? i_input_data[492 % IN_WIDTH] : pong_storage_data_804 ^ i_input_data[492 % IN_WIDTH];
                761 / IN_WIDTH: pong_storage_data_804 <= (fillup_transition == 1'b1) ? i_input_data[761 % IN_WIDTH] : pong_storage_data_804 ^ i_input_data[761 % IN_WIDTH];
                1137 / IN_WIDTH: pong_storage_data_804 <= (fillup_transition == 1'b1) ? i_input_data[1137 % IN_WIDTH] : pong_storage_data_804 ^ i_input_data[1137 % IN_WIDTH];
                default: pong_storage_data_804 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_804;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_804 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_804;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_804 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_804;
            end
        end
    end
end

logic ping_storage_data_805;
logic pong_storage_data_805;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_805 <= 1'b0;
        pong_storage_data_805 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                25 / IN_WIDTH: ping_storage_data_805 <= (fillup_transition == 1'b1) ? i_input_data[25 % IN_WIDTH] : ping_storage_data_805 ^ i_input_data[25 % IN_WIDTH];
                434 / IN_WIDTH: ping_storage_data_805 <= (fillup_transition == 1'b1) ? i_input_data[434 % IN_WIDTH] : ping_storage_data_805 ^ i_input_data[434 % IN_WIDTH];
                493 / IN_WIDTH: ping_storage_data_805 <= (fillup_transition == 1'b1) ? i_input_data[493 % IN_WIDTH] : ping_storage_data_805 ^ i_input_data[493 % IN_WIDTH];
                762 / IN_WIDTH: ping_storage_data_805 <= (fillup_transition == 1'b1) ? i_input_data[762 % IN_WIDTH] : ping_storage_data_805 ^ i_input_data[762 % IN_WIDTH];
                1138 / IN_WIDTH: ping_storage_data_805 <= (fillup_transition == 1'b1) ? i_input_data[1138 % IN_WIDTH] : ping_storage_data_805 ^ i_input_data[1138 % IN_WIDTH];
                default: ping_storage_data_805 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_805;
                endcase
            end else begin
                case (input_count)
                25 / IN_WIDTH: pong_storage_data_805 <= (fillup_transition == 1'b1) ? i_input_data[25 % IN_WIDTH] : pong_storage_data_805 ^ i_input_data[25 % IN_WIDTH];
                434 / IN_WIDTH: pong_storage_data_805 <= (fillup_transition == 1'b1) ? i_input_data[434 % IN_WIDTH] : pong_storage_data_805 ^ i_input_data[434 % IN_WIDTH];
                493 / IN_WIDTH: pong_storage_data_805 <= (fillup_transition == 1'b1) ? i_input_data[493 % IN_WIDTH] : pong_storage_data_805 ^ i_input_data[493 % IN_WIDTH];
                762 / IN_WIDTH: pong_storage_data_805 <= (fillup_transition == 1'b1) ? i_input_data[762 % IN_WIDTH] : pong_storage_data_805 ^ i_input_data[762 % IN_WIDTH];
                1138 / IN_WIDTH: pong_storage_data_805 <= (fillup_transition == 1'b1) ? i_input_data[1138 % IN_WIDTH] : pong_storage_data_805 ^ i_input_data[1138 % IN_WIDTH];
                default: pong_storage_data_805 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_805;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_805 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_805;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_805 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_805;
            end
        end
    end
end

logic ping_storage_data_806;
logic pong_storage_data_806;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_806 <= 1'b0;
        pong_storage_data_806 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                26 / IN_WIDTH: ping_storage_data_806 <= (fillup_transition == 1'b1) ? i_input_data[26 % IN_WIDTH] : ping_storage_data_806 ^ i_input_data[26 % IN_WIDTH];
                435 / IN_WIDTH: ping_storage_data_806 <= (fillup_transition == 1'b1) ? i_input_data[435 % IN_WIDTH] : ping_storage_data_806 ^ i_input_data[435 % IN_WIDTH];
                494 / IN_WIDTH: ping_storage_data_806 <= (fillup_transition == 1'b1) ? i_input_data[494 % IN_WIDTH] : ping_storage_data_806 ^ i_input_data[494 % IN_WIDTH];
                763 / IN_WIDTH: ping_storage_data_806 <= (fillup_transition == 1'b1) ? i_input_data[763 % IN_WIDTH] : ping_storage_data_806 ^ i_input_data[763 % IN_WIDTH];
                1139 / IN_WIDTH: ping_storage_data_806 <= (fillup_transition == 1'b1) ? i_input_data[1139 % IN_WIDTH] : ping_storage_data_806 ^ i_input_data[1139 % IN_WIDTH];
                default: ping_storage_data_806 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_806;
                endcase
            end else begin
                case (input_count)
                26 / IN_WIDTH: pong_storage_data_806 <= (fillup_transition == 1'b1) ? i_input_data[26 % IN_WIDTH] : pong_storage_data_806 ^ i_input_data[26 % IN_WIDTH];
                435 / IN_WIDTH: pong_storage_data_806 <= (fillup_transition == 1'b1) ? i_input_data[435 % IN_WIDTH] : pong_storage_data_806 ^ i_input_data[435 % IN_WIDTH];
                494 / IN_WIDTH: pong_storage_data_806 <= (fillup_transition == 1'b1) ? i_input_data[494 % IN_WIDTH] : pong_storage_data_806 ^ i_input_data[494 % IN_WIDTH];
                763 / IN_WIDTH: pong_storage_data_806 <= (fillup_transition == 1'b1) ? i_input_data[763 % IN_WIDTH] : pong_storage_data_806 ^ i_input_data[763 % IN_WIDTH];
                1139 / IN_WIDTH: pong_storage_data_806 <= (fillup_transition == 1'b1) ? i_input_data[1139 % IN_WIDTH] : pong_storage_data_806 ^ i_input_data[1139 % IN_WIDTH];
                default: pong_storage_data_806 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_806;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_806 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_806;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_806 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_806;
            end
        end
    end
end

logic ping_storage_data_807;
logic pong_storage_data_807;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_807 <= 1'b0;
        pong_storage_data_807 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                27 / IN_WIDTH: ping_storage_data_807 <= (fillup_transition == 1'b1) ? i_input_data[27 % IN_WIDTH] : ping_storage_data_807 ^ i_input_data[27 % IN_WIDTH];
                436 / IN_WIDTH: ping_storage_data_807 <= (fillup_transition == 1'b1) ? i_input_data[436 % IN_WIDTH] : ping_storage_data_807 ^ i_input_data[436 % IN_WIDTH];
                495 / IN_WIDTH: ping_storage_data_807 <= (fillup_transition == 1'b1) ? i_input_data[495 % IN_WIDTH] : ping_storage_data_807 ^ i_input_data[495 % IN_WIDTH];
                764 / IN_WIDTH: ping_storage_data_807 <= (fillup_transition == 1'b1) ? i_input_data[764 % IN_WIDTH] : ping_storage_data_807 ^ i_input_data[764 % IN_WIDTH];
                1140 / IN_WIDTH: ping_storage_data_807 <= (fillup_transition == 1'b1) ? i_input_data[1140 % IN_WIDTH] : ping_storage_data_807 ^ i_input_data[1140 % IN_WIDTH];
                default: ping_storage_data_807 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_807;
                endcase
            end else begin
                case (input_count)
                27 / IN_WIDTH: pong_storage_data_807 <= (fillup_transition == 1'b1) ? i_input_data[27 % IN_WIDTH] : pong_storage_data_807 ^ i_input_data[27 % IN_WIDTH];
                436 / IN_WIDTH: pong_storage_data_807 <= (fillup_transition == 1'b1) ? i_input_data[436 % IN_WIDTH] : pong_storage_data_807 ^ i_input_data[436 % IN_WIDTH];
                495 / IN_WIDTH: pong_storage_data_807 <= (fillup_transition == 1'b1) ? i_input_data[495 % IN_WIDTH] : pong_storage_data_807 ^ i_input_data[495 % IN_WIDTH];
                764 / IN_WIDTH: pong_storage_data_807 <= (fillup_transition == 1'b1) ? i_input_data[764 % IN_WIDTH] : pong_storage_data_807 ^ i_input_data[764 % IN_WIDTH];
                1140 / IN_WIDTH: pong_storage_data_807 <= (fillup_transition == 1'b1) ? i_input_data[1140 % IN_WIDTH] : pong_storage_data_807 ^ i_input_data[1140 % IN_WIDTH];
                default: pong_storage_data_807 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_807;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_807 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_807;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_807 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_807;
            end
        end
    end
end

logic ping_storage_data_808;
logic pong_storage_data_808;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_808 <= 1'b0;
        pong_storage_data_808 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                28 / IN_WIDTH: ping_storage_data_808 <= (fillup_transition == 1'b1) ? i_input_data[28 % IN_WIDTH] : ping_storage_data_808 ^ i_input_data[28 % IN_WIDTH];
                437 / IN_WIDTH: ping_storage_data_808 <= (fillup_transition == 1'b1) ? i_input_data[437 % IN_WIDTH] : ping_storage_data_808 ^ i_input_data[437 % IN_WIDTH];
                496 / IN_WIDTH: ping_storage_data_808 <= (fillup_transition == 1'b1) ? i_input_data[496 % IN_WIDTH] : ping_storage_data_808 ^ i_input_data[496 % IN_WIDTH];
                765 / IN_WIDTH: ping_storage_data_808 <= (fillup_transition == 1'b1) ? i_input_data[765 % IN_WIDTH] : ping_storage_data_808 ^ i_input_data[765 % IN_WIDTH];
                1141 / IN_WIDTH: ping_storage_data_808 <= (fillup_transition == 1'b1) ? i_input_data[1141 % IN_WIDTH] : ping_storage_data_808 ^ i_input_data[1141 % IN_WIDTH];
                default: ping_storage_data_808 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_808;
                endcase
            end else begin
                case (input_count)
                28 / IN_WIDTH: pong_storage_data_808 <= (fillup_transition == 1'b1) ? i_input_data[28 % IN_WIDTH] : pong_storage_data_808 ^ i_input_data[28 % IN_WIDTH];
                437 / IN_WIDTH: pong_storage_data_808 <= (fillup_transition == 1'b1) ? i_input_data[437 % IN_WIDTH] : pong_storage_data_808 ^ i_input_data[437 % IN_WIDTH];
                496 / IN_WIDTH: pong_storage_data_808 <= (fillup_transition == 1'b1) ? i_input_data[496 % IN_WIDTH] : pong_storage_data_808 ^ i_input_data[496 % IN_WIDTH];
                765 / IN_WIDTH: pong_storage_data_808 <= (fillup_transition == 1'b1) ? i_input_data[765 % IN_WIDTH] : pong_storage_data_808 ^ i_input_data[765 % IN_WIDTH];
                1141 / IN_WIDTH: pong_storage_data_808 <= (fillup_transition == 1'b1) ? i_input_data[1141 % IN_WIDTH] : pong_storage_data_808 ^ i_input_data[1141 % IN_WIDTH];
                default: pong_storage_data_808 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_808;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_808 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_808;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_808 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_808;
            end
        end
    end
end

logic ping_storage_data_809;
logic pong_storage_data_809;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_809 <= 1'b0;
        pong_storage_data_809 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                29 / IN_WIDTH: ping_storage_data_809 <= (fillup_transition == 1'b1) ? i_input_data[29 % IN_WIDTH] : ping_storage_data_809 ^ i_input_data[29 % IN_WIDTH];
                438 / IN_WIDTH: ping_storage_data_809 <= (fillup_transition == 1'b1) ? i_input_data[438 % IN_WIDTH] : ping_storage_data_809 ^ i_input_data[438 % IN_WIDTH];
                497 / IN_WIDTH: ping_storage_data_809 <= (fillup_transition == 1'b1) ? i_input_data[497 % IN_WIDTH] : ping_storage_data_809 ^ i_input_data[497 % IN_WIDTH];
                766 / IN_WIDTH: ping_storage_data_809 <= (fillup_transition == 1'b1) ? i_input_data[766 % IN_WIDTH] : ping_storage_data_809 ^ i_input_data[766 % IN_WIDTH];
                1142 / IN_WIDTH: ping_storage_data_809 <= (fillup_transition == 1'b1) ? i_input_data[1142 % IN_WIDTH] : ping_storage_data_809 ^ i_input_data[1142 % IN_WIDTH];
                default: ping_storage_data_809 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_809;
                endcase
            end else begin
                case (input_count)
                29 / IN_WIDTH: pong_storage_data_809 <= (fillup_transition == 1'b1) ? i_input_data[29 % IN_WIDTH] : pong_storage_data_809 ^ i_input_data[29 % IN_WIDTH];
                438 / IN_WIDTH: pong_storage_data_809 <= (fillup_transition == 1'b1) ? i_input_data[438 % IN_WIDTH] : pong_storage_data_809 ^ i_input_data[438 % IN_WIDTH];
                497 / IN_WIDTH: pong_storage_data_809 <= (fillup_transition == 1'b1) ? i_input_data[497 % IN_WIDTH] : pong_storage_data_809 ^ i_input_data[497 % IN_WIDTH];
                766 / IN_WIDTH: pong_storage_data_809 <= (fillup_transition == 1'b1) ? i_input_data[766 % IN_WIDTH] : pong_storage_data_809 ^ i_input_data[766 % IN_WIDTH];
                1142 / IN_WIDTH: pong_storage_data_809 <= (fillup_transition == 1'b1) ? i_input_data[1142 % IN_WIDTH] : pong_storage_data_809 ^ i_input_data[1142 % IN_WIDTH];
                default: pong_storage_data_809 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_809;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_809 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_809;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_809 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_809;
            end
        end
    end
end

logic ping_storage_data_810;
logic pong_storage_data_810;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_810 <= 1'b0;
        pong_storage_data_810 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                30 / IN_WIDTH: ping_storage_data_810 <= (fillup_transition == 1'b1) ? i_input_data[30 % IN_WIDTH] : ping_storage_data_810 ^ i_input_data[30 % IN_WIDTH];
                439 / IN_WIDTH: ping_storage_data_810 <= (fillup_transition == 1'b1) ? i_input_data[439 % IN_WIDTH] : ping_storage_data_810 ^ i_input_data[439 % IN_WIDTH];
                498 / IN_WIDTH: ping_storage_data_810 <= (fillup_transition == 1'b1) ? i_input_data[498 % IN_WIDTH] : ping_storage_data_810 ^ i_input_data[498 % IN_WIDTH];
                767 / IN_WIDTH: ping_storage_data_810 <= (fillup_transition == 1'b1) ? i_input_data[767 % IN_WIDTH] : ping_storage_data_810 ^ i_input_data[767 % IN_WIDTH];
                1143 / IN_WIDTH: ping_storage_data_810 <= (fillup_transition == 1'b1) ? i_input_data[1143 % IN_WIDTH] : ping_storage_data_810 ^ i_input_data[1143 % IN_WIDTH];
                default: ping_storage_data_810 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_810;
                endcase
            end else begin
                case (input_count)
                30 / IN_WIDTH: pong_storage_data_810 <= (fillup_transition == 1'b1) ? i_input_data[30 % IN_WIDTH] : pong_storage_data_810 ^ i_input_data[30 % IN_WIDTH];
                439 / IN_WIDTH: pong_storage_data_810 <= (fillup_transition == 1'b1) ? i_input_data[439 % IN_WIDTH] : pong_storage_data_810 ^ i_input_data[439 % IN_WIDTH];
                498 / IN_WIDTH: pong_storage_data_810 <= (fillup_transition == 1'b1) ? i_input_data[498 % IN_WIDTH] : pong_storage_data_810 ^ i_input_data[498 % IN_WIDTH];
                767 / IN_WIDTH: pong_storage_data_810 <= (fillup_transition == 1'b1) ? i_input_data[767 % IN_WIDTH] : pong_storage_data_810 ^ i_input_data[767 % IN_WIDTH];
                1143 / IN_WIDTH: pong_storage_data_810 <= (fillup_transition == 1'b1) ? i_input_data[1143 % IN_WIDTH] : pong_storage_data_810 ^ i_input_data[1143 % IN_WIDTH];
                default: pong_storage_data_810 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_810;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_810 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_810;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_810 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_810;
            end
        end
    end
end

logic ping_storage_data_811;
logic pong_storage_data_811;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_811 <= 1'b0;
        pong_storage_data_811 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                31 / IN_WIDTH: ping_storage_data_811 <= (fillup_transition == 1'b1) ? i_input_data[31 % IN_WIDTH] : ping_storage_data_811 ^ i_input_data[31 % IN_WIDTH];
                440 / IN_WIDTH: ping_storage_data_811 <= (fillup_transition == 1'b1) ? i_input_data[440 % IN_WIDTH] : ping_storage_data_811 ^ i_input_data[440 % IN_WIDTH];
                499 / IN_WIDTH: ping_storage_data_811 <= (fillup_transition == 1'b1) ? i_input_data[499 % IN_WIDTH] : ping_storage_data_811 ^ i_input_data[499 % IN_WIDTH];
                672 / IN_WIDTH: ping_storage_data_811 <= (fillup_transition == 1'b1) ? i_input_data[672 % IN_WIDTH] : ping_storage_data_811 ^ i_input_data[672 % IN_WIDTH];
                1144 / IN_WIDTH: ping_storage_data_811 <= (fillup_transition == 1'b1) ? i_input_data[1144 % IN_WIDTH] : ping_storage_data_811 ^ i_input_data[1144 % IN_WIDTH];
                default: ping_storage_data_811 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_811;
                endcase
            end else begin
                case (input_count)
                31 / IN_WIDTH: pong_storage_data_811 <= (fillup_transition == 1'b1) ? i_input_data[31 % IN_WIDTH] : pong_storage_data_811 ^ i_input_data[31 % IN_WIDTH];
                440 / IN_WIDTH: pong_storage_data_811 <= (fillup_transition == 1'b1) ? i_input_data[440 % IN_WIDTH] : pong_storage_data_811 ^ i_input_data[440 % IN_WIDTH];
                499 / IN_WIDTH: pong_storage_data_811 <= (fillup_transition == 1'b1) ? i_input_data[499 % IN_WIDTH] : pong_storage_data_811 ^ i_input_data[499 % IN_WIDTH];
                672 / IN_WIDTH: pong_storage_data_811 <= (fillup_transition == 1'b1) ? i_input_data[672 % IN_WIDTH] : pong_storage_data_811 ^ i_input_data[672 % IN_WIDTH];
                1144 / IN_WIDTH: pong_storage_data_811 <= (fillup_transition == 1'b1) ? i_input_data[1144 % IN_WIDTH] : pong_storage_data_811 ^ i_input_data[1144 % IN_WIDTH];
                default: pong_storage_data_811 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_811;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_811 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_811;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_811 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_811;
            end
        end
    end
end

logic ping_storage_data_812;
logic pong_storage_data_812;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_812 <= 1'b0;
        pong_storage_data_812 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                32 / IN_WIDTH: ping_storage_data_812 <= (fillup_transition == 1'b1) ? i_input_data[32 % IN_WIDTH] : ping_storage_data_812 ^ i_input_data[32 % IN_WIDTH];
                441 / IN_WIDTH: ping_storage_data_812 <= (fillup_transition == 1'b1) ? i_input_data[441 % IN_WIDTH] : ping_storage_data_812 ^ i_input_data[441 % IN_WIDTH];
                500 / IN_WIDTH: ping_storage_data_812 <= (fillup_transition == 1'b1) ? i_input_data[500 % IN_WIDTH] : ping_storage_data_812 ^ i_input_data[500 % IN_WIDTH];
                673 / IN_WIDTH: ping_storage_data_812 <= (fillup_transition == 1'b1) ? i_input_data[673 % IN_WIDTH] : ping_storage_data_812 ^ i_input_data[673 % IN_WIDTH];
                1145 / IN_WIDTH: ping_storage_data_812 <= (fillup_transition == 1'b1) ? i_input_data[1145 % IN_WIDTH] : ping_storage_data_812 ^ i_input_data[1145 % IN_WIDTH];
                default: ping_storage_data_812 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_812;
                endcase
            end else begin
                case (input_count)
                32 / IN_WIDTH: pong_storage_data_812 <= (fillup_transition == 1'b1) ? i_input_data[32 % IN_WIDTH] : pong_storage_data_812 ^ i_input_data[32 % IN_WIDTH];
                441 / IN_WIDTH: pong_storage_data_812 <= (fillup_transition == 1'b1) ? i_input_data[441 % IN_WIDTH] : pong_storage_data_812 ^ i_input_data[441 % IN_WIDTH];
                500 / IN_WIDTH: pong_storage_data_812 <= (fillup_transition == 1'b1) ? i_input_data[500 % IN_WIDTH] : pong_storage_data_812 ^ i_input_data[500 % IN_WIDTH];
                673 / IN_WIDTH: pong_storage_data_812 <= (fillup_transition == 1'b1) ? i_input_data[673 % IN_WIDTH] : pong_storage_data_812 ^ i_input_data[673 % IN_WIDTH];
                1145 / IN_WIDTH: pong_storage_data_812 <= (fillup_transition == 1'b1) ? i_input_data[1145 % IN_WIDTH] : pong_storage_data_812 ^ i_input_data[1145 % IN_WIDTH];
                default: pong_storage_data_812 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_812;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_812 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_812;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_812 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_812;
            end
        end
    end
end

logic ping_storage_data_813;
logic pong_storage_data_813;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_813 <= 1'b0;
        pong_storage_data_813 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                33 / IN_WIDTH: ping_storage_data_813 <= (fillup_transition == 1'b1) ? i_input_data[33 % IN_WIDTH] : ping_storage_data_813 ^ i_input_data[33 % IN_WIDTH];
                442 / IN_WIDTH: ping_storage_data_813 <= (fillup_transition == 1'b1) ? i_input_data[442 % IN_WIDTH] : ping_storage_data_813 ^ i_input_data[442 % IN_WIDTH];
                501 / IN_WIDTH: ping_storage_data_813 <= (fillup_transition == 1'b1) ? i_input_data[501 % IN_WIDTH] : ping_storage_data_813 ^ i_input_data[501 % IN_WIDTH];
                674 / IN_WIDTH: ping_storage_data_813 <= (fillup_transition == 1'b1) ? i_input_data[674 % IN_WIDTH] : ping_storage_data_813 ^ i_input_data[674 % IN_WIDTH];
                1146 / IN_WIDTH: ping_storage_data_813 <= (fillup_transition == 1'b1) ? i_input_data[1146 % IN_WIDTH] : ping_storage_data_813 ^ i_input_data[1146 % IN_WIDTH];
                default: ping_storage_data_813 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_813;
                endcase
            end else begin
                case (input_count)
                33 / IN_WIDTH: pong_storage_data_813 <= (fillup_transition == 1'b1) ? i_input_data[33 % IN_WIDTH] : pong_storage_data_813 ^ i_input_data[33 % IN_WIDTH];
                442 / IN_WIDTH: pong_storage_data_813 <= (fillup_transition == 1'b1) ? i_input_data[442 % IN_WIDTH] : pong_storage_data_813 ^ i_input_data[442 % IN_WIDTH];
                501 / IN_WIDTH: pong_storage_data_813 <= (fillup_transition == 1'b1) ? i_input_data[501 % IN_WIDTH] : pong_storage_data_813 ^ i_input_data[501 % IN_WIDTH];
                674 / IN_WIDTH: pong_storage_data_813 <= (fillup_transition == 1'b1) ? i_input_data[674 % IN_WIDTH] : pong_storage_data_813 ^ i_input_data[674 % IN_WIDTH];
                1146 / IN_WIDTH: pong_storage_data_813 <= (fillup_transition == 1'b1) ? i_input_data[1146 % IN_WIDTH] : pong_storage_data_813 ^ i_input_data[1146 % IN_WIDTH];
                default: pong_storage_data_813 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_813;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_813 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_813;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_813 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_813;
            end
        end
    end
end

logic ping_storage_data_814;
logic pong_storage_data_814;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_814 <= 1'b0;
        pong_storage_data_814 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                34 / IN_WIDTH: ping_storage_data_814 <= (fillup_transition == 1'b1) ? i_input_data[34 % IN_WIDTH] : ping_storage_data_814 ^ i_input_data[34 % IN_WIDTH];
                443 / IN_WIDTH: ping_storage_data_814 <= (fillup_transition == 1'b1) ? i_input_data[443 % IN_WIDTH] : ping_storage_data_814 ^ i_input_data[443 % IN_WIDTH];
                502 / IN_WIDTH: ping_storage_data_814 <= (fillup_transition == 1'b1) ? i_input_data[502 % IN_WIDTH] : ping_storage_data_814 ^ i_input_data[502 % IN_WIDTH];
                675 / IN_WIDTH: ping_storage_data_814 <= (fillup_transition == 1'b1) ? i_input_data[675 % IN_WIDTH] : ping_storage_data_814 ^ i_input_data[675 % IN_WIDTH];
                1147 / IN_WIDTH: ping_storage_data_814 <= (fillup_transition == 1'b1) ? i_input_data[1147 % IN_WIDTH] : ping_storage_data_814 ^ i_input_data[1147 % IN_WIDTH];
                default: ping_storage_data_814 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_814;
                endcase
            end else begin
                case (input_count)
                34 / IN_WIDTH: pong_storage_data_814 <= (fillup_transition == 1'b1) ? i_input_data[34 % IN_WIDTH] : pong_storage_data_814 ^ i_input_data[34 % IN_WIDTH];
                443 / IN_WIDTH: pong_storage_data_814 <= (fillup_transition == 1'b1) ? i_input_data[443 % IN_WIDTH] : pong_storage_data_814 ^ i_input_data[443 % IN_WIDTH];
                502 / IN_WIDTH: pong_storage_data_814 <= (fillup_transition == 1'b1) ? i_input_data[502 % IN_WIDTH] : pong_storage_data_814 ^ i_input_data[502 % IN_WIDTH];
                675 / IN_WIDTH: pong_storage_data_814 <= (fillup_transition == 1'b1) ? i_input_data[675 % IN_WIDTH] : pong_storage_data_814 ^ i_input_data[675 % IN_WIDTH];
                1147 / IN_WIDTH: pong_storage_data_814 <= (fillup_transition == 1'b1) ? i_input_data[1147 % IN_WIDTH] : pong_storage_data_814 ^ i_input_data[1147 % IN_WIDTH];
                default: pong_storage_data_814 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_814;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_814 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_814;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_814 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_814;
            end
        end
    end
end

logic ping_storage_data_815;
logic pong_storage_data_815;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_815 <= 1'b0;
        pong_storage_data_815 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                35 / IN_WIDTH: ping_storage_data_815 <= (fillup_transition == 1'b1) ? i_input_data[35 % IN_WIDTH] : ping_storage_data_815 ^ i_input_data[35 % IN_WIDTH];
                444 / IN_WIDTH: ping_storage_data_815 <= (fillup_transition == 1'b1) ? i_input_data[444 % IN_WIDTH] : ping_storage_data_815 ^ i_input_data[444 % IN_WIDTH];
                503 / IN_WIDTH: ping_storage_data_815 <= (fillup_transition == 1'b1) ? i_input_data[503 % IN_WIDTH] : ping_storage_data_815 ^ i_input_data[503 % IN_WIDTH];
                676 / IN_WIDTH: ping_storage_data_815 <= (fillup_transition == 1'b1) ? i_input_data[676 % IN_WIDTH] : ping_storage_data_815 ^ i_input_data[676 % IN_WIDTH];
                1148 / IN_WIDTH: ping_storage_data_815 <= (fillup_transition == 1'b1) ? i_input_data[1148 % IN_WIDTH] : ping_storage_data_815 ^ i_input_data[1148 % IN_WIDTH];
                default: ping_storage_data_815 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_815;
                endcase
            end else begin
                case (input_count)
                35 / IN_WIDTH: pong_storage_data_815 <= (fillup_transition == 1'b1) ? i_input_data[35 % IN_WIDTH] : pong_storage_data_815 ^ i_input_data[35 % IN_WIDTH];
                444 / IN_WIDTH: pong_storage_data_815 <= (fillup_transition == 1'b1) ? i_input_data[444 % IN_WIDTH] : pong_storage_data_815 ^ i_input_data[444 % IN_WIDTH];
                503 / IN_WIDTH: pong_storage_data_815 <= (fillup_transition == 1'b1) ? i_input_data[503 % IN_WIDTH] : pong_storage_data_815 ^ i_input_data[503 % IN_WIDTH];
                676 / IN_WIDTH: pong_storage_data_815 <= (fillup_transition == 1'b1) ? i_input_data[676 % IN_WIDTH] : pong_storage_data_815 ^ i_input_data[676 % IN_WIDTH];
                1148 / IN_WIDTH: pong_storage_data_815 <= (fillup_transition == 1'b1) ? i_input_data[1148 % IN_WIDTH] : pong_storage_data_815 ^ i_input_data[1148 % IN_WIDTH];
                default: pong_storage_data_815 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_815;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_815 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_815;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_815 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_815;
            end
        end
    end
end

logic ping_storage_data_816;
logic pong_storage_data_816;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_816 <= 1'b0;
        pong_storage_data_816 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                36 / IN_WIDTH: ping_storage_data_816 <= (fillup_transition == 1'b1) ? i_input_data[36 % IN_WIDTH] : ping_storage_data_816 ^ i_input_data[36 % IN_WIDTH];
                445 / IN_WIDTH: ping_storage_data_816 <= (fillup_transition == 1'b1) ? i_input_data[445 % IN_WIDTH] : ping_storage_data_816 ^ i_input_data[445 % IN_WIDTH];
                504 / IN_WIDTH: ping_storage_data_816 <= (fillup_transition == 1'b1) ? i_input_data[504 % IN_WIDTH] : ping_storage_data_816 ^ i_input_data[504 % IN_WIDTH];
                677 / IN_WIDTH: ping_storage_data_816 <= (fillup_transition == 1'b1) ? i_input_data[677 % IN_WIDTH] : ping_storage_data_816 ^ i_input_data[677 % IN_WIDTH];
                1149 / IN_WIDTH: ping_storage_data_816 <= (fillup_transition == 1'b1) ? i_input_data[1149 % IN_WIDTH] : ping_storage_data_816 ^ i_input_data[1149 % IN_WIDTH];
                default: ping_storage_data_816 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_816;
                endcase
            end else begin
                case (input_count)
                36 / IN_WIDTH: pong_storage_data_816 <= (fillup_transition == 1'b1) ? i_input_data[36 % IN_WIDTH] : pong_storage_data_816 ^ i_input_data[36 % IN_WIDTH];
                445 / IN_WIDTH: pong_storage_data_816 <= (fillup_transition == 1'b1) ? i_input_data[445 % IN_WIDTH] : pong_storage_data_816 ^ i_input_data[445 % IN_WIDTH];
                504 / IN_WIDTH: pong_storage_data_816 <= (fillup_transition == 1'b1) ? i_input_data[504 % IN_WIDTH] : pong_storage_data_816 ^ i_input_data[504 % IN_WIDTH];
                677 / IN_WIDTH: pong_storage_data_816 <= (fillup_transition == 1'b1) ? i_input_data[677 % IN_WIDTH] : pong_storage_data_816 ^ i_input_data[677 % IN_WIDTH];
                1149 / IN_WIDTH: pong_storage_data_816 <= (fillup_transition == 1'b1) ? i_input_data[1149 % IN_WIDTH] : pong_storage_data_816 ^ i_input_data[1149 % IN_WIDTH];
                default: pong_storage_data_816 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_816;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_816 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_816;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_816 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_816;
            end
        end
    end
end

logic ping_storage_data_817;
logic pong_storage_data_817;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_817 <= 1'b0;
        pong_storage_data_817 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                37 / IN_WIDTH: ping_storage_data_817 <= (fillup_transition == 1'b1) ? i_input_data[37 % IN_WIDTH] : ping_storage_data_817 ^ i_input_data[37 % IN_WIDTH];
                446 / IN_WIDTH: ping_storage_data_817 <= (fillup_transition == 1'b1) ? i_input_data[446 % IN_WIDTH] : ping_storage_data_817 ^ i_input_data[446 % IN_WIDTH];
                505 / IN_WIDTH: ping_storage_data_817 <= (fillup_transition == 1'b1) ? i_input_data[505 % IN_WIDTH] : ping_storage_data_817 ^ i_input_data[505 % IN_WIDTH];
                678 / IN_WIDTH: ping_storage_data_817 <= (fillup_transition == 1'b1) ? i_input_data[678 % IN_WIDTH] : ping_storage_data_817 ^ i_input_data[678 % IN_WIDTH];
                1150 / IN_WIDTH: ping_storage_data_817 <= (fillup_transition == 1'b1) ? i_input_data[1150 % IN_WIDTH] : ping_storage_data_817 ^ i_input_data[1150 % IN_WIDTH];
                default: ping_storage_data_817 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_817;
                endcase
            end else begin
                case (input_count)
                37 / IN_WIDTH: pong_storage_data_817 <= (fillup_transition == 1'b1) ? i_input_data[37 % IN_WIDTH] : pong_storage_data_817 ^ i_input_data[37 % IN_WIDTH];
                446 / IN_WIDTH: pong_storage_data_817 <= (fillup_transition == 1'b1) ? i_input_data[446 % IN_WIDTH] : pong_storage_data_817 ^ i_input_data[446 % IN_WIDTH];
                505 / IN_WIDTH: pong_storage_data_817 <= (fillup_transition == 1'b1) ? i_input_data[505 % IN_WIDTH] : pong_storage_data_817 ^ i_input_data[505 % IN_WIDTH];
                678 / IN_WIDTH: pong_storage_data_817 <= (fillup_transition == 1'b1) ? i_input_data[678 % IN_WIDTH] : pong_storage_data_817 ^ i_input_data[678 % IN_WIDTH];
                1150 / IN_WIDTH: pong_storage_data_817 <= (fillup_transition == 1'b1) ? i_input_data[1150 % IN_WIDTH] : pong_storage_data_817 ^ i_input_data[1150 % IN_WIDTH];
                default: pong_storage_data_817 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_817;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_817 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_817;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_817 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_817;
            end
        end
    end
end

logic ping_storage_data_818;
logic pong_storage_data_818;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_818 <= 1'b0;
        pong_storage_data_818 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                38 / IN_WIDTH: ping_storage_data_818 <= (fillup_transition == 1'b1) ? i_input_data[38 % IN_WIDTH] : ping_storage_data_818 ^ i_input_data[38 % IN_WIDTH];
                447 / IN_WIDTH: ping_storage_data_818 <= (fillup_transition == 1'b1) ? i_input_data[447 % IN_WIDTH] : ping_storage_data_818 ^ i_input_data[447 % IN_WIDTH];
                506 / IN_WIDTH: ping_storage_data_818 <= (fillup_transition == 1'b1) ? i_input_data[506 % IN_WIDTH] : ping_storage_data_818 ^ i_input_data[506 % IN_WIDTH];
                679 / IN_WIDTH: ping_storage_data_818 <= (fillup_transition == 1'b1) ? i_input_data[679 % IN_WIDTH] : ping_storage_data_818 ^ i_input_data[679 % IN_WIDTH];
                1151 / IN_WIDTH: ping_storage_data_818 <= (fillup_transition == 1'b1) ? i_input_data[1151 % IN_WIDTH] : ping_storage_data_818 ^ i_input_data[1151 % IN_WIDTH];
                default: ping_storage_data_818 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_818;
                endcase
            end else begin
                case (input_count)
                38 / IN_WIDTH: pong_storage_data_818 <= (fillup_transition == 1'b1) ? i_input_data[38 % IN_WIDTH] : pong_storage_data_818 ^ i_input_data[38 % IN_WIDTH];
                447 / IN_WIDTH: pong_storage_data_818 <= (fillup_transition == 1'b1) ? i_input_data[447 % IN_WIDTH] : pong_storage_data_818 ^ i_input_data[447 % IN_WIDTH];
                506 / IN_WIDTH: pong_storage_data_818 <= (fillup_transition == 1'b1) ? i_input_data[506 % IN_WIDTH] : pong_storage_data_818 ^ i_input_data[506 % IN_WIDTH];
                679 / IN_WIDTH: pong_storage_data_818 <= (fillup_transition == 1'b1) ? i_input_data[679 % IN_WIDTH] : pong_storage_data_818 ^ i_input_data[679 % IN_WIDTH];
                1151 / IN_WIDTH: pong_storage_data_818 <= (fillup_transition == 1'b1) ? i_input_data[1151 % IN_WIDTH] : pong_storage_data_818 ^ i_input_data[1151 % IN_WIDTH];
                default: pong_storage_data_818 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_818;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_818 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_818;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_818 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_818;
            end
        end
    end
end

logic ping_storage_data_819;
logic pong_storage_data_819;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_819 <= 1'b0;
        pong_storage_data_819 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                39 / IN_WIDTH: ping_storage_data_819 <= (fillup_transition == 1'b1) ? i_input_data[39 % IN_WIDTH] : ping_storage_data_819 ^ i_input_data[39 % IN_WIDTH];
                448 / IN_WIDTH: ping_storage_data_819 <= (fillup_transition == 1'b1) ? i_input_data[448 % IN_WIDTH] : ping_storage_data_819 ^ i_input_data[448 % IN_WIDTH];
                507 / IN_WIDTH: ping_storage_data_819 <= (fillup_transition == 1'b1) ? i_input_data[507 % IN_WIDTH] : ping_storage_data_819 ^ i_input_data[507 % IN_WIDTH];
                680 / IN_WIDTH: ping_storage_data_819 <= (fillup_transition == 1'b1) ? i_input_data[680 % IN_WIDTH] : ping_storage_data_819 ^ i_input_data[680 % IN_WIDTH];
                1056 / IN_WIDTH: ping_storage_data_819 <= (fillup_transition == 1'b1) ? i_input_data[1056 % IN_WIDTH] : ping_storage_data_819 ^ i_input_data[1056 % IN_WIDTH];
                default: ping_storage_data_819 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_819;
                endcase
            end else begin
                case (input_count)
                39 / IN_WIDTH: pong_storage_data_819 <= (fillup_transition == 1'b1) ? i_input_data[39 % IN_WIDTH] : pong_storage_data_819 ^ i_input_data[39 % IN_WIDTH];
                448 / IN_WIDTH: pong_storage_data_819 <= (fillup_transition == 1'b1) ? i_input_data[448 % IN_WIDTH] : pong_storage_data_819 ^ i_input_data[448 % IN_WIDTH];
                507 / IN_WIDTH: pong_storage_data_819 <= (fillup_transition == 1'b1) ? i_input_data[507 % IN_WIDTH] : pong_storage_data_819 ^ i_input_data[507 % IN_WIDTH];
                680 / IN_WIDTH: pong_storage_data_819 <= (fillup_transition == 1'b1) ? i_input_data[680 % IN_WIDTH] : pong_storage_data_819 ^ i_input_data[680 % IN_WIDTH];
                1056 / IN_WIDTH: pong_storage_data_819 <= (fillup_transition == 1'b1) ? i_input_data[1056 % IN_WIDTH] : pong_storage_data_819 ^ i_input_data[1056 % IN_WIDTH];
                default: pong_storage_data_819 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_819;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_819 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_819;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_819 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_819;
            end
        end
    end
end

logic ping_storage_data_820;
logic pong_storage_data_820;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_820 <= 1'b0;
        pong_storage_data_820 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                40 / IN_WIDTH: ping_storage_data_820 <= (fillup_transition == 1'b1) ? i_input_data[40 % IN_WIDTH] : ping_storage_data_820 ^ i_input_data[40 % IN_WIDTH];
                449 / IN_WIDTH: ping_storage_data_820 <= (fillup_transition == 1'b1) ? i_input_data[449 % IN_WIDTH] : ping_storage_data_820 ^ i_input_data[449 % IN_WIDTH];
                508 / IN_WIDTH: ping_storage_data_820 <= (fillup_transition == 1'b1) ? i_input_data[508 % IN_WIDTH] : ping_storage_data_820 ^ i_input_data[508 % IN_WIDTH];
                681 / IN_WIDTH: ping_storage_data_820 <= (fillup_transition == 1'b1) ? i_input_data[681 % IN_WIDTH] : ping_storage_data_820 ^ i_input_data[681 % IN_WIDTH];
                1057 / IN_WIDTH: ping_storage_data_820 <= (fillup_transition == 1'b1) ? i_input_data[1057 % IN_WIDTH] : ping_storage_data_820 ^ i_input_data[1057 % IN_WIDTH];
                default: ping_storage_data_820 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_820;
                endcase
            end else begin
                case (input_count)
                40 / IN_WIDTH: pong_storage_data_820 <= (fillup_transition == 1'b1) ? i_input_data[40 % IN_WIDTH] : pong_storage_data_820 ^ i_input_data[40 % IN_WIDTH];
                449 / IN_WIDTH: pong_storage_data_820 <= (fillup_transition == 1'b1) ? i_input_data[449 % IN_WIDTH] : pong_storage_data_820 ^ i_input_data[449 % IN_WIDTH];
                508 / IN_WIDTH: pong_storage_data_820 <= (fillup_transition == 1'b1) ? i_input_data[508 % IN_WIDTH] : pong_storage_data_820 ^ i_input_data[508 % IN_WIDTH];
                681 / IN_WIDTH: pong_storage_data_820 <= (fillup_transition == 1'b1) ? i_input_data[681 % IN_WIDTH] : pong_storage_data_820 ^ i_input_data[681 % IN_WIDTH];
                1057 / IN_WIDTH: pong_storage_data_820 <= (fillup_transition == 1'b1) ? i_input_data[1057 % IN_WIDTH] : pong_storage_data_820 ^ i_input_data[1057 % IN_WIDTH];
                default: pong_storage_data_820 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_820;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_820 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_820;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_820 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_820;
            end
        end
    end
end

logic ping_storage_data_821;
logic pong_storage_data_821;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_821 <= 1'b0;
        pong_storage_data_821 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                41 / IN_WIDTH: ping_storage_data_821 <= (fillup_transition == 1'b1) ? i_input_data[41 % IN_WIDTH] : ping_storage_data_821 ^ i_input_data[41 % IN_WIDTH];
                450 / IN_WIDTH: ping_storage_data_821 <= (fillup_transition == 1'b1) ? i_input_data[450 % IN_WIDTH] : ping_storage_data_821 ^ i_input_data[450 % IN_WIDTH];
                509 / IN_WIDTH: ping_storage_data_821 <= (fillup_transition == 1'b1) ? i_input_data[509 % IN_WIDTH] : ping_storage_data_821 ^ i_input_data[509 % IN_WIDTH];
                682 / IN_WIDTH: ping_storage_data_821 <= (fillup_transition == 1'b1) ? i_input_data[682 % IN_WIDTH] : ping_storage_data_821 ^ i_input_data[682 % IN_WIDTH];
                1058 / IN_WIDTH: ping_storage_data_821 <= (fillup_transition == 1'b1) ? i_input_data[1058 % IN_WIDTH] : ping_storage_data_821 ^ i_input_data[1058 % IN_WIDTH];
                default: ping_storage_data_821 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_821;
                endcase
            end else begin
                case (input_count)
                41 / IN_WIDTH: pong_storage_data_821 <= (fillup_transition == 1'b1) ? i_input_data[41 % IN_WIDTH] : pong_storage_data_821 ^ i_input_data[41 % IN_WIDTH];
                450 / IN_WIDTH: pong_storage_data_821 <= (fillup_transition == 1'b1) ? i_input_data[450 % IN_WIDTH] : pong_storage_data_821 ^ i_input_data[450 % IN_WIDTH];
                509 / IN_WIDTH: pong_storage_data_821 <= (fillup_transition == 1'b1) ? i_input_data[509 % IN_WIDTH] : pong_storage_data_821 ^ i_input_data[509 % IN_WIDTH];
                682 / IN_WIDTH: pong_storage_data_821 <= (fillup_transition == 1'b1) ? i_input_data[682 % IN_WIDTH] : pong_storage_data_821 ^ i_input_data[682 % IN_WIDTH];
                1058 / IN_WIDTH: pong_storage_data_821 <= (fillup_transition == 1'b1) ? i_input_data[1058 % IN_WIDTH] : pong_storage_data_821 ^ i_input_data[1058 % IN_WIDTH];
                default: pong_storage_data_821 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_821;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_821 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_821;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_821 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_821;
            end
        end
    end
end

logic ping_storage_data_822;
logic pong_storage_data_822;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_822 <= 1'b0;
        pong_storage_data_822 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                42 / IN_WIDTH: ping_storage_data_822 <= (fillup_transition == 1'b1) ? i_input_data[42 % IN_WIDTH] : ping_storage_data_822 ^ i_input_data[42 % IN_WIDTH];
                451 / IN_WIDTH: ping_storage_data_822 <= (fillup_transition == 1'b1) ? i_input_data[451 % IN_WIDTH] : ping_storage_data_822 ^ i_input_data[451 % IN_WIDTH];
                510 / IN_WIDTH: ping_storage_data_822 <= (fillup_transition == 1'b1) ? i_input_data[510 % IN_WIDTH] : ping_storage_data_822 ^ i_input_data[510 % IN_WIDTH];
                683 / IN_WIDTH: ping_storage_data_822 <= (fillup_transition == 1'b1) ? i_input_data[683 % IN_WIDTH] : ping_storage_data_822 ^ i_input_data[683 % IN_WIDTH];
                1059 / IN_WIDTH: ping_storage_data_822 <= (fillup_transition == 1'b1) ? i_input_data[1059 % IN_WIDTH] : ping_storage_data_822 ^ i_input_data[1059 % IN_WIDTH];
                default: ping_storage_data_822 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_822;
                endcase
            end else begin
                case (input_count)
                42 / IN_WIDTH: pong_storage_data_822 <= (fillup_transition == 1'b1) ? i_input_data[42 % IN_WIDTH] : pong_storage_data_822 ^ i_input_data[42 % IN_WIDTH];
                451 / IN_WIDTH: pong_storage_data_822 <= (fillup_transition == 1'b1) ? i_input_data[451 % IN_WIDTH] : pong_storage_data_822 ^ i_input_data[451 % IN_WIDTH];
                510 / IN_WIDTH: pong_storage_data_822 <= (fillup_transition == 1'b1) ? i_input_data[510 % IN_WIDTH] : pong_storage_data_822 ^ i_input_data[510 % IN_WIDTH];
                683 / IN_WIDTH: pong_storage_data_822 <= (fillup_transition == 1'b1) ? i_input_data[683 % IN_WIDTH] : pong_storage_data_822 ^ i_input_data[683 % IN_WIDTH];
                1059 / IN_WIDTH: pong_storage_data_822 <= (fillup_transition == 1'b1) ? i_input_data[1059 % IN_WIDTH] : pong_storage_data_822 ^ i_input_data[1059 % IN_WIDTH];
                default: pong_storage_data_822 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_822;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_822 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_822;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_822 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_822;
            end
        end
    end
end

logic ping_storage_data_823;
logic pong_storage_data_823;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_823 <= 1'b0;
        pong_storage_data_823 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                43 / IN_WIDTH: ping_storage_data_823 <= (fillup_transition == 1'b1) ? i_input_data[43 % IN_WIDTH] : ping_storage_data_823 ^ i_input_data[43 % IN_WIDTH];
                452 / IN_WIDTH: ping_storage_data_823 <= (fillup_transition == 1'b1) ? i_input_data[452 % IN_WIDTH] : ping_storage_data_823 ^ i_input_data[452 % IN_WIDTH];
                511 / IN_WIDTH: ping_storage_data_823 <= (fillup_transition == 1'b1) ? i_input_data[511 % IN_WIDTH] : ping_storage_data_823 ^ i_input_data[511 % IN_WIDTH];
                684 / IN_WIDTH: ping_storage_data_823 <= (fillup_transition == 1'b1) ? i_input_data[684 % IN_WIDTH] : ping_storage_data_823 ^ i_input_data[684 % IN_WIDTH];
                1060 / IN_WIDTH: ping_storage_data_823 <= (fillup_transition == 1'b1) ? i_input_data[1060 % IN_WIDTH] : ping_storage_data_823 ^ i_input_data[1060 % IN_WIDTH];
                default: ping_storage_data_823 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_823;
                endcase
            end else begin
                case (input_count)
                43 / IN_WIDTH: pong_storage_data_823 <= (fillup_transition == 1'b1) ? i_input_data[43 % IN_WIDTH] : pong_storage_data_823 ^ i_input_data[43 % IN_WIDTH];
                452 / IN_WIDTH: pong_storage_data_823 <= (fillup_transition == 1'b1) ? i_input_data[452 % IN_WIDTH] : pong_storage_data_823 ^ i_input_data[452 % IN_WIDTH];
                511 / IN_WIDTH: pong_storage_data_823 <= (fillup_transition == 1'b1) ? i_input_data[511 % IN_WIDTH] : pong_storage_data_823 ^ i_input_data[511 % IN_WIDTH];
                684 / IN_WIDTH: pong_storage_data_823 <= (fillup_transition == 1'b1) ? i_input_data[684 % IN_WIDTH] : pong_storage_data_823 ^ i_input_data[684 % IN_WIDTH];
                1060 / IN_WIDTH: pong_storage_data_823 <= (fillup_transition == 1'b1) ? i_input_data[1060 % IN_WIDTH] : pong_storage_data_823 ^ i_input_data[1060 % IN_WIDTH];
                default: pong_storage_data_823 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_823;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_823 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_823;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_823 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_823;
            end
        end
    end
end

logic ping_storage_data_824;
logic pong_storage_data_824;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_824 <= 1'b0;
        pong_storage_data_824 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                44 / IN_WIDTH: ping_storage_data_824 <= (fillup_transition == 1'b1) ? i_input_data[44 % IN_WIDTH] : ping_storage_data_824 ^ i_input_data[44 % IN_WIDTH];
                453 / IN_WIDTH: ping_storage_data_824 <= (fillup_transition == 1'b1) ? i_input_data[453 % IN_WIDTH] : ping_storage_data_824 ^ i_input_data[453 % IN_WIDTH];
                512 / IN_WIDTH: ping_storage_data_824 <= (fillup_transition == 1'b1) ? i_input_data[512 % IN_WIDTH] : ping_storage_data_824 ^ i_input_data[512 % IN_WIDTH];
                685 / IN_WIDTH: ping_storage_data_824 <= (fillup_transition == 1'b1) ? i_input_data[685 % IN_WIDTH] : ping_storage_data_824 ^ i_input_data[685 % IN_WIDTH];
                1061 / IN_WIDTH: ping_storage_data_824 <= (fillup_transition == 1'b1) ? i_input_data[1061 % IN_WIDTH] : ping_storage_data_824 ^ i_input_data[1061 % IN_WIDTH];
                default: ping_storage_data_824 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_824;
                endcase
            end else begin
                case (input_count)
                44 / IN_WIDTH: pong_storage_data_824 <= (fillup_transition == 1'b1) ? i_input_data[44 % IN_WIDTH] : pong_storage_data_824 ^ i_input_data[44 % IN_WIDTH];
                453 / IN_WIDTH: pong_storage_data_824 <= (fillup_transition == 1'b1) ? i_input_data[453 % IN_WIDTH] : pong_storage_data_824 ^ i_input_data[453 % IN_WIDTH];
                512 / IN_WIDTH: pong_storage_data_824 <= (fillup_transition == 1'b1) ? i_input_data[512 % IN_WIDTH] : pong_storage_data_824 ^ i_input_data[512 % IN_WIDTH];
                685 / IN_WIDTH: pong_storage_data_824 <= (fillup_transition == 1'b1) ? i_input_data[685 % IN_WIDTH] : pong_storage_data_824 ^ i_input_data[685 % IN_WIDTH];
                1061 / IN_WIDTH: pong_storage_data_824 <= (fillup_transition == 1'b1) ? i_input_data[1061 % IN_WIDTH] : pong_storage_data_824 ^ i_input_data[1061 % IN_WIDTH];
                default: pong_storage_data_824 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_824;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_824 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_824;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_824 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_824;
            end
        end
    end
end

logic ping_storage_data_825;
logic pong_storage_data_825;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_825 <= 1'b0;
        pong_storage_data_825 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                45 / IN_WIDTH: ping_storage_data_825 <= (fillup_transition == 1'b1) ? i_input_data[45 % IN_WIDTH] : ping_storage_data_825 ^ i_input_data[45 % IN_WIDTH];
                454 / IN_WIDTH: ping_storage_data_825 <= (fillup_transition == 1'b1) ? i_input_data[454 % IN_WIDTH] : ping_storage_data_825 ^ i_input_data[454 % IN_WIDTH];
                513 / IN_WIDTH: ping_storage_data_825 <= (fillup_transition == 1'b1) ? i_input_data[513 % IN_WIDTH] : ping_storage_data_825 ^ i_input_data[513 % IN_WIDTH];
                686 / IN_WIDTH: ping_storage_data_825 <= (fillup_transition == 1'b1) ? i_input_data[686 % IN_WIDTH] : ping_storage_data_825 ^ i_input_data[686 % IN_WIDTH];
                1062 / IN_WIDTH: ping_storage_data_825 <= (fillup_transition == 1'b1) ? i_input_data[1062 % IN_WIDTH] : ping_storage_data_825 ^ i_input_data[1062 % IN_WIDTH];
                default: ping_storage_data_825 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_825;
                endcase
            end else begin
                case (input_count)
                45 / IN_WIDTH: pong_storage_data_825 <= (fillup_transition == 1'b1) ? i_input_data[45 % IN_WIDTH] : pong_storage_data_825 ^ i_input_data[45 % IN_WIDTH];
                454 / IN_WIDTH: pong_storage_data_825 <= (fillup_transition == 1'b1) ? i_input_data[454 % IN_WIDTH] : pong_storage_data_825 ^ i_input_data[454 % IN_WIDTH];
                513 / IN_WIDTH: pong_storage_data_825 <= (fillup_transition == 1'b1) ? i_input_data[513 % IN_WIDTH] : pong_storage_data_825 ^ i_input_data[513 % IN_WIDTH];
                686 / IN_WIDTH: pong_storage_data_825 <= (fillup_transition == 1'b1) ? i_input_data[686 % IN_WIDTH] : pong_storage_data_825 ^ i_input_data[686 % IN_WIDTH];
                1062 / IN_WIDTH: pong_storage_data_825 <= (fillup_transition == 1'b1) ? i_input_data[1062 % IN_WIDTH] : pong_storage_data_825 ^ i_input_data[1062 % IN_WIDTH];
                default: pong_storage_data_825 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_825;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_825 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_825;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_825 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_825;
            end
        end
    end
end

logic ping_storage_data_826;
logic pong_storage_data_826;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_826 <= 1'b0;
        pong_storage_data_826 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                46 / IN_WIDTH: ping_storage_data_826 <= (fillup_transition == 1'b1) ? i_input_data[46 % IN_WIDTH] : ping_storage_data_826 ^ i_input_data[46 % IN_WIDTH];
                455 / IN_WIDTH: ping_storage_data_826 <= (fillup_transition == 1'b1) ? i_input_data[455 % IN_WIDTH] : ping_storage_data_826 ^ i_input_data[455 % IN_WIDTH];
                514 / IN_WIDTH: ping_storage_data_826 <= (fillup_transition == 1'b1) ? i_input_data[514 % IN_WIDTH] : ping_storage_data_826 ^ i_input_data[514 % IN_WIDTH];
                687 / IN_WIDTH: ping_storage_data_826 <= (fillup_transition == 1'b1) ? i_input_data[687 % IN_WIDTH] : ping_storage_data_826 ^ i_input_data[687 % IN_WIDTH];
                1063 / IN_WIDTH: ping_storage_data_826 <= (fillup_transition == 1'b1) ? i_input_data[1063 % IN_WIDTH] : ping_storage_data_826 ^ i_input_data[1063 % IN_WIDTH];
                default: ping_storage_data_826 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_826;
                endcase
            end else begin
                case (input_count)
                46 / IN_WIDTH: pong_storage_data_826 <= (fillup_transition == 1'b1) ? i_input_data[46 % IN_WIDTH] : pong_storage_data_826 ^ i_input_data[46 % IN_WIDTH];
                455 / IN_WIDTH: pong_storage_data_826 <= (fillup_transition == 1'b1) ? i_input_data[455 % IN_WIDTH] : pong_storage_data_826 ^ i_input_data[455 % IN_WIDTH];
                514 / IN_WIDTH: pong_storage_data_826 <= (fillup_transition == 1'b1) ? i_input_data[514 % IN_WIDTH] : pong_storage_data_826 ^ i_input_data[514 % IN_WIDTH];
                687 / IN_WIDTH: pong_storage_data_826 <= (fillup_transition == 1'b1) ? i_input_data[687 % IN_WIDTH] : pong_storage_data_826 ^ i_input_data[687 % IN_WIDTH];
                1063 / IN_WIDTH: pong_storage_data_826 <= (fillup_transition == 1'b1) ? i_input_data[1063 % IN_WIDTH] : pong_storage_data_826 ^ i_input_data[1063 % IN_WIDTH];
                default: pong_storage_data_826 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_826;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_826 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_826;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_826 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_826;
            end
        end
    end
end

logic ping_storage_data_827;
logic pong_storage_data_827;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_827 <= 1'b0;
        pong_storage_data_827 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                47 / IN_WIDTH: ping_storage_data_827 <= (fillup_transition == 1'b1) ? i_input_data[47 % IN_WIDTH] : ping_storage_data_827 ^ i_input_data[47 % IN_WIDTH];
                456 / IN_WIDTH: ping_storage_data_827 <= (fillup_transition == 1'b1) ? i_input_data[456 % IN_WIDTH] : ping_storage_data_827 ^ i_input_data[456 % IN_WIDTH];
                515 / IN_WIDTH: ping_storage_data_827 <= (fillup_transition == 1'b1) ? i_input_data[515 % IN_WIDTH] : ping_storage_data_827 ^ i_input_data[515 % IN_WIDTH];
                688 / IN_WIDTH: ping_storage_data_827 <= (fillup_transition == 1'b1) ? i_input_data[688 % IN_WIDTH] : ping_storage_data_827 ^ i_input_data[688 % IN_WIDTH];
                1064 / IN_WIDTH: ping_storage_data_827 <= (fillup_transition == 1'b1) ? i_input_data[1064 % IN_WIDTH] : ping_storage_data_827 ^ i_input_data[1064 % IN_WIDTH];
                default: ping_storage_data_827 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_827;
                endcase
            end else begin
                case (input_count)
                47 / IN_WIDTH: pong_storage_data_827 <= (fillup_transition == 1'b1) ? i_input_data[47 % IN_WIDTH] : pong_storage_data_827 ^ i_input_data[47 % IN_WIDTH];
                456 / IN_WIDTH: pong_storage_data_827 <= (fillup_transition == 1'b1) ? i_input_data[456 % IN_WIDTH] : pong_storage_data_827 ^ i_input_data[456 % IN_WIDTH];
                515 / IN_WIDTH: pong_storage_data_827 <= (fillup_transition == 1'b1) ? i_input_data[515 % IN_WIDTH] : pong_storage_data_827 ^ i_input_data[515 % IN_WIDTH];
                688 / IN_WIDTH: pong_storage_data_827 <= (fillup_transition == 1'b1) ? i_input_data[688 % IN_WIDTH] : pong_storage_data_827 ^ i_input_data[688 % IN_WIDTH];
                1064 / IN_WIDTH: pong_storage_data_827 <= (fillup_transition == 1'b1) ? i_input_data[1064 % IN_WIDTH] : pong_storage_data_827 ^ i_input_data[1064 % IN_WIDTH];
                default: pong_storage_data_827 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_827;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_827 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_827;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_827 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_827;
            end
        end
    end
end

logic ping_storage_data_828;
logic pong_storage_data_828;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_828 <= 1'b0;
        pong_storage_data_828 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                48 / IN_WIDTH: ping_storage_data_828 <= (fillup_transition == 1'b1) ? i_input_data[48 % IN_WIDTH] : ping_storage_data_828 ^ i_input_data[48 % IN_WIDTH];
                457 / IN_WIDTH: ping_storage_data_828 <= (fillup_transition == 1'b1) ? i_input_data[457 % IN_WIDTH] : ping_storage_data_828 ^ i_input_data[457 % IN_WIDTH];
                516 / IN_WIDTH: ping_storage_data_828 <= (fillup_transition == 1'b1) ? i_input_data[516 % IN_WIDTH] : ping_storage_data_828 ^ i_input_data[516 % IN_WIDTH];
                689 / IN_WIDTH: ping_storage_data_828 <= (fillup_transition == 1'b1) ? i_input_data[689 % IN_WIDTH] : ping_storage_data_828 ^ i_input_data[689 % IN_WIDTH];
                1065 / IN_WIDTH: ping_storage_data_828 <= (fillup_transition == 1'b1) ? i_input_data[1065 % IN_WIDTH] : ping_storage_data_828 ^ i_input_data[1065 % IN_WIDTH];
                default: ping_storage_data_828 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_828;
                endcase
            end else begin
                case (input_count)
                48 / IN_WIDTH: pong_storage_data_828 <= (fillup_transition == 1'b1) ? i_input_data[48 % IN_WIDTH] : pong_storage_data_828 ^ i_input_data[48 % IN_WIDTH];
                457 / IN_WIDTH: pong_storage_data_828 <= (fillup_transition == 1'b1) ? i_input_data[457 % IN_WIDTH] : pong_storage_data_828 ^ i_input_data[457 % IN_WIDTH];
                516 / IN_WIDTH: pong_storage_data_828 <= (fillup_transition == 1'b1) ? i_input_data[516 % IN_WIDTH] : pong_storage_data_828 ^ i_input_data[516 % IN_WIDTH];
                689 / IN_WIDTH: pong_storage_data_828 <= (fillup_transition == 1'b1) ? i_input_data[689 % IN_WIDTH] : pong_storage_data_828 ^ i_input_data[689 % IN_WIDTH];
                1065 / IN_WIDTH: pong_storage_data_828 <= (fillup_transition == 1'b1) ? i_input_data[1065 % IN_WIDTH] : pong_storage_data_828 ^ i_input_data[1065 % IN_WIDTH];
                default: pong_storage_data_828 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_828;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_828 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_828;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_828 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_828;
            end
        end
    end
end

logic ping_storage_data_829;
logic pong_storage_data_829;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_829 <= 1'b0;
        pong_storage_data_829 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                49 / IN_WIDTH: ping_storage_data_829 <= (fillup_transition == 1'b1) ? i_input_data[49 % IN_WIDTH] : ping_storage_data_829 ^ i_input_data[49 % IN_WIDTH];
                458 / IN_WIDTH: ping_storage_data_829 <= (fillup_transition == 1'b1) ? i_input_data[458 % IN_WIDTH] : ping_storage_data_829 ^ i_input_data[458 % IN_WIDTH];
                517 / IN_WIDTH: ping_storage_data_829 <= (fillup_transition == 1'b1) ? i_input_data[517 % IN_WIDTH] : ping_storage_data_829 ^ i_input_data[517 % IN_WIDTH];
                690 / IN_WIDTH: ping_storage_data_829 <= (fillup_transition == 1'b1) ? i_input_data[690 % IN_WIDTH] : ping_storage_data_829 ^ i_input_data[690 % IN_WIDTH];
                1066 / IN_WIDTH: ping_storage_data_829 <= (fillup_transition == 1'b1) ? i_input_data[1066 % IN_WIDTH] : ping_storage_data_829 ^ i_input_data[1066 % IN_WIDTH];
                default: ping_storage_data_829 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_829;
                endcase
            end else begin
                case (input_count)
                49 / IN_WIDTH: pong_storage_data_829 <= (fillup_transition == 1'b1) ? i_input_data[49 % IN_WIDTH] : pong_storage_data_829 ^ i_input_data[49 % IN_WIDTH];
                458 / IN_WIDTH: pong_storage_data_829 <= (fillup_transition == 1'b1) ? i_input_data[458 % IN_WIDTH] : pong_storage_data_829 ^ i_input_data[458 % IN_WIDTH];
                517 / IN_WIDTH: pong_storage_data_829 <= (fillup_transition == 1'b1) ? i_input_data[517 % IN_WIDTH] : pong_storage_data_829 ^ i_input_data[517 % IN_WIDTH];
                690 / IN_WIDTH: pong_storage_data_829 <= (fillup_transition == 1'b1) ? i_input_data[690 % IN_WIDTH] : pong_storage_data_829 ^ i_input_data[690 % IN_WIDTH];
                1066 / IN_WIDTH: pong_storage_data_829 <= (fillup_transition == 1'b1) ? i_input_data[1066 % IN_WIDTH] : pong_storage_data_829 ^ i_input_data[1066 % IN_WIDTH];
                default: pong_storage_data_829 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_829;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_829 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_829;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_829 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_829;
            end
        end
    end
end

logic ping_storage_data_830;
logic pong_storage_data_830;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_830 <= 1'b0;
        pong_storage_data_830 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                50 / IN_WIDTH: ping_storage_data_830 <= (fillup_transition == 1'b1) ? i_input_data[50 % IN_WIDTH] : ping_storage_data_830 ^ i_input_data[50 % IN_WIDTH];
                459 / IN_WIDTH: ping_storage_data_830 <= (fillup_transition == 1'b1) ? i_input_data[459 % IN_WIDTH] : ping_storage_data_830 ^ i_input_data[459 % IN_WIDTH];
                518 / IN_WIDTH: ping_storage_data_830 <= (fillup_transition == 1'b1) ? i_input_data[518 % IN_WIDTH] : ping_storage_data_830 ^ i_input_data[518 % IN_WIDTH];
                691 / IN_WIDTH: ping_storage_data_830 <= (fillup_transition == 1'b1) ? i_input_data[691 % IN_WIDTH] : ping_storage_data_830 ^ i_input_data[691 % IN_WIDTH];
                1067 / IN_WIDTH: ping_storage_data_830 <= (fillup_transition == 1'b1) ? i_input_data[1067 % IN_WIDTH] : ping_storage_data_830 ^ i_input_data[1067 % IN_WIDTH];
                default: ping_storage_data_830 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_830;
                endcase
            end else begin
                case (input_count)
                50 / IN_WIDTH: pong_storage_data_830 <= (fillup_transition == 1'b1) ? i_input_data[50 % IN_WIDTH] : pong_storage_data_830 ^ i_input_data[50 % IN_WIDTH];
                459 / IN_WIDTH: pong_storage_data_830 <= (fillup_transition == 1'b1) ? i_input_data[459 % IN_WIDTH] : pong_storage_data_830 ^ i_input_data[459 % IN_WIDTH];
                518 / IN_WIDTH: pong_storage_data_830 <= (fillup_transition == 1'b1) ? i_input_data[518 % IN_WIDTH] : pong_storage_data_830 ^ i_input_data[518 % IN_WIDTH];
                691 / IN_WIDTH: pong_storage_data_830 <= (fillup_transition == 1'b1) ? i_input_data[691 % IN_WIDTH] : pong_storage_data_830 ^ i_input_data[691 % IN_WIDTH];
                1067 / IN_WIDTH: pong_storage_data_830 <= (fillup_transition == 1'b1) ? i_input_data[1067 % IN_WIDTH] : pong_storage_data_830 ^ i_input_data[1067 % IN_WIDTH];
                default: pong_storage_data_830 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_830;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_830 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_830;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_830 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_830;
            end
        end
    end
end

logic ping_storage_data_831;
logic pong_storage_data_831;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_831 <= 1'b0;
        pong_storage_data_831 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                51 / IN_WIDTH: ping_storage_data_831 <= (fillup_transition == 1'b1) ? i_input_data[51 % IN_WIDTH] : ping_storage_data_831 ^ i_input_data[51 % IN_WIDTH];
                460 / IN_WIDTH: ping_storage_data_831 <= (fillup_transition == 1'b1) ? i_input_data[460 % IN_WIDTH] : ping_storage_data_831 ^ i_input_data[460 % IN_WIDTH];
                519 / IN_WIDTH: ping_storage_data_831 <= (fillup_transition == 1'b1) ? i_input_data[519 % IN_WIDTH] : ping_storage_data_831 ^ i_input_data[519 % IN_WIDTH];
                692 / IN_WIDTH: ping_storage_data_831 <= (fillup_transition == 1'b1) ? i_input_data[692 % IN_WIDTH] : ping_storage_data_831 ^ i_input_data[692 % IN_WIDTH];
                1068 / IN_WIDTH: ping_storage_data_831 <= (fillup_transition == 1'b1) ? i_input_data[1068 % IN_WIDTH] : ping_storage_data_831 ^ i_input_data[1068 % IN_WIDTH];
                default: ping_storage_data_831 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_831;
                endcase
            end else begin
                case (input_count)
                51 / IN_WIDTH: pong_storage_data_831 <= (fillup_transition == 1'b1) ? i_input_data[51 % IN_WIDTH] : pong_storage_data_831 ^ i_input_data[51 % IN_WIDTH];
                460 / IN_WIDTH: pong_storage_data_831 <= (fillup_transition == 1'b1) ? i_input_data[460 % IN_WIDTH] : pong_storage_data_831 ^ i_input_data[460 % IN_WIDTH];
                519 / IN_WIDTH: pong_storage_data_831 <= (fillup_transition == 1'b1) ? i_input_data[519 % IN_WIDTH] : pong_storage_data_831 ^ i_input_data[519 % IN_WIDTH];
                692 / IN_WIDTH: pong_storage_data_831 <= (fillup_transition == 1'b1) ? i_input_data[692 % IN_WIDTH] : pong_storage_data_831 ^ i_input_data[692 % IN_WIDTH];
                1068 / IN_WIDTH: pong_storage_data_831 <= (fillup_transition == 1'b1) ? i_input_data[1068 % IN_WIDTH] : pong_storage_data_831 ^ i_input_data[1068 % IN_WIDTH];
                default: pong_storage_data_831 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_831;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_831 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_831;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_831 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_831;
            end
        end
    end
end

logic ping_storage_data_832;
logic pong_storage_data_832;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_832 <= 1'b0;
        pong_storage_data_832 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                52 / IN_WIDTH: ping_storage_data_832 <= (fillup_transition == 1'b1) ? i_input_data[52 % IN_WIDTH] : ping_storage_data_832 ^ i_input_data[52 % IN_WIDTH];
                461 / IN_WIDTH: ping_storage_data_832 <= (fillup_transition == 1'b1) ? i_input_data[461 % IN_WIDTH] : ping_storage_data_832 ^ i_input_data[461 % IN_WIDTH];
                520 / IN_WIDTH: ping_storage_data_832 <= (fillup_transition == 1'b1) ? i_input_data[520 % IN_WIDTH] : ping_storage_data_832 ^ i_input_data[520 % IN_WIDTH];
                693 / IN_WIDTH: ping_storage_data_832 <= (fillup_transition == 1'b1) ? i_input_data[693 % IN_WIDTH] : ping_storage_data_832 ^ i_input_data[693 % IN_WIDTH];
                1069 / IN_WIDTH: ping_storage_data_832 <= (fillup_transition == 1'b1) ? i_input_data[1069 % IN_WIDTH] : ping_storage_data_832 ^ i_input_data[1069 % IN_WIDTH];
                default: ping_storage_data_832 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_832;
                endcase
            end else begin
                case (input_count)
                52 / IN_WIDTH: pong_storage_data_832 <= (fillup_transition == 1'b1) ? i_input_data[52 % IN_WIDTH] : pong_storage_data_832 ^ i_input_data[52 % IN_WIDTH];
                461 / IN_WIDTH: pong_storage_data_832 <= (fillup_transition == 1'b1) ? i_input_data[461 % IN_WIDTH] : pong_storage_data_832 ^ i_input_data[461 % IN_WIDTH];
                520 / IN_WIDTH: pong_storage_data_832 <= (fillup_transition == 1'b1) ? i_input_data[520 % IN_WIDTH] : pong_storage_data_832 ^ i_input_data[520 % IN_WIDTH];
                693 / IN_WIDTH: pong_storage_data_832 <= (fillup_transition == 1'b1) ? i_input_data[693 % IN_WIDTH] : pong_storage_data_832 ^ i_input_data[693 % IN_WIDTH];
                1069 / IN_WIDTH: pong_storage_data_832 <= (fillup_transition == 1'b1) ? i_input_data[1069 % IN_WIDTH] : pong_storage_data_832 ^ i_input_data[1069 % IN_WIDTH];
                default: pong_storage_data_832 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_832;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_832 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_832;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_832 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_832;
            end
        end
    end
end

logic ping_storage_data_833;
logic pong_storage_data_833;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_833 <= 1'b0;
        pong_storage_data_833 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                53 / IN_WIDTH: ping_storage_data_833 <= (fillup_transition == 1'b1) ? i_input_data[53 % IN_WIDTH] : ping_storage_data_833 ^ i_input_data[53 % IN_WIDTH];
                462 / IN_WIDTH: ping_storage_data_833 <= (fillup_transition == 1'b1) ? i_input_data[462 % IN_WIDTH] : ping_storage_data_833 ^ i_input_data[462 % IN_WIDTH];
                521 / IN_WIDTH: ping_storage_data_833 <= (fillup_transition == 1'b1) ? i_input_data[521 % IN_WIDTH] : ping_storage_data_833 ^ i_input_data[521 % IN_WIDTH];
                694 / IN_WIDTH: ping_storage_data_833 <= (fillup_transition == 1'b1) ? i_input_data[694 % IN_WIDTH] : ping_storage_data_833 ^ i_input_data[694 % IN_WIDTH];
                1070 / IN_WIDTH: ping_storage_data_833 <= (fillup_transition == 1'b1) ? i_input_data[1070 % IN_WIDTH] : ping_storage_data_833 ^ i_input_data[1070 % IN_WIDTH];
                default: ping_storage_data_833 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_833;
                endcase
            end else begin
                case (input_count)
                53 / IN_WIDTH: pong_storage_data_833 <= (fillup_transition == 1'b1) ? i_input_data[53 % IN_WIDTH] : pong_storage_data_833 ^ i_input_data[53 % IN_WIDTH];
                462 / IN_WIDTH: pong_storage_data_833 <= (fillup_transition == 1'b1) ? i_input_data[462 % IN_WIDTH] : pong_storage_data_833 ^ i_input_data[462 % IN_WIDTH];
                521 / IN_WIDTH: pong_storage_data_833 <= (fillup_transition == 1'b1) ? i_input_data[521 % IN_WIDTH] : pong_storage_data_833 ^ i_input_data[521 % IN_WIDTH];
                694 / IN_WIDTH: pong_storage_data_833 <= (fillup_transition == 1'b1) ? i_input_data[694 % IN_WIDTH] : pong_storage_data_833 ^ i_input_data[694 % IN_WIDTH];
                1070 / IN_WIDTH: pong_storage_data_833 <= (fillup_transition == 1'b1) ? i_input_data[1070 % IN_WIDTH] : pong_storage_data_833 ^ i_input_data[1070 % IN_WIDTH];
                default: pong_storage_data_833 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_833;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_833 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_833;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_833 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_833;
            end
        end
    end
end

logic ping_storage_data_834;
logic pong_storage_data_834;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_834 <= 1'b0;
        pong_storage_data_834 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                54 / IN_WIDTH: ping_storage_data_834 <= (fillup_transition == 1'b1) ? i_input_data[54 % IN_WIDTH] : ping_storage_data_834 ^ i_input_data[54 % IN_WIDTH];
                463 / IN_WIDTH: ping_storage_data_834 <= (fillup_transition == 1'b1) ? i_input_data[463 % IN_WIDTH] : ping_storage_data_834 ^ i_input_data[463 % IN_WIDTH];
                522 / IN_WIDTH: ping_storage_data_834 <= (fillup_transition == 1'b1) ? i_input_data[522 % IN_WIDTH] : ping_storage_data_834 ^ i_input_data[522 % IN_WIDTH];
                695 / IN_WIDTH: ping_storage_data_834 <= (fillup_transition == 1'b1) ? i_input_data[695 % IN_WIDTH] : ping_storage_data_834 ^ i_input_data[695 % IN_WIDTH];
                1071 / IN_WIDTH: ping_storage_data_834 <= (fillup_transition == 1'b1) ? i_input_data[1071 % IN_WIDTH] : ping_storage_data_834 ^ i_input_data[1071 % IN_WIDTH];
                default: ping_storage_data_834 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_834;
                endcase
            end else begin
                case (input_count)
                54 / IN_WIDTH: pong_storage_data_834 <= (fillup_transition == 1'b1) ? i_input_data[54 % IN_WIDTH] : pong_storage_data_834 ^ i_input_data[54 % IN_WIDTH];
                463 / IN_WIDTH: pong_storage_data_834 <= (fillup_transition == 1'b1) ? i_input_data[463 % IN_WIDTH] : pong_storage_data_834 ^ i_input_data[463 % IN_WIDTH];
                522 / IN_WIDTH: pong_storage_data_834 <= (fillup_transition == 1'b1) ? i_input_data[522 % IN_WIDTH] : pong_storage_data_834 ^ i_input_data[522 % IN_WIDTH];
                695 / IN_WIDTH: pong_storage_data_834 <= (fillup_transition == 1'b1) ? i_input_data[695 % IN_WIDTH] : pong_storage_data_834 ^ i_input_data[695 % IN_WIDTH];
                1071 / IN_WIDTH: pong_storage_data_834 <= (fillup_transition == 1'b1) ? i_input_data[1071 % IN_WIDTH] : pong_storage_data_834 ^ i_input_data[1071 % IN_WIDTH];
                default: pong_storage_data_834 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_834;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_834 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_834;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_834 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_834;
            end
        end
    end
end

logic ping_storage_data_835;
logic pong_storage_data_835;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_835 <= 1'b0;
        pong_storage_data_835 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                55 / IN_WIDTH: ping_storage_data_835 <= (fillup_transition == 1'b1) ? i_input_data[55 % IN_WIDTH] : ping_storage_data_835 ^ i_input_data[55 % IN_WIDTH];
                464 / IN_WIDTH: ping_storage_data_835 <= (fillup_transition == 1'b1) ? i_input_data[464 % IN_WIDTH] : ping_storage_data_835 ^ i_input_data[464 % IN_WIDTH];
                523 / IN_WIDTH: ping_storage_data_835 <= (fillup_transition == 1'b1) ? i_input_data[523 % IN_WIDTH] : ping_storage_data_835 ^ i_input_data[523 % IN_WIDTH];
                696 / IN_WIDTH: ping_storage_data_835 <= (fillup_transition == 1'b1) ? i_input_data[696 % IN_WIDTH] : ping_storage_data_835 ^ i_input_data[696 % IN_WIDTH];
                1072 / IN_WIDTH: ping_storage_data_835 <= (fillup_transition == 1'b1) ? i_input_data[1072 % IN_WIDTH] : ping_storage_data_835 ^ i_input_data[1072 % IN_WIDTH];
                default: ping_storage_data_835 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_835;
                endcase
            end else begin
                case (input_count)
                55 / IN_WIDTH: pong_storage_data_835 <= (fillup_transition == 1'b1) ? i_input_data[55 % IN_WIDTH] : pong_storage_data_835 ^ i_input_data[55 % IN_WIDTH];
                464 / IN_WIDTH: pong_storage_data_835 <= (fillup_transition == 1'b1) ? i_input_data[464 % IN_WIDTH] : pong_storage_data_835 ^ i_input_data[464 % IN_WIDTH];
                523 / IN_WIDTH: pong_storage_data_835 <= (fillup_transition == 1'b1) ? i_input_data[523 % IN_WIDTH] : pong_storage_data_835 ^ i_input_data[523 % IN_WIDTH];
                696 / IN_WIDTH: pong_storage_data_835 <= (fillup_transition == 1'b1) ? i_input_data[696 % IN_WIDTH] : pong_storage_data_835 ^ i_input_data[696 % IN_WIDTH];
                1072 / IN_WIDTH: pong_storage_data_835 <= (fillup_transition == 1'b1) ? i_input_data[1072 % IN_WIDTH] : pong_storage_data_835 ^ i_input_data[1072 % IN_WIDTH];
                default: pong_storage_data_835 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_835;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_835 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_835;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_835 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_835;
            end
        end
    end
end

logic ping_storage_data_836;
logic pong_storage_data_836;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_836 <= 1'b0;
        pong_storage_data_836 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                56 / IN_WIDTH: ping_storage_data_836 <= (fillup_transition == 1'b1) ? i_input_data[56 % IN_WIDTH] : ping_storage_data_836 ^ i_input_data[56 % IN_WIDTH];
                465 / IN_WIDTH: ping_storage_data_836 <= (fillup_transition == 1'b1) ? i_input_data[465 % IN_WIDTH] : ping_storage_data_836 ^ i_input_data[465 % IN_WIDTH];
                524 / IN_WIDTH: ping_storage_data_836 <= (fillup_transition == 1'b1) ? i_input_data[524 % IN_WIDTH] : ping_storage_data_836 ^ i_input_data[524 % IN_WIDTH];
                697 / IN_WIDTH: ping_storage_data_836 <= (fillup_transition == 1'b1) ? i_input_data[697 % IN_WIDTH] : ping_storage_data_836 ^ i_input_data[697 % IN_WIDTH];
                1073 / IN_WIDTH: ping_storage_data_836 <= (fillup_transition == 1'b1) ? i_input_data[1073 % IN_WIDTH] : ping_storage_data_836 ^ i_input_data[1073 % IN_WIDTH];
                default: ping_storage_data_836 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_836;
                endcase
            end else begin
                case (input_count)
                56 / IN_WIDTH: pong_storage_data_836 <= (fillup_transition == 1'b1) ? i_input_data[56 % IN_WIDTH] : pong_storage_data_836 ^ i_input_data[56 % IN_WIDTH];
                465 / IN_WIDTH: pong_storage_data_836 <= (fillup_transition == 1'b1) ? i_input_data[465 % IN_WIDTH] : pong_storage_data_836 ^ i_input_data[465 % IN_WIDTH];
                524 / IN_WIDTH: pong_storage_data_836 <= (fillup_transition == 1'b1) ? i_input_data[524 % IN_WIDTH] : pong_storage_data_836 ^ i_input_data[524 % IN_WIDTH];
                697 / IN_WIDTH: pong_storage_data_836 <= (fillup_transition == 1'b1) ? i_input_data[697 % IN_WIDTH] : pong_storage_data_836 ^ i_input_data[697 % IN_WIDTH];
                1073 / IN_WIDTH: pong_storage_data_836 <= (fillup_transition == 1'b1) ? i_input_data[1073 % IN_WIDTH] : pong_storage_data_836 ^ i_input_data[1073 % IN_WIDTH];
                default: pong_storage_data_836 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_836;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_836 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_836;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_836 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_836;
            end
        end
    end
end

logic ping_storage_data_837;
logic pong_storage_data_837;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_837 <= 1'b0;
        pong_storage_data_837 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                57 / IN_WIDTH: ping_storage_data_837 <= (fillup_transition == 1'b1) ? i_input_data[57 % IN_WIDTH] : ping_storage_data_837 ^ i_input_data[57 % IN_WIDTH];
                466 / IN_WIDTH: ping_storage_data_837 <= (fillup_transition == 1'b1) ? i_input_data[466 % IN_WIDTH] : ping_storage_data_837 ^ i_input_data[466 % IN_WIDTH];
                525 / IN_WIDTH: ping_storage_data_837 <= (fillup_transition == 1'b1) ? i_input_data[525 % IN_WIDTH] : ping_storage_data_837 ^ i_input_data[525 % IN_WIDTH];
                698 / IN_WIDTH: ping_storage_data_837 <= (fillup_transition == 1'b1) ? i_input_data[698 % IN_WIDTH] : ping_storage_data_837 ^ i_input_data[698 % IN_WIDTH];
                1074 / IN_WIDTH: ping_storage_data_837 <= (fillup_transition == 1'b1) ? i_input_data[1074 % IN_WIDTH] : ping_storage_data_837 ^ i_input_data[1074 % IN_WIDTH];
                default: ping_storage_data_837 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_837;
                endcase
            end else begin
                case (input_count)
                57 / IN_WIDTH: pong_storage_data_837 <= (fillup_transition == 1'b1) ? i_input_data[57 % IN_WIDTH] : pong_storage_data_837 ^ i_input_data[57 % IN_WIDTH];
                466 / IN_WIDTH: pong_storage_data_837 <= (fillup_transition == 1'b1) ? i_input_data[466 % IN_WIDTH] : pong_storage_data_837 ^ i_input_data[466 % IN_WIDTH];
                525 / IN_WIDTH: pong_storage_data_837 <= (fillup_transition == 1'b1) ? i_input_data[525 % IN_WIDTH] : pong_storage_data_837 ^ i_input_data[525 % IN_WIDTH];
                698 / IN_WIDTH: pong_storage_data_837 <= (fillup_transition == 1'b1) ? i_input_data[698 % IN_WIDTH] : pong_storage_data_837 ^ i_input_data[698 % IN_WIDTH];
                1074 / IN_WIDTH: pong_storage_data_837 <= (fillup_transition == 1'b1) ? i_input_data[1074 % IN_WIDTH] : pong_storage_data_837 ^ i_input_data[1074 % IN_WIDTH];
                default: pong_storage_data_837 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_837;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_837 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_837;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_837 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_837;
            end
        end
    end
end

logic ping_storage_data_838;
logic pong_storage_data_838;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_838 <= 1'b0;
        pong_storage_data_838 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                58 / IN_WIDTH: ping_storage_data_838 <= (fillup_transition == 1'b1) ? i_input_data[58 % IN_WIDTH] : ping_storage_data_838 ^ i_input_data[58 % IN_WIDTH];
                467 / IN_WIDTH: ping_storage_data_838 <= (fillup_transition == 1'b1) ? i_input_data[467 % IN_WIDTH] : ping_storage_data_838 ^ i_input_data[467 % IN_WIDTH];
                526 / IN_WIDTH: ping_storage_data_838 <= (fillup_transition == 1'b1) ? i_input_data[526 % IN_WIDTH] : ping_storage_data_838 ^ i_input_data[526 % IN_WIDTH];
                699 / IN_WIDTH: ping_storage_data_838 <= (fillup_transition == 1'b1) ? i_input_data[699 % IN_WIDTH] : ping_storage_data_838 ^ i_input_data[699 % IN_WIDTH];
                1075 / IN_WIDTH: ping_storage_data_838 <= (fillup_transition == 1'b1) ? i_input_data[1075 % IN_WIDTH] : ping_storage_data_838 ^ i_input_data[1075 % IN_WIDTH];
                default: ping_storage_data_838 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_838;
                endcase
            end else begin
                case (input_count)
                58 / IN_WIDTH: pong_storage_data_838 <= (fillup_transition == 1'b1) ? i_input_data[58 % IN_WIDTH] : pong_storage_data_838 ^ i_input_data[58 % IN_WIDTH];
                467 / IN_WIDTH: pong_storage_data_838 <= (fillup_transition == 1'b1) ? i_input_data[467 % IN_WIDTH] : pong_storage_data_838 ^ i_input_data[467 % IN_WIDTH];
                526 / IN_WIDTH: pong_storage_data_838 <= (fillup_transition == 1'b1) ? i_input_data[526 % IN_WIDTH] : pong_storage_data_838 ^ i_input_data[526 % IN_WIDTH];
                699 / IN_WIDTH: pong_storage_data_838 <= (fillup_transition == 1'b1) ? i_input_data[699 % IN_WIDTH] : pong_storage_data_838 ^ i_input_data[699 % IN_WIDTH];
                1075 / IN_WIDTH: pong_storage_data_838 <= (fillup_transition == 1'b1) ? i_input_data[1075 % IN_WIDTH] : pong_storage_data_838 ^ i_input_data[1075 % IN_WIDTH];
                default: pong_storage_data_838 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_838;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_838 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_838;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_838 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_838;
            end
        end
    end
end

logic ping_storage_data_839;
logic pong_storage_data_839;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_839 <= 1'b0;
        pong_storage_data_839 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                59 / IN_WIDTH: ping_storage_data_839 <= (fillup_transition == 1'b1) ? i_input_data[59 % IN_WIDTH] : ping_storage_data_839 ^ i_input_data[59 % IN_WIDTH];
                468 / IN_WIDTH: ping_storage_data_839 <= (fillup_transition == 1'b1) ? i_input_data[468 % IN_WIDTH] : ping_storage_data_839 ^ i_input_data[468 % IN_WIDTH];
                527 / IN_WIDTH: ping_storage_data_839 <= (fillup_transition == 1'b1) ? i_input_data[527 % IN_WIDTH] : ping_storage_data_839 ^ i_input_data[527 % IN_WIDTH];
                700 / IN_WIDTH: ping_storage_data_839 <= (fillup_transition == 1'b1) ? i_input_data[700 % IN_WIDTH] : ping_storage_data_839 ^ i_input_data[700 % IN_WIDTH];
                1076 / IN_WIDTH: ping_storage_data_839 <= (fillup_transition == 1'b1) ? i_input_data[1076 % IN_WIDTH] : ping_storage_data_839 ^ i_input_data[1076 % IN_WIDTH];
                default: ping_storage_data_839 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_839;
                endcase
            end else begin
                case (input_count)
                59 / IN_WIDTH: pong_storage_data_839 <= (fillup_transition == 1'b1) ? i_input_data[59 % IN_WIDTH] : pong_storage_data_839 ^ i_input_data[59 % IN_WIDTH];
                468 / IN_WIDTH: pong_storage_data_839 <= (fillup_transition == 1'b1) ? i_input_data[468 % IN_WIDTH] : pong_storage_data_839 ^ i_input_data[468 % IN_WIDTH];
                527 / IN_WIDTH: pong_storage_data_839 <= (fillup_transition == 1'b1) ? i_input_data[527 % IN_WIDTH] : pong_storage_data_839 ^ i_input_data[527 % IN_WIDTH];
                700 / IN_WIDTH: pong_storage_data_839 <= (fillup_transition == 1'b1) ? i_input_data[700 % IN_WIDTH] : pong_storage_data_839 ^ i_input_data[700 % IN_WIDTH];
                1076 / IN_WIDTH: pong_storage_data_839 <= (fillup_transition == 1'b1) ? i_input_data[1076 % IN_WIDTH] : pong_storage_data_839 ^ i_input_data[1076 % IN_WIDTH];
                default: pong_storage_data_839 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_839;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_839 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_839;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_839 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_839;
            end
        end
    end
end

logic ping_storage_data_840;
logic pong_storage_data_840;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_840 <= 1'b0;
        pong_storage_data_840 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                60 / IN_WIDTH: ping_storage_data_840 <= (fillup_transition == 1'b1) ? i_input_data[60 % IN_WIDTH] : ping_storage_data_840 ^ i_input_data[60 % IN_WIDTH];
                469 / IN_WIDTH: ping_storage_data_840 <= (fillup_transition == 1'b1) ? i_input_data[469 % IN_WIDTH] : ping_storage_data_840 ^ i_input_data[469 % IN_WIDTH];
                528 / IN_WIDTH: ping_storage_data_840 <= (fillup_transition == 1'b1) ? i_input_data[528 % IN_WIDTH] : ping_storage_data_840 ^ i_input_data[528 % IN_WIDTH];
                701 / IN_WIDTH: ping_storage_data_840 <= (fillup_transition == 1'b1) ? i_input_data[701 % IN_WIDTH] : ping_storage_data_840 ^ i_input_data[701 % IN_WIDTH];
                1077 / IN_WIDTH: ping_storage_data_840 <= (fillup_transition == 1'b1) ? i_input_data[1077 % IN_WIDTH] : ping_storage_data_840 ^ i_input_data[1077 % IN_WIDTH];
                default: ping_storage_data_840 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_840;
                endcase
            end else begin
                case (input_count)
                60 / IN_WIDTH: pong_storage_data_840 <= (fillup_transition == 1'b1) ? i_input_data[60 % IN_WIDTH] : pong_storage_data_840 ^ i_input_data[60 % IN_WIDTH];
                469 / IN_WIDTH: pong_storage_data_840 <= (fillup_transition == 1'b1) ? i_input_data[469 % IN_WIDTH] : pong_storage_data_840 ^ i_input_data[469 % IN_WIDTH];
                528 / IN_WIDTH: pong_storage_data_840 <= (fillup_transition == 1'b1) ? i_input_data[528 % IN_WIDTH] : pong_storage_data_840 ^ i_input_data[528 % IN_WIDTH];
                701 / IN_WIDTH: pong_storage_data_840 <= (fillup_transition == 1'b1) ? i_input_data[701 % IN_WIDTH] : pong_storage_data_840 ^ i_input_data[701 % IN_WIDTH];
                1077 / IN_WIDTH: pong_storage_data_840 <= (fillup_transition == 1'b1) ? i_input_data[1077 % IN_WIDTH] : pong_storage_data_840 ^ i_input_data[1077 % IN_WIDTH];
                default: pong_storage_data_840 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_840;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_840 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_840;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_840 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_840;
            end
        end
    end
end

logic ping_storage_data_841;
logic pong_storage_data_841;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_841 <= 1'b0;
        pong_storage_data_841 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                61 / IN_WIDTH: ping_storage_data_841 <= (fillup_transition == 1'b1) ? i_input_data[61 % IN_WIDTH] : ping_storage_data_841 ^ i_input_data[61 % IN_WIDTH];
                470 / IN_WIDTH: ping_storage_data_841 <= (fillup_transition == 1'b1) ? i_input_data[470 % IN_WIDTH] : ping_storage_data_841 ^ i_input_data[470 % IN_WIDTH];
                529 / IN_WIDTH: ping_storage_data_841 <= (fillup_transition == 1'b1) ? i_input_data[529 % IN_WIDTH] : ping_storage_data_841 ^ i_input_data[529 % IN_WIDTH];
                702 / IN_WIDTH: ping_storage_data_841 <= (fillup_transition == 1'b1) ? i_input_data[702 % IN_WIDTH] : ping_storage_data_841 ^ i_input_data[702 % IN_WIDTH];
                1078 / IN_WIDTH: ping_storage_data_841 <= (fillup_transition == 1'b1) ? i_input_data[1078 % IN_WIDTH] : ping_storage_data_841 ^ i_input_data[1078 % IN_WIDTH];
                default: ping_storage_data_841 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_841;
                endcase
            end else begin
                case (input_count)
                61 / IN_WIDTH: pong_storage_data_841 <= (fillup_transition == 1'b1) ? i_input_data[61 % IN_WIDTH] : pong_storage_data_841 ^ i_input_data[61 % IN_WIDTH];
                470 / IN_WIDTH: pong_storage_data_841 <= (fillup_transition == 1'b1) ? i_input_data[470 % IN_WIDTH] : pong_storage_data_841 ^ i_input_data[470 % IN_WIDTH];
                529 / IN_WIDTH: pong_storage_data_841 <= (fillup_transition == 1'b1) ? i_input_data[529 % IN_WIDTH] : pong_storage_data_841 ^ i_input_data[529 % IN_WIDTH];
                702 / IN_WIDTH: pong_storage_data_841 <= (fillup_transition == 1'b1) ? i_input_data[702 % IN_WIDTH] : pong_storage_data_841 ^ i_input_data[702 % IN_WIDTH];
                1078 / IN_WIDTH: pong_storage_data_841 <= (fillup_transition == 1'b1) ? i_input_data[1078 % IN_WIDTH] : pong_storage_data_841 ^ i_input_data[1078 % IN_WIDTH];
                default: pong_storage_data_841 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_841;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_841 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_841;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_841 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_841;
            end
        end
    end
end

logic ping_storage_data_842;
logic pong_storage_data_842;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_842 <= 1'b0;
        pong_storage_data_842 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                62 / IN_WIDTH: ping_storage_data_842 <= (fillup_transition == 1'b1) ? i_input_data[62 % IN_WIDTH] : ping_storage_data_842 ^ i_input_data[62 % IN_WIDTH];
                471 / IN_WIDTH: ping_storage_data_842 <= (fillup_transition == 1'b1) ? i_input_data[471 % IN_WIDTH] : ping_storage_data_842 ^ i_input_data[471 % IN_WIDTH];
                530 / IN_WIDTH: ping_storage_data_842 <= (fillup_transition == 1'b1) ? i_input_data[530 % IN_WIDTH] : ping_storage_data_842 ^ i_input_data[530 % IN_WIDTH];
                703 / IN_WIDTH: ping_storage_data_842 <= (fillup_transition == 1'b1) ? i_input_data[703 % IN_WIDTH] : ping_storage_data_842 ^ i_input_data[703 % IN_WIDTH];
                1079 / IN_WIDTH: ping_storage_data_842 <= (fillup_transition == 1'b1) ? i_input_data[1079 % IN_WIDTH] : ping_storage_data_842 ^ i_input_data[1079 % IN_WIDTH];
                default: ping_storage_data_842 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_842;
                endcase
            end else begin
                case (input_count)
                62 / IN_WIDTH: pong_storage_data_842 <= (fillup_transition == 1'b1) ? i_input_data[62 % IN_WIDTH] : pong_storage_data_842 ^ i_input_data[62 % IN_WIDTH];
                471 / IN_WIDTH: pong_storage_data_842 <= (fillup_transition == 1'b1) ? i_input_data[471 % IN_WIDTH] : pong_storage_data_842 ^ i_input_data[471 % IN_WIDTH];
                530 / IN_WIDTH: pong_storage_data_842 <= (fillup_transition == 1'b1) ? i_input_data[530 % IN_WIDTH] : pong_storage_data_842 ^ i_input_data[530 % IN_WIDTH];
                703 / IN_WIDTH: pong_storage_data_842 <= (fillup_transition == 1'b1) ? i_input_data[703 % IN_WIDTH] : pong_storage_data_842 ^ i_input_data[703 % IN_WIDTH];
                1079 / IN_WIDTH: pong_storage_data_842 <= (fillup_transition == 1'b1) ? i_input_data[1079 % IN_WIDTH] : pong_storage_data_842 ^ i_input_data[1079 % IN_WIDTH];
                default: pong_storage_data_842 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_842;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_842 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_842;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_842 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_842;
            end
        end
    end
end

logic ping_storage_data_843;
logic pong_storage_data_843;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_843 <= 1'b0;
        pong_storage_data_843 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                63 / IN_WIDTH: ping_storage_data_843 <= (fillup_transition == 1'b1) ? i_input_data[63 % IN_WIDTH] : ping_storage_data_843 ^ i_input_data[63 % IN_WIDTH];
                472 / IN_WIDTH: ping_storage_data_843 <= (fillup_transition == 1'b1) ? i_input_data[472 % IN_WIDTH] : ping_storage_data_843 ^ i_input_data[472 % IN_WIDTH];
                531 / IN_WIDTH: ping_storage_data_843 <= (fillup_transition == 1'b1) ? i_input_data[531 % IN_WIDTH] : ping_storage_data_843 ^ i_input_data[531 % IN_WIDTH];
                704 / IN_WIDTH: ping_storage_data_843 <= (fillup_transition == 1'b1) ? i_input_data[704 % IN_WIDTH] : ping_storage_data_843 ^ i_input_data[704 % IN_WIDTH];
                1080 / IN_WIDTH: ping_storage_data_843 <= (fillup_transition == 1'b1) ? i_input_data[1080 % IN_WIDTH] : ping_storage_data_843 ^ i_input_data[1080 % IN_WIDTH];
                default: ping_storage_data_843 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_843;
                endcase
            end else begin
                case (input_count)
                63 / IN_WIDTH: pong_storage_data_843 <= (fillup_transition == 1'b1) ? i_input_data[63 % IN_WIDTH] : pong_storage_data_843 ^ i_input_data[63 % IN_WIDTH];
                472 / IN_WIDTH: pong_storage_data_843 <= (fillup_transition == 1'b1) ? i_input_data[472 % IN_WIDTH] : pong_storage_data_843 ^ i_input_data[472 % IN_WIDTH];
                531 / IN_WIDTH: pong_storage_data_843 <= (fillup_transition == 1'b1) ? i_input_data[531 % IN_WIDTH] : pong_storage_data_843 ^ i_input_data[531 % IN_WIDTH];
                704 / IN_WIDTH: pong_storage_data_843 <= (fillup_transition == 1'b1) ? i_input_data[704 % IN_WIDTH] : pong_storage_data_843 ^ i_input_data[704 % IN_WIDTH];
                1080 / IN_WIDTH: pong_storage_data_843 <= (fillup_transition == 1'b1) ? i_input_data[1080 % IN_WIDTH] : pong_storage_data_843 ^ i_input_data[1080 % IN_WIDTH];
                default: pong_storage_data_843 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_843;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_843 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_843;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_843 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_843;
            end
        end
    end
end

logic ping_storage_data_844;
logic pong_storage_data_844;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_844 <= 1'b0;
        pong_storage_data_844 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                64 / IN_WIDTH: ping_storage_data_844 <= (fillup_transition == 1'b1) ? i_input_data[64 % IN_WIDTH] : ping_storage_data_844 ^ i_input_data[64 % IN_WIDTH];
                473 / IN_WIDTH: ping_storage_data_844 <= (fillup_transition == 1'b1) ? i_input_data[473 % IN_WIDTH] : ping_storage_data_844 ^ i_input_data[473 % IN_WIDTH];
                532 / IN_WIDTH: ping_storage_data_844 <= (fillup_transition == 1'b1) ? i_input_data[532 % IN_WIDTH] : ping_storage_data_844 ^ i_input_data[532 % IN_WIDTH];
                705 / IN_WIDTH: ping_storage_data_844 <= (fillup_transition == 1'b1) ? i_input_data[705 % IN_WIDTH] : ping_storage_data_844 ^ i_input_data[705 % IN_WIDTH];
                1081 / IN_WIDTH: ping_storage_data_844 <= (fillup_transition == 1'b1) ? i_input_data[1081 % IN_WIDTH] : ping_storage_data_844 ^ i_input_data[1081 % IN_WIDTH];
                default: ping_storage_data_844 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_844;
                endcase
            end else begin
                case (input_count)
                64 / IN_WIDTH: pong_storage_data_844 <= (fillup_transition == 1'b1) ? i_input_data[64 % IN_WIDTH] : pong_storage_data_844 ^ i_input_data[64 % IN_WIDTH];
                473 / IN_WIDTH: pong_storage_data_844 <= (fillup_transition == 1'b1) ? i_input_data[473 % IN_WIDTH] : pong_storage_data_844 ^ i_input_data[473 % IN_WIDTH];
                532 / IN_WIDTH: pong_storage_data_844 <= (fillup_transition == 1'b1) ? i_input_data[532 % IN_WIDTH] : pong_storage_data_844 ^ i_input_data[532 % IN_WIDTH];
                705 / IN_WIDTH: pong_storage_data_844 <= (fillup_transition == 1'b1) ? i_input_data[705 % IN_WIDTH] : pong_storage_data_844 ^ i_input_data[705 % IN_WIDTH];
                1081 / IN_WIDTH: pong_storage_data_844 <= (fillup_transition == 1'b1) ? i_input_data[1081 % IN_WIDTH] : pong_storage_data_844 ^ i_input_data[1081 % IN_WIDTH];
                default: pong_storage_data_844 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_844;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_844 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_844;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_844 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_844;
            end
        end
    end
end

logic ping_storage_data_845;
logic pong_storage_data_845;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_845 <= 1'b0;
        pong_storage_data_845 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                65 / IN_WIDTH: ping_storage_data_845 <= (fillup_transition == 1'b1) ? i_input_data[65 % IN_WIDTH] : ping_storage_data_845 ^ i_input_data[65 % IN_WIDTH];
                474 / IN_WIDTH: ping_storage_data_845 <= (fillup_transition == 1'b1) ? i_input_data[474 % IN_WIDTH] : ping_storage_data_845 ^ i_input_data[474 % IN_WIDTH];
                533 / IN_WIDTH: ping_storage_data_845 <= (fillup_transition == 1'b1) ? i_input_data[533 % IN_WIDTH] : ping_storage_data_845 ^ i_input_data[533 % IN_WIDTH];
                706 / IN_WIDTH: ping_storage_data_845 <= (fillup_transition == 1'b1) ? i_input_data[706 % IN_WIDTH] : ping_storage_data_845 ^ i_input_data[706 % IN_WIDTH];
                1082 / IN_WIDTH: ping_storage_data_845 <= (fillup_transition == 1'b1) ? i_input_data[1082 % IN_WIDTH] : ping_storage_data_845 ^ i_input_data[1082 % IN_WIDTH];
                default: ping_storage_data_845 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_845;
                endcase
            end else begin
                case (input_count)
                65 / IN_WIDTH: pong_storage_data_845 <= (fillup_transition == 1'b1) ? i_input_data[65 % IN_WIDTH] : pong_storage_data_845 ^ i_input_data[65 % IN_WIDTH];
                474 / IN_WIDTH: pong_storage_data_845 <= (fillup_transition == 1'b1) ? i_input_data[474 % IN_WIDTH] : pong_storage_data_845 ^ i_input_data[474 % IN_WIDTH];
                533 / IN_WIDTH: pong_storage_data_845 <= (fillup_transition == 1'b1) ? i_input_data[533 % IN_WIDTH] : pong_storage_data_845 ^ i_input_data[533 % IN_WIDTH];
                706 / IN_WIDTH: pong_storage_data_845 <= (fillup_transition == 1'b1) ? i_input_data[706 % IN_WIDTH] : pong_storage_data_845 ^ i_input_data[706 % IN_WIDTH];
                1082 / IN_WIDTH: pong_storage_data_845 <= (fillup_transition == 1'b1) ? i_input_data[1082 % IN_WIDTH] : pong_storage_data_845 ^ i_input_data[1082 % IN_WIDTH];
                default: pong_storage_data_845 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_845;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_845 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_845;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_845 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_845;
            end
        end
    end
end

logic ping_storage_data_846;
logic pong_storage_data_846;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_846 <= 1'b0;
        pong_storage_data_846 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                66 / IN_WIDTH: ping_storage_data_846 <= (fillup_transition == 1'b1) ? i_input_data[66 % IN_WIDTH] : ping_storage_data_846 ^ i_input_data[66 % IN_WIDTH];
                475 / IN_WIDTH: ping_storage_data_846 <= (fillup_transition == 1'b1) ? i_input_data[475 % IN_WIDTH] : ping_storage_data_846 ^ i_input_data[475 % IN_WIDTH];
                534 / IN_WIDTH: ping_storage_data_846 <= (fillup_transition == 1'b1) ? i_input_data[534 % IN_WIDTH] : ping_storage_data_846 ^ i_input_data[534 % IN_WIDTH];
                707 / IN_WIDTH: ping_storage_data_846 <= (fillup_transition == 1'b1) ? i_input_data[707 % IN_WIDTH] : ping_storage_data_846 ^ i_input_data[707 % IN_WIDTH];
                1083 / IN_WIDTH: ping_storage_data_846 <= (fillup_transition == 1'b1) ? i_input_data[1083 % IN_WIDTH] : ping_storage_data_846 ^ i_input_data[1083 % IN_WIDTH];
                default: ping_storage_data_846 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_846;
                endcase
            end else begin
                case (input_count)
                66 / IN_WIDTH: pong_storage_data_846 <= (fillup_transition == 1'b1) ? i_input_data[66 % IN_WIDTH] : pong_storage_data_846 ^ i_input_data[66 % IN_WIDTH];
                475 / IN_WIDTH: pong_storage_data_846 <= (fillup_transition == 1'b1) ? i_input_data[475 % IN_WIDTH] : pong_storage_data_846 ^ i_input_data[475 % IN_WIDTH];
                534 / IN_WIDTH: pong_storage_data_846 <= (fillup_transition == 1'b1) ? i_input_data[534 % IN_WIDTH] : pong_storage_data_846 ^ i_input_data[534 % IN_WIDTH];
                707 / IN_WIDTH: pong_storage_data_846 <= (fillup_transition == 1'b1) ? i_input_data[707 % IN_WIDTH] : pong_storage_data_846 ^ i_input_data[707 % IN_WIDTH];
                1083 / IN_WIDTH: pong_storage_data_846 <= (fillup_transition == 1'b1) ? i_input_data[1083 % IN_WIDTH] : pong_storage_data_846 ^ i_input_data[1083 % IN_WIDTH];
                default: pong_storage_data_846 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_846;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_846 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_846;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_846 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_846;
            end
        end
    end
end

logic ping_storage_data_847;
logic pong_storage_data_847;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_847 <= 1'b0;
        pong_storage_data_847 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                67 / IN_WIDTH: ping_storage_data_847 <= (fillup_transition == 1'b1) ? i_input_data[67 % IN_WIDTH] : ping_storage_data_847 ^ i_input_data[67 % IN_WIDTH];
                476 / IN_WIDTH: ping_storage_data_847 <= (fillup_transition == 1'b1) ? i_input_data[476 % IN_WIDTH] : ping_storage_data_847 ^ i_input_data[476 % IN_WIDTH];
                535 / IN_WIDTH: ping_storage_data_847 <= (fillup_transition == 1'b1) ? i_input_data[535 % IN_WIDTH] : ping_storage_data_847 ^ i_input_data[535 % IN_WIDTH];
                708 / IN_WIDTH: ping_storage_data_847 <= (fillup_transition == 1'b1) ? i_input_data[708 % IN_WIDTH] : ping_storage_data_847 ^ i_input_data[708 % IN_WIDTH];
                1084 / IN_WIDTH: ping_storage_data_847 <= (fillup_transition == 1'b1) ? i_input_data[1084 % IN_WIDTH] : ping_storage_data_847 ^ i_input_data[1084 % IN_WIDTH];
                default: ping_storage_data_847 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_847;
                endcase
            end else begin
                case (input_count)
                67 / IN_WIDTH: pong_storage_data_847 <= (fillup_transition == 1'b1) ? i_input_data[67 % IN_WIDTH] : pong_storage_data_847 ^ i_input_data[67 % IN_WIDTH];
                476 / IN_WIDTH: pong_storage_data_847 <= (fillup_transition == 1'b1) ? i_input_data[476 % IN_WIDTH] : pong_storage_data_847 ^ i_input_data[476 % IN_WIDTH];
                535 / IN_WIDTH: pong_storage_data_847 <= (fillup_transition == 1'b1) ? i_input_data[535 % IN_WIDTH] : pong_storage_data_847 ^ i_input_data[535 % IN_WIDTH];
                708 / IN_WIDTH: pong_storage_data_847 <= (fillup_transition == 1'b1) ? i_input_data[708 % IN_WIDTH] : pong_storage_data_847 ^ i_input_data[708 % IN_WIDTH];
                1084 / IN_WIDTH: pong_storage_data_847 <= (fillup_transition == 1'b1) ? i_input_data[1084 % IN_WIDTH] : pong_storage_data_847 ^ i_input_data[1084 % IN_WIDTH];
                default: pong_storage_data_847 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_847;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_847 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_847;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_847 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_847;
            end
        end
    end
end

logic ping_storage_data_848;
logic pong_storage_data_848;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_848 <= 1'b0;
        pong_storage_data_848 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                68 / IN_WIDTH: ping_storage_data_848 <= (fillup_transition == 1'b1) ? i_input_data[68 % IN_WIDTH] : ping_storage_data_848 ^ i_input_data[68 % IN_WIDTH];
                477 / IN_WIDTH: ping_storage_data_848 <= (fillup_transition == 1'b1) ? i_input_data[477 % IN_WIDTH] : ping_storage_data_848 ^ i_input_data[477 % IN_WIDTH];
                536 / IN_WIDTH: ping_storage_data_848 <= (fillup_transition == 1'b1) ? i_input_data[536 % IN_WIDTH] : ping_storage_data_848 ^ i_input_data[536 % IN_WIDTH];
                709 / IN_WIDTH: ping_storage_data_848 <= (fillup_transition == 1'b1) ? i_input_data[709 % IN_WIDTH] : ping_storage_data_848 ^ i_input_data[709 % IN_WIDTH];
                1085 / IN_WIDTH: ping_storage_data_848 <= (fillup_transition == 1'b1) ? i_input_data[1085 % IN_WIDTH] : ping_storage_data_848 ^ i_input_data[1085 % IN_WIDTH];
                default: ping_storage_data_848 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_848;
                endcase
            end else begin
                case (input_count)
                68 / IN_WIDTH: pong_storage_data_848 <= (fillup_transition == 1'b1) ? i_input_data[68 % IN_WIDTH] : pong_storage_data_848 ^ i_input_data[68 % IN_WIDTH];
                477 / IN_WIDTH: pong_storage_data_848 <= (fillup_transition == 1'b1) ? i_input_data[477 % IN_WIDTH] : pong_storage_data_848 ^ i_input_data[477 % IN_WIDTH];
                536 / IN_WIDTH: pong_storage_data_848 <= (fillup_transition == 1'b1) ? i_input_data[536 % IN_WIDTH] : pong_storage_data_848 ^ i_input_data[536 % IN_WIDTH];
                709 / IN_WIDTH: pong_storage_data_848 <= (fillup_transition == 1'b1) ? i_input_data[709 % IN_WIDTH] : pong_storage_data_848 ^ i_input_data[709 % IN_WIDTH];
                1085 / IN_WIDTH: pong_storage_data_848 <= (fillup_transition == 1'b1) ? i_input_data[1085 % IN_WIDTH] : pong_storage_data_848 ^ i_input_data[1085 % IN_WIDTH];
                default: pong_storage_data_848 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_848;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_848 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_848;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_848 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_848;
            end
        end
    end
end

logic ping_storage_data_849;
logic pong_storage_data_849;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_849 <= 1'b0;
        pong_storage_data_849 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                69 / IN_WIDTH: ping_storage_data_849 <= (fillup_transition == 1'b1) ? i_input_data[69 % IN_WIDTH] : ping_storage_data_849 ^ i_input_data[69 % IN_WIDTH];
                478 / IN_WIDTH: ping_storage_data_849 <= (fillup_transition == 1'b1) ? i_input_data[478 % IN_WIDTH] : ping_storage_data_849 ^ i_input_data[478 % IN_WIDTH];
                537 / IN_WIDTH: ping_storage_data_849 <= (fillup_transition == 1'b1) ? i_input_data[537 % IN_WIDTH] : ping_storage_data_849 ^ i_input_data[537 % IN_WIDTH];
                710 / IN_WIDTH: ping_storage_data_849 <= (fillup_transition == 1'b1) ? i_input_data[710 % IN_WIDTH] : ping_storage_data_849 ^ i_input_data[710 % IN_WIDTH];
                1086 / IN_WIDTH: ping_storage_data_849 <= (fillup_transition == 1'b1) ? i_input_data[1086 % IN_WIDTH] : ping_storage_data_849 ^ i_input_data[1086 % IN_WIDTH];
                default: ping_storage_data_849 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_849;
                endcase
            end else begin
                case (input_count)
                69 / IN_WIDTH: pong_storage_data_849 <= (fillup_transition == 1'b1) ? i_input_data[69 % IN_WIDTH] : pong_storage_data_849 ^ i_input_data[69 % IN_WIDTH];
                478 / IN_WIDTH: pong_storage_data_849 <= (fillup_transition == 1'b1) ? i_input_data[478 % IN_WIDTH] : pong_storage_data_849 ^ i_input_data[478 % IN_WIDTH];
                537 / IN_WIDTH: pong_storage_data_849 <= (fillup_transition == 1'b1) ? i_input_data[537 % IN_WIDTH] : pong_storage_data_849 ^ i_input_data[537 % IN_WIDTH];
                710 / IN_WIDTH: pong_storage_data_849 <= (fillup_transition == 1'b1) ? i_input_data[710 % IN_WIDTH] : pong_storage_data_849 ^ i_input_data[710 % IN_WIDTH];
                1086 / IN_WIDTH: pong_storage_data_849 <= (fillup_transition == 1'b1) ? i_input_data[1086 % IN_WIDTH] : pong_storage_data_849 ^ i_input_data[1086 % IN_WIDTH];
                default: pong_storage_data_849 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_849;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_849 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_849;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_849 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_849;
            end
        end
    end
end

logic ping_storage_data_850;
logic pong_storage_data_850;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_850 <= 1'b0;
        pong_storage_data_850 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                70 / IN_WIDTH: ping_storage_data_850 <= (fillup_transition == 1'b1) ? i_input_data[70 % IN_WIDTH] : ping_storage_data_850 ^ i_input_data[70 % IN_WIDTH];
                479 / IN_WIDTH: ping_storage_data_850 <= (fillup_transition == 1'b1) ? i_input_data[479 % IN_WIDTH] : ping_storage_data_850 ^ i_input_data[479 % IN_WIDTH];
                538 / IN_WIDTH: ping_storage_data_850 <= (fillup_transition == 1'b1) ? i_input_data[538 % IN_WIDTH] : ping_storage_data_850 ^ i_input_data[538 % IN_WIDTH];
                711 / IN_WIDTH: ping_storage_data_850 <= (fillup_transition == 1'b1) ? i_input_data[711 % IN_WIDTH] : ping_storage_data_850 ^ i_input_data[711 % IN_WIDTH];
                1087 / IN_WIDTH: ping_storage_data_850 <= (fillup_transition == 1'b1) ? i_input_data[1087 % IN_WIDTH] : ping_storage_data_850 ^ i_input_data[1087 % IN_WIDTH];
                default: ping_storage_data_850 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_850;
                endcase
            end else begin
                case (input_count)
                70 / IN_WIDTH: pong_storage_data_850 <= (fillup_transition == 1'b1) ? i_input_data[70 % IN_WIDTH] : pong_storage_data_850 ^ i_input_data[70 % IN_WIDTH];
                479 / IN_WIDTH: pong_storage_data_850 <= (fillup_transition == 1'b1) ? i_input_data[479 % IN_WIDTH] : pong_storage_data_850 ^ i_input_data[479 % IN_WIDTH];
                538 / IN_WIDTH: pong_storage_data_850 <= (fillup_transition == 1'b1) ? i_input_data[538 % IN_WIDTH] : pong_storage_data_850 ^ i_input_data[538 % IN_WIDTH];
                711 / IN_WIDTH: pong_storage_data_850 <= (fillup_transition == 1'b1) ? i_input_data[711 % IN_WIDTH] : pong_storage_data_850 ^ i_input_data[711 % IN_WIDTH];
                1087 / IN_WIDTH: pong_storage_data_850 <= (fillup_transition == 1'b1) ? i_input_data[1087 % IN_WIDTH] : pong_storage_data_850 ^ i_input_data[1087 % IN_WIDTH];
                default: pong_storage_data_850 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_850;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_850 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_850;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_850 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_850;
            end
        end
    end
end

logic ping_storage_data_851;
logic pong_storage_data_851;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_851 <= 1'b0;
        pong_storage_data_851 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                71 / IN_WIDTH: ping_storage_data_851 <= (fillup_transition == 1'b1) ? i_input_data[71 % IN_WIDTH] : ping_storage_data_851 ^ i_input_data[71 % IN_WIDTH];
                384 / IN_WIDTH: ping_storage_data_851 <= (fillup_transition == 1'b1) ? i_input_data[384 % IN_WIDTH] : ping_storage_data_851 ^ i_input_data[384 % IN_WIDTH];
                539 / IN_WIDTH: ping_storage_data_851 <= (fillup_transition == 1'b1) ? i_input_data[539 % IN_WIDTH] : ping_storage_data_851 ^ i_input_data[539 % IN_WIDTH];
                712 / IN_WIDTH: ping_storage_data_851 <= (fillup_transition == 1'b1) ? i_input_data[712 % IN_WIDTH] : ping_storage_data_851 ^ i_input_data[712 % IN_WIDTH];
                1088 / IN_WIDTH: ping_storage_data_851 <= (fillup_transition == 1'b1) ? i_input_data[1088 % IN_WIDTH] : ping_storage_data_851 ^ i_input_data[1088 % IN_WIDTH];
                default: ping_storage_data_851 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_851;
                endcase
            end else begin
                case (input_count)
                71 / IN_WIDTH: pong_storage_data_851 <= (fillup_transition == 1'b1) ? i_input_data[71 % IN_WIDTH] : pong_storage_data_851 ^ i_input_data[71 % IN_WIDTH];
                384 / IN_WIDTH: pong_storage_data_851 <= (fillup_transition == 1'b1) ? i_input_data[384 % IN_WIDTH] : pong_storage_data_851 ^ i_input_data[384 % IN_WIDTH];
                539 / IN_WIDTH: pong_storage_data_851 <= (fillup_transition == 1'b1) ? i_input_data[539 % IN_WIDTH] : pong_storage_data_851 ^ i_input_data[539 % IN_WIDTH];
                712 / IN_WIDTH: pong_storage_data_851 <= (fillup_transition == 1'b1) ? i_input_data[712 % IN_WIDTH] : pong_storage_data_851 ^ i_input_data[712 % IN_WIDTH];
                1088 / IN_WIDTH: pong_storage_data_851 <= (fillup_transition == 1'b1) ? i_input_data[1088 % IN_WIDTH] : pong_storage_data_851 ^ i_input_data[1088 % IN_WIDTH];
                default: pong_storage_data_851 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_851;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_851 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_851;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_851 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_851;
            end
        end
    end
end

logic ping_storage_data_852;
logic pong_storage_data_852;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_852 <= 1'b0;
        pong_storage_data_852 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                72 / IN_WIDTH: ping_storage_data_852 <= (fillup_transition == 1'b1) ? i_input_data[72 % IN_WIDTH] : ping_storage_data_852 ^ i_input_data[72 % IN_WIDTH];
                385 / IN_WIDTH: ping_storage_data_852 <= (fillup_transition == 1'b1) ? i_input_data[385 % IN_WIDTH] : ping_storage_data_852 ^ i_input_data[385 % IN_WIDTH];
                540 / IN_WIDTH: ping_storage_data_852 <= (fillup_transition == 1'b1) ? i_input_data[540 % IN_WIDTH] : ping_storage_data_852 ^ i_input_data[540 % IN_WIDTH];
                713 / IN_WIDTH: ping_storage_data_852 <= (fillup_transition == 1'b1) ? i_input_data[713 % IN_WIDTH] : ping_storage_data_852 ^ i_input_data[713 % IN_WIDTH];
                1089 / IN_WIDTH: ping_storage_data_852 <= (fillup_transition == 1'b1) ? i_input_data[1089 % IN_WIDTH] : ping_storage_data_852 ^ i_input_data[1089 % IN_WIDTH];
                default: ping_storage_data_852 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_852;
                endcase
            end else begin
                case (input_count)
                72 / IN_WIDTH: pong_storage_data_852 <= (fillup_transition == 1'b1) ? i_input_data[72 % IN_WIDTH] : pong_storage_data_852 ^ i_input_data[72 % IN_WIDTH];
                385 / IN_WIDTH: pong_storage_data_852 <= (fillup_transition == 1'b1) ? i_input_data[385 % IN_WIDTH] : pong_storage_data_852 ^ i_input_data[385 % IN_WIDTH];
                540 / IN_WIDTH: pong_storage_data_852 <= (fillup_transition == 1'b1) ? i_input_data[540 % IN_WIDTH] : pong_storage_data_852 ^ i_input_data[540 % IN_WIDTH];
                713 / IN_WIDTH: pong_storage_data_852 <= (fillup_transition == 1'b1) ? i_input_data[713 % IN_WIDTH] : pong_storage_data_852 ^ i_input_data[713 % IN_WIDTH];
                1089 / IN_WIDTH: pong_storage_data_852 <= (fillup_transition == 1'b1) ? i_input_data[1089 % IN_WIDTH] : pong_storage_data_852 ^ i_input_data[1089 % IN_WIDTH];
                default: pong_storage_data_852 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_852;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_852 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_852;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_852 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_852;
            end
        end
    end
end

logic ping_storage_data_853;
logic pong_storage_data_853;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_853 <= 1'b0;
        pong_storage_data_853 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                73 / IN_WIDTH: ping_storage_data_853 <= (fillup_transition == 1'b1) ? i_input_data[73 % IN_WIDTH] : ping_storage_data_853 ^ i_input_data[73 % IN_WIDTH];
                386 / IN_WIDTH: ping_storage_data_853 <= (fillup_transition == 1'b1) ? i_input_data[386 % IN_WIDTH] : ping_storage_data_853 ^ i_input_data[386 % IN_WIDTH];
                541 / IN_WIDTH: ping_storage_data_853 <= (fillup_transition == 1'b1) ? i_input_data[541 % IN_WIDTH] : ping_storage_data_853 ^ i_input_data[541 % IN_WIDTH];
                714 / IN_WIDTH: ping_storage_data_853 <= (fillup_transition == 1'b1) ? i_input_data[714 % IN_WIDTH] : ping_storage_data_853 ^ i_input_data[714 % IN_WIDTH];
                1090 / IN_WIDTH: ping_storage_data_853 <= (fillup_transition == 1'b1) ? i_input_data[1090 % IN_WIDTH] : ping_storage_data_853 ^ i_input_data[1090 % IN_WIDTH];
                default: ping_storage_data_853 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_853;
                endcase
            end else begin
                case (input_count)
                73 / IN_WIDTH: pong_storage_data_853 <= (fillup_transition == 1'b1) ? i_input_data[73 % IN_WIDTH] : pong_storage_data_853 ^ i_input_data[73 % IN_WIDTH];
                386 / IN_WIDTH: pong_storage_data_853 <= (fillup_transition == 1'b1) ? i_input_data[386 % IN_WIDTH] : pong_storage_data_853 ^ i_input_data[386 % IN_WIDTH];
                541 / IN_WIDTH: pong_storage_data_853 <= (fillup_transition == 1'b1) ? i_input_data[541 % IN_WIDTH] : pong_storage_data_853 ^ i_input_data[541 % IN_WIDTH];
                714 / IN_WIDTH: pong_storage_data_853 <= (fillup_transition == 1'b1) ? i_input_data[714 % IN_WIDTH] : pong_storage_data_853 ^ i_input_data[714 % IN_WIDTH];
                1090 / IN_WIDTH: pong_storage_data_853 <= (fillup_transition == 1'b1) ? i_input_data[1090 % IN_WIDTH] : pong_storage_data_853 ^ i_input_data[1090 % IN_WIDTH];
                default: pong_storage_data_853 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_853;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_853 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_853;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_853 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_853;
            end
        end
    end
end

logic ping_storage_data_854;
logic pong_storage_data_854;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_854 <= 1'b0;
        pong_storage_data_854 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                74 / IN_WIDTH: ping_storage_data_854 <= (fillup_transition == 1'b1) ? i_input_data[74 % IN_WIDTH] : ping_storage_data_854 ^ i_input_data[74 % IN_WIDTH];
                387 / IN_WIDTH: ping_storage_data_854 <= (fillup_transition == 1'b1) ? i_input_data[387 % IN_WIDTH] : ping_storage_data_854 ^ i_input_data[387 % IN_WIDTH];
                542 / IN_WIDTH: ping_storage_data_854 <= (fillup_transition == 1'b1) ? i_input_data[542 % IN_WIDTH] : ping_storage_data_854 ^ i_input_data[542 % IN_WIDTH];
                715 / IN_WIDTH: ping_storage_data_854 <= (fillup_transition == 1'b1) ? i_input_data[715 % IN_WIDTH] : ping_storage_data_854 ^ i_input_data[715 % IN_WIDTH];
                1091 / IN_WIDTH: ping_storage_data_854 <= (fillup_transition == 1'b1) ? i_input_data[1091 % IN_WIDTH] : ping_storage_data_854 ^ i_input_data[1091 % IN_WIDTH];
                default: ping_storage_data_854 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_854;
                endcase
            end else begin
                case (input_count)
                74 / IN_WIDTH: pong_storage_data_854 <= (fillup_transition == 1'b1) ? i_input_data[74 % IN_WIDTH] : pong_storage_data_854 ^ i_input_data[74 % IN_WIDTH];
                387 / IN_WIDTH: pong_storage_data_854 <= (fillup_transition == 1'b1) ? i_input_data[387 % IN_WIDTH] : pong_storage_data_854 ^ i_input_data[387 % IN_WIDTH];
                542 / IN_WIDTH: pong_storage_data_854 <= (fillup_transition == 1'b1) ? i_input_data[542 % IN_WIDTH] : pong_storage_data_854 ^ i_input_data[542 % IN_WIDTH];
                715 / IN_WIDTH: pong_storage_data_854 <= (fillup_transition == 1'b1) ? i_input_data[715 % IN_WIDTH] : pong_storage_data_854 ^ i_input_data[715 % IN_WIDTH];
                1091 / IN_WIDTH: pong_storage_data_854 <= (fillup_transition == 1'b1) ? i_input_data[1091 % IN_WIDTH] : pong_storage_data_854 ^ i_input_data[1091 % IN_WIDTH];
                default: pong_storage_data_854 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_854;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_854 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_854;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_854 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_854;
            end
        end
    end
end

logic ping_storage_data_855;
logic pong_storage_data_855;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_855 <= 1'b0;
        pong_storage_data_855 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                75 / IN_WIDTH: ping_storage_data_855 <= (fillup_transition == 1'b1) ? i_input_data[75 % IN_WIDTH] : ping_storage_data_855 ^ i_input_data[75 % IN_WIDTH];
                388 / IN_WIDTH: ping_storage_data_855 <= (fillup_transition == 1'b1) ? i_input_data[388 % IN_WIDTH] : ping_storage_data_855 ^ i_input_data[388 % IN_WIDTH];
                543 / IN_WIDTH: ping_storage_data_855 <= (fillup_transition == 1'b1) ? i_input_data[543 % IN_WIDTH] : ping_storage_data_855 ^ i_input_data[543 % IN_WIDTH];
                716 / IN_WIDTH: ping_storage_data_855 <= (fillup_transition == 1'b1) ? i_input_data[716 % IN_WIDTH] : ping_storage_data_855 ^ i_input_data[716 % IN_WIDTH];
                1092 / IN_WIDTH: ping_storage_data_855 <= (fillup_transition == 1'b1) ? i_input_data[1092 % IN_WIDTH] : ping_storage_data_855 ^ i_input_data[1092 % IN_WIDTH];
                default: ping_storage_data_855 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_855;
                endcase
            end else begin
                case (input_count)
                75 / IN_WIDTH: pong_storage_data_855 <= (fillup_transition == 1'b1) ? i_input_data[75 % IN_WIDTH] : pong_storage_data_855 ^ i_input_data[75 % IN_WIDTH];
                388 / IN_WIDTH: pong_storage_data_855 <= (fillup_transition == 1'b1) ? i_input_data[388 % IN_WIDTH] : pong_storage_data_855 ^ i_input_data[388 % IN_WIDTH];
                543 / IN_WIDTH: pong_storage_data_855 <= (fillup_transition == 1'b1) ? i_input_data[543 % IN_WIDTH] : pong_storage_data_855 ^ i_input_data[543 % IN_WIDTH];
                716 / IN_WIDTH: pong_storage_data_855 <= (fillup_transition == 1'b1) ? i_input_data[716 % IN_WIDTH] : pong_storage_data_855 ^ i_input_data[716 % IN_WIDTH];
                1092 / IN_WIDTH: pong_storage_data_855 <= (fillup_transition == 1'b1) ? i_input_data[1092 % IN_WIDTH] : pong_storage_data_855 ^ i_input_data[1092 % IN_WIDTH];
                default: pong_storage_data_855 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_855;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_855 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_855;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_855 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_855;
            end
        end
    end
end

logic ping_storage_data_856;
logic pong_storage_data_856;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_856 <= 1'b0;
        pong_storage_data_856 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                76 / IN_WIDTH: ping_storage_data_856 <= (fillup_transition == 1'b1) ? i_input_data[76 % IN_WIDTH] : ping_storage_data_856 ^ i_input_data[76 % IN_WIDTH];
                389 / IN_WIDTH: ping_storage_data_856 <= (fillup_transition == 1'b1) ? i_input_data[389 % IN_WIDTH] : ping_storage_data_856 ^ i_input_data[389 % IN_WIDTH];
                544 / IN_WIDTH: ping_storage_data_856 <= (fillup_transition == 1'b1) ? i_input_data[544 % IN_WIDTH] : ping_storage_data_856 ^ i_input_data[544 % IN_WIDTH];
                717 / IN_WIDTH: ping_storage_data_856 <= (fillup_transition == 1'b1) ? i_input_data[717 % IN_WIDTH] : ping_storage_data_856 ^ i_input_data[717 % IN_WIDTH];
                1093 / IN_WIDTH: ping_storage_data_856 <= (fillup_transition == 1'b1) ? i_input_data[1093 % IN_WIDTH] : ping_storage_data_856 ^ i_input_data[1093 % IN_WIDTH];
                default: ping_storage_data_856 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_856;
                endcase
            end else begin
                case (input_count)
                76 / IN_WIDTH: pong_storage_data_856 <= (fillup_transition == 1'b1) ? i_input_data[76 % IN_WIDTH] : pong_storage_data_856 ^ i_input_data[76 % IN_WIDTH];
                389 / IN_WIDTH: pong_storage_data_856 <= (fillup_transition == 1'b1) ? i_input_data[389 % IN_WIDTH] : pong_storage_data_856 ^ i_input_data[389 % IN_WIDTH];
                544 / IN_WIDTH: pong_storage_data_856 <= (fillup_transition == 1'b1) ? i_input_data[544 % IN_WIDTH] : pong_storage_data_856 ^ i_input_data[544 % IN_WIDTH];
                717 / IN_WIDTH: pong_storage_data_856 <= (fillup_transition == 1'b1) ? i_input_data[717 % IN_WIDTH] : pong_storage_data_856 ^ i_input_data[717 % IN_WIDTH];
                1093 / IN_WIDTH: pong_storage_data_856 <= (fillup_transition == 1'b1) ? i_input_data[1093 % IN_WIDTH] : pong_storage_data_856 ^ i_input_data[1093 % IN_WIDTH];
                default: pong_storage_data_856 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_856;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_856 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_856;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_856 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_856;
            end
        end
    end
end

logic ping_storage_data_857;
logic pong_storage_data_857;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_857 <= 1'b0;
        pong_storage_data_857 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                77 / IN_WIDTH: ping_storage_data_857 <= (fillup_transition == 1'b1) ? i_input_data[77 % IN_WIDTH] : ping_storage_data_857 ^ i_input_data[77 % IN_WIDTH];
                390 / IN_WIDTH: ping_storage_data_857 <= (fillup_transition == 1'b1) ? i_input_data[390 % IN_WIDTH] : ping_storage_data_857 ^ i_input_data[390 % IN_WIDTH];
                545 / IN_WIDTH: ping_storage_data_857 <= (fillup_transition == 1'b1) ? i_input_data[545 % IN_WIDTH] : ping_storage_data_857 ^ i_input_data[545 % IN_WIDTH];
                718 / IN_WIDTH: ping_storage_data_857 <= (fillup_transition == 1'b1) ? i_input_data[718 % IN_WIDTH] : ping_storage_data_857 ^ i_input_data[718 % IN_WIDTH];
                1094 / IN_WIDTH: ping_storage_data_857 <= (fillup_transition == 1'b1) ? i_input_data[1094 % IN_WIDTH] : ping_storage_data_857 ^ i_input_data[1094 % IN_WIDTH];
                default: ping_storage_data_857 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_857;
                endcase
            end else begin
                case (input_count)
                77 / IN_WIDTH: pong_storage_data_857 <= (fillup_transition == 1'b1) ? i_input_data[77 % IN_WIDTH] : pong_storage_data_857 ^ i_input_data[77 % IN_WIDTH];
                390 / IN_WIDTH: pong_storage_data_857 <= (fillup_transition == 1'b1) ? i_input_data[390 % IN_WIDTH] : pong_storage_data_857 ^ i_input_data[390 % IN_WIDTH];
                545 / IN_WIDTH: pong_storage_data_857 <= (fillup_transition == 1'b1) ? i_input_data[545 % IN_WIDTH] : pong_storage_data_857 ^ i_input_data[545 % IN_WIDTH];
                718 / IN_WIDTH: pong_storage_data_857 <= (fillup_transition == 1'b1) ? i_input_data[718 % IN_WIDTH] : pong_storage_data_857 ^ i_input_data[718 % IN_WIDTH];
                1094 / IN_WIDTH: pong_storage_data_857 <= (fillup_transition == 1'b1) ? i_input_data[1094 % IN_WIDTH] : pong_storage_data_857 ^ i_input_data[1094 % IN_WIDTH];
                default: pong_storage_data_857 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_857;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_857 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_857;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_857 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_857;
            end
        end
    end
end

logic ping_storage_data_858;
logic pong_storage_data_858;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_858 <= 1'b0;
        pong_storage_data_858 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                78 / IN_WIDTH: ping_storage_data_858 <= (fillup_transition == 1'b1) ? i_input_data[78 % IN_WIDTH] : ping_storage_data_858 ^ i_input_data[78 % IN_WIDTH];
                391 / IN_WIDTH: ping_storage_data_858 <= (fillup_transition == 1'b1) ? i_input_data[391 % IN_WIDTH] : ping_storage_data_858 ^ i_input_data[391 % IN_WIDTH];
                546 / IN_WIDTH: ping_storage_data_858 <= (fillup_transition == 1'b1) ? i_input_data[546 % IN_WIDTH] : ping_storage_data_858 ^ i_input_data[546 % IN_WIDTH];
                719 / IN_WIDTH: ping_storage_data_858 <= (fillup_transition == 1'b1) ? i_input_data[719 % IN_WIDTH] : ping_storage_data_858 ^ i_input_data[719 % IN_WIDTH];
                1095 / IN_WIDTH: ping_storage_data_858 <= (fillup_transition == 1'b1) ? i_input_data[1095 % IN_WIDTH] : ping_storage_data_858 ^ i_input_data[1095 % IN_WIDTH];
                default: ping_storage_data_858 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_858;
                endcase
            end else begin
                case (input_count)
                78 / IN_WIDTH: pong_storage_data_858 <= (fillup_transition == 1'b1) ? i_input_data[78 % IN_WIDTH] : pong_storage_data_858 ^ i_input_data[78 % IN_WIDTH];
                391 / IN_WIDTH: pong_storage_data_858 <= (fillup_transition == 1'b1) ? i_input_data[391 % IN_WIDTH] : pong_storage_data_858 ^ i_input_data[391 % IN_WIDTH];
                546 / IN_WIDTH: pong_storage_data_858 <= (fillup_transition == 1'b1) ? i_input_data[546 % IN_WIDTH] : pong_storage_data_858 ^ i_input_data[546 % IN_WIDTH];
                719 / IN_WIDTH: pong_storage_data_858 <= (fillup_transition == 1'b1) ? i_input_data[719 % IN_WIDTH] : pong_storage_data_858 ^ i_input_data[719 % IN_WIDTH];
                1095 / IN_WIDTH: pong_storage_data_858 <= (fillup_transition == 1'b1) ? i_input_data[1095 % IN_WIDTH] : pong_storage_data_858 ^ i_input_data[1095 % IN_WIDTH];
                default: pong_storage_data_858 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_858;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_858 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_858;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_858 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_858;
            end
        end
    end
end

logic ping_storage_data_859;
logic pong_storage_data_859;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_859 <= 1'b0;
        pong_storage_data_859 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                79 / IN_WIDTH: ping_storage_data_859 <= (fillup_transition == 1'b1) ? i_input_data[79 % IN_WIDTH] : ping_storage_data_859 ^ i_input_data[79 % IN_WIDTH];
                392 / IN_WIDTH: ping_storage_data_859 <= (fillup_transition == 1'b1) ? i_input_data[392 % IN_WIDTH] : ping_storage_data_859 ^ i_input_data[392 % IN_WIDTH];
                547 / IN_WIDTH: ping_storage_data_859 <= (fillup_transition == 1'b1) ? i_input_data[547 % IN_WIDTH] : ping_storage_data_859 ^ i_input_data[547 % IN_WIDTH];
                720 / IN_WIDTH: ping_storage_data_859 <= (fillup_transition == 1'b1) ? i_input_data[720 % IN_WIDTH] : ping_storage_data_859 ^ i_input_data[720 % IN_WIDTH];
                1096 / IN_WIDTH: ping_storage_data_859 <= (fillup_transition == 1'b1) ? i_input_data[1096 % IN_WIDTH] : ping_storage_data_859 ^ i_input_data[1096 % IN_WIDTH];
                default: ping_storage_data_859 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_859;
                endcase
            end else begin
                case (input_count)
                79 / IN_WIDTH: pong_storage_data_859 <= (fillup_transition == 1'b1) ? i_input_data[79 % IN_WIDTH] : pong_storage_data_859 ^ i_input_data[79 % IN_WIDTH];
                392 / IN_WIDTH: pong_storage_data_859 <= (fillup_transition == 1'b1) ? i_input_data[392 % IN_WIDTH] : pong_storage_data_859 ^ i_input_data[392 % IN_WIDTH];
                547 / IN_WIDTH: pong_storage_data_859 <= (fillup_transition == 1'b1) ? i_input_data[547 % IN_WIDTH] : pong_storage_data_859 ^ i_input_data[547 % IN_WIDTH];
                720 / IN_WIDTH: pong_storage_data_859 <= (fillup_transition == 1'b1) ? i_input_data[720 % IN_WIDTH] : pong_storage_data_859 ^ i_input_data[720 % IN_WIDTH];
                1096 / IN_WIDTH: pong_storage_data_859 <= (fillup_transition == 1'b1) ? i_input_data[1096 % IN_WIDTH] : pong_storage_data_859 ^ i_input_data[1096 % IN_WIDTH];
                default: pong_storage_data_859 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_859;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_859 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_859;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_859 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_859;
            end
        end
    end
end

logic ping_storage_data_860;
logic pong_storage_data_860;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_860 <= 1'b0;
        pong_storage_data_860 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                80 / IN_WIDTH: ping_storage_data_860 <= (fillup_transition == 1'b1) ? i_input_data[80 % IN_WIDTH] : ping_storage_data_860 ^ i_input_data[80 % IN_WIDTH];
                393 / IN_WIDTH: ping_storage_data_860 <= (fillup_transition == 1'b1) ? i_input_data[393 % IN_WIDTH] : ping_storage_data_860 ^ i_input_data[393 % IN_WIDTH];
                548 / IN_WIDTH: ping_storage_data_860 <= (fillup_transition == 1'b1) ? i_input_data[548 % IN_WIDTH] : ping_storage_data_860 ^ i_input_data[548 % IN_WIDTH];
                721 / IN_WIDTH: ping_storage_data_860 <= (fillup_transition == 1'b1) ? i_input_data[721 % IN_WIDTH] : ping_storage_data_860 ^ i_input_data[721 % IN_WIDTH];
                1097 / IN_WIDTH: ping_storage_data_860 <= (fillup_transition == 1'b1) ? i_input_data[1097 % IN_WIDTH] : ping_storage_data_860 ^ i_input_data[1097 % IN_WIDTH];
                default: ping_storage_data_860 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_860;
                endcase
            end else begin
                case (input_count)
                80 / IN_WIDTH: pong_storage_data_860 <= (fillup_transition == 1'b1) ? i_input_data[80 % IN_WIDTH] : pong_storage_data_860 ^ i_input_data[80 % IN_WIDTH];
                393 / IN_WIDTH: pong_storage_data_860 <= (fillup_transition == 1'b1) ? i_input_data[393 % IN_WIDTH] : pong_storage_data_860 ^ i_input_data[393 % IN_WIDTH];
                548 / IN_WIDTH: pong_storage_data_860 <= (fillup_transition == 1'b1) ? i_input_data[548 % IN_WIDTH] : pong_storage_data_860 ^ i_input_data[548 % IN_WIDTH];
                721 / IN_WIDTH: pong_storage_data_860 <= (fillup_transition == 1'b1) ? i_input_data[721 % IN_WIDTH] : pong_storage_data_860 ^ i_input_data[721 % IN_WIDTH];
                1097 / IN_WIDTH: pong_storage_data_860 <= (fillup_transition == 1'b1) ? i_input_data[1097 % IN_WIDTH] : pong_storage_data_860 ^ i_input_data[1097 % IN_WIDTH];
                default: pong_storage_data_860 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_860;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_860 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_860;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_860 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_860;
            end
        end
    end
end

logic ping_storage_data_861;
logic pong_storage_data_861;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_861 <= 1'b0;
        pong_storage_data_861 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                81 / IN_WIDTH: ping_storage_data_861 <= (fillup_transition == 1'b1) ? i_input_data[81 % IN_WIDTH] : ping_storage_data_861 ^ i_input_data[81 % IN_WIDTH];
                394 / IN_WIDTH: ping_storage_data_861 <= (fillup_transition == 1'b1) ? i_input_data[394 % IN_WIDTH] : ping_storage_data_861 ^ i_input_data[394 % IN_WIDTH];
                549 / IN_WIDTH: ping_storage_data_861 <= (fillup_transition == 1'b1) ? i_input_data[549 % IN_WIDTH] : ping_storage_data_861 ^ i_input_data[549 % IN_WIDTH];
                722 / IN_WIDTH: ping_storage_data_861 <= (fillup_transition == 1'b1) ? i_input_data[722 % IN_WIDTH] : ping_storage_data_861 ^ i_input_data[722 % IN_WIDTH];
                1098 / IN_WIDTH: ping_storage_data_861 <= (fillup_transition == 1'b1) ? i_input_data[1098 % IN_WIDTH] : ping_storage_data_861 ^ i_input_data[1098 % IN_WIDTH];
                default: ping_storage_data_861 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_861;
                endcase
            end else begin
                case (input_count)
                81 / IN_WIDTH: pong_storage_data_861 <= (fillup_transition == 1'b1) ? i_input_data[81 % IN_WIDTH] : pong_storage_data_861 ^ i_input_data[81 % IN_WIDTH];
                394 / IN_WIDTH: pong_storage_data_861 <= (fillup_transition == 1'b1) ? i_input_data[394 % IN_WIDTH] : pong_storage_data_861 ^ i_input_data[394 % IN_WIDTH];
                549 / IN_WIDTH: pong_storage_data_861 <= (fillup_transition == 1'b1) ? i_input_data[549 % IN_WIDTH] : pong_storage_data_861 ^ i_input_data[549 % IN_WIDTH];
                722 / IN_WIDTH: pong_storage_data_861 <= (fillup_transition == 1'b1) ? i_input_data[722 % IN_WIDTH] : pong_storage_data_861 ^ i_input_data[722 % IN_WIDTH];
                1098 / IN_WIDTH: pong_storage_data_861 <= (fillup_transition == 1'b1) ? i_input_data[1098 % IN_WIDTH] : pong_storage_data_861 ^ i_input_data[1098 % IN_WIDTH];
                default: pong_storage_data_861 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_861;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_861 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_861;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_861 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_861;
            end
        end
    end
end

logic ping_storage_data_862;
logic pong_storage_data_862;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_862 <= 1'b0;
        pong_storage_data_862 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                82 / IN_WIDTH: ping_storage_data_862 <= (fillup_transition == 1'b1) ? i_input_data[82 % IN_WIDTH] : ping_storage_data_862 ^ i_input_data[82 % IN_WIDTH];
                395 / IN_WIDTH: ping_storage_data_862 <= (fillup_transition == 1'b1) ? i_input_data[395 % IN_WIDTH] : ping_storage_data_862 ^ i_input_data[395 % IN_WIDTH];
                550 / IN_WIDTH: ping_storage_data_862 <= (fillup_transition == 1'b1) ? i_input_data[550 % IN_WIDTH] : ping_storage_data_862 ^ i_input_data[550 % IN_WIDTH];
                723 / IN_WIDTH: ping_storage_data_862 <= (fillup_transition == 1'b1) ? i_input_data[723 % IN_WIDTH] : ping_storage_data_862 ^ i_input_data[723 % IN_WIDTH];
                1099 / IN_WIDTH: ping_storage_data_862 <= (fillup_transition == 1'b1) ? i_input_data[1099 % IN_WIDTH] : ping_storage_data_862 ^ i_input_data[1099 % IN_WIDTH];
                default: ping_storage_data_862 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_862;
                endcase
            end else begin
                case (input_count)
                82 / IN_WIDTH: pong_storage_data_862 <= (fillup_transition == 1'b1) ? i_input_data[82 % IN_WIDTH] : pong_storage_data_862 ^ i_input_data[82 % IN_WIDTH];
                395 / IN_WIDTH: pong_storage_data_862 <= (fillup_transition == 1'b1) ? i_input_data[395 % IN_WIDTH] : pong_storage_data_862 ^ i_input_data[395 % IN_WIDTH];
                550 / IN_WIDTH: pong_storage_data_862 <= (fillup_transition == 1'b1) ? i_input_data[550 % IN_WIDTH] : pong_storage_data_862 ^ i_input_data[550 % IN_WIDTH];
                723 / IN_WIDTH: pong_storage_data_862 <= (fillup_transition == 1'b1) ? i_input_data[723 % IN_WIDTH] : pong_storage_data_862 ^ i_input_data[723 % IN_WIDTH];
                1099 / IN_WIDTH: pong_storage_data_862 <= (fillup_transition == 1'b1) ? i_input_data[1099 % IN_WIDTH] : pong_storage_data_862 ^ i_input_data[1099 % IN_WIDTH];
                default: pong_storage_data_862 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_862;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_862 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_862;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_862 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_862;
            end
        end
    end
end

logic ping_storage_data_863;
logic pong_storage_data_863;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_863 <= 1'b0;
        pong_storage_data_863 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                83 / IN_WIDTH: ping_storage_data_863 <= (fillup_transition == 1'b1) ? i_input_data[83 % IN_WIDTH] : ping_storage_data_863 ^ i_input_data[83 % IN_WIDTH];
                396 / IN_WIDTH: ping_storage_data_863 <= (fillup_transition == 1'b1) ? i_input_data[396 % IN_WIDTH] : ping_storage_data_863 ^ i_input_data[396 % IN_WIDTH];
                551 / IN_WIDTH: ping_storage_data_863 <= (fillup_transition == 1'b1) ? i_input_data[551 % IN_WIDTH] : ping_storage_data_863 ^ i_input_data[551 % IN_WIDTH];
                724 / IN_WIDTH: ping_storage_data_863 <= (fillup_transition == 1'b1) ? i_input_data[724 % IN_WIDTH] : ping_storage_data_863 ^ i_input_data[724 % IN_WIDTH];
                1100 / IN_WIDTH: ping_storage_data_863 <= (fillup_transition == 1'b1) ? i_input_data[1100 % IN_WIDTH] : ping_storage_data_863 ^ i_input_data[1100 % IN_WIDTH];
                default: ping_storage_data_863 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_863;
                endcase
            end else begin
                case (input_count)
                83 / IN_WIDTH: pong_storage_data_863 <= (fillup_transition == 1'b1) ? i_input_data[83 % IN_WIDTH] : pong_storage_data_863 ^ i_input_data[83 % IN_WIDTH];
                396 / IN_WIDTH: pong_storage_data_863 <= (fillup_transition == 1'b1) ? i_input_data[396 % IN_WIDTH] : pong_storage_data_863 ^ i_input_data[396 % IN_WIDTH];
                551 / IN_WIDTH: pong_storage_data_863 <= (fillup_transition == 1'b1) ? i_input_data[551 % IN_WIDTH] : pong_storage_data_863 ^ i_input_data[551 % IN_WIDTH];
                724 / IN_WIDTH: pong_storage_data_863 <= (fillup_transition == 1'b1) ? i_input_data[724 % IN_WIDTH] : pong_storage_data_863 ^ i_input_data[724 % IN_WIDTH];
                1100 / IN_WIDTH: pong_storage_data_863 <= (fillup_transition == 1'b1) ? i_input_data[1100 % IN_WIDTH] : pong_storage_data_863 ^ i_input_data[1100 % IN_WIDTH];
                default: pong_storage_data_863 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_863;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_863 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_863;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_863 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_863;
            end
        end
    end
end

logic ping_storage_data_864;
logic pong_storage_data_864;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_864 <= 1'b0;
        pong_storage_data_864 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                482 / IN_WIDTH: ping_storage_data_864 <= (fillup_transition == 1'b1) ? i_input_data[482 % IN_WIDTH] : ping_storage_data_864 ^ i_input_data[482 % IN_WIDTH];
                709 / IN_WIDTH: ping_storage_data_864 <= (fillup_transition == 1'b1) ? i_input_data[709 % IN_WIDTH] : ping_storage_data_864 ^ i_input_data[709 % IN_WIDTH];
                986 / IN_WIDTH: ping_storage_data_864 <= (fillup_transition == 1'b1) ? i_input_data[986 % IN_WIDTH] : ping_storage_data_864 ^ i_input_data[986 % IN_WIDTH];
                1080 / IN_WIDTH: ping_storage_data_864 <= (fillup_transition == 1'b1) ? i_input_data[1080 % IN_WIDTH] : ping_storage_data_864 ^ i_input_data[1080 % IN_WIDTH];
                default: ping_storage_data_864 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_864;
                endcase
            end else begin
                case (input_count)
                482 / IN_WIDTH: pong_storage_data_864 <= (fillup_transition == 1'b1) ? i_input_data[482 % IN_WIDTH] : pong_storage_data_864 ^ i_input_data[482 % IN_WIDTH];
                709 / IN_WIDTH: pong_storage_data_864 <= (fillup_transition == 1'b1) ? i_input_data[709 % IN_WIDTH] : pong_storage_data_864 ^ i_input_data[709 % IN_WIDTH];
                986 / IN_WIDTH: pong_storage_data_864 <= (fillup_transition == 1'b1) ? i_input_data[986 % IN_WIDTH] : pong_storage_data_864 ^ i_input_data[986 % IN_WIDTH];
                1080 / IN_WIDTH: pong_storage_data_864 <= (fillup_transition == 1'b1) ? i_input_data[1080 % IN_WIDTH] : pong_storage_data_864 ^ i_input_data[1080 % IN_WIDTH];
                default: pong_storage_data_864 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_864;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_864 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_864;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_864 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_864;
            end
        end
    end
end

logic ping_storage_data_865;
logic pong_storage_data_865;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_865 <= 1'b0;
        pong_storage_data_865 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                483 / IN_WIDTH: ping_storage_data_865 <= (fillup_transition == 1'b1) ? i_input_data[483 % IN_WIDTH] : ping_storage_data_865 ^ i_input_data[483 % IN_WIDTH];
                710 / IN_WIDTH: ping_storage_data_865 <= (fillup_transition == 1'b1) ? i_input_data[710 % IN_WIDTH] : ping_storage_data_865 ^ i_input_data[710 % IN_WIDTH];
                987 / IN_WIDTH: ping_storage_data_865 <= (fillup_transition == 1'b1) ? i_input_data[987 % IN_WIDTH] : ping_storage_data_865 ^ i_input_data[987 % IN_WIDTH];
                1081 / IN_WIDTH: ping_storage_data_865 <= (fillup_transition == 1'b1) ? i_input_data[1081 % IN_WIDTH] : ping_storage_data_865 ^ i_input_data[1081 % IN_WIDTH];
                default: ping_storage_data_865 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_865;
                endcase
            end else begin
                case (input_count)
                483 / IN_WIDTH: pong_storage_data_865 <= (fillup_transition == 1'b1) ? i_input_data[483 % IN_WIDTH] : pong_storage_data_865 ^ i_input_data[483 % IN_WIDTH];
                710 / IN_WIDTH: pong_storage_data_865 <= (fillup_transition == 1'b1) ? i_input_data[710 % IN_WIDTH] : pong_storage_data_865 ^ i_input_data[710 % IN_WIDTH];
                987 / IN_WIDTH: pong_storage_data_865 <= (fillup_transition == 1'b1) ? i_input_data[987 % IN_WIDTH] : pong_storage_data_865 ^ i_input_data[987 % IN_WIDTH];
                1081 / IN_WIDTH: pong_storage_data_865 <= (fillup_transition == 1'b1) ? i_input_data[1081 % IN_WIDTH] : pong_storage_data_865 ^ i_input_data[1081 % IN_WIDTH];
                default: pong_storage_data_865 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_865;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_865 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_865;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_865 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_865;
            end
        end
    end
end

logic ping_storage_data_866;
logic pong_storage_data_866;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_866 <= 1'b0;
        pong_storage_data_866 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                484 / IN_WIDTH: ping_storage_data_866 <= (fillup_transition == 1'b1) ? i_input_data[484 % IN_WIDTH] : ping_storage_data_866 ^ i_input_data[484 % IN_WIDTH];
                711 / IN_WIDTH: ping_storage_data_866 <= (fillup_transition == 1'b1) ? i_input_data[711 % IN_WIDTH] : ping_storage_data_866 ^ i_input_data[711 % IN_WIDTH];
                988 / IN_WIDTH: ping_storage_data_866 <= (fillup_transition == 1'b1) ? i_input_data[988 % IN_WIDTH] : ping_storage_data_866 ^ i_input_data[988 % IN_WIDTH];
                1082 / IN_WIDTH: ping_storage_data_866 <= (fillup_transition == 1'b1) ? i_input_data[1082 % IN_WIDTH] : ping_storage_data_866 ^ i_input_data[1082 % IN_WIDTH];
                default: ping_storage_data_866 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_866;
                endcase
            end else begin
                case (input_count)
                484 / IN_WIDTH: pong_storage_data_866 <= (fillup_transition == 1'b1) ? i_input_data[484 % IN_WIDTH] : pong_storage_data_866 ^ i_input_data[484 % IN_WIDTH];
                711 / IN_WIDTH: pong_storage_data_866 <= (fillup_transition == 1'b1) ? i_input_data[711 % IN_WIDTH] : pong_storage_data_866 ^ i_input_data[711 % IN_WIDTH];
                988 / IN_WIDTH: pong_storage_data_866 <= (fillup_transition == 1'b1) ? i_input_data[988 % IN_WIDTH] : pong_storage_data_866 ^ i_input_data[988 % IN_WIDTH];
                1082 / IN_WIDTH: pong_storage_data_866 <= (fillup_transition == 1'b1) ? i_input_data[1082 % IN_WIDTH] : pong_storage_data_866 ^ i_input_data[1082 % IN_WIDTH];
                default: pong_storage_data_866 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_866;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_866 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_866;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_866 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_866;
            end
        end
    end
end

logic ping_storage_data_867;
logic pong_storage_data_867;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_867 <= 1'b0;
        pong_storage_data_867 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                485 / IN_WIDTH: ping_storage_data_867 <= (fillup_transition == 1'b1) ? i_input_data[485 % IN_WIDTH] : ping_storage_data_867 ^ i_input_data[485 % IN_WIDTH];
                712 / IN_WIDTH: ping_storage_data_867 <= (fillup_transition == 1'b1) ? i_input_data[712 % IN_WIDTH] : ping_storage_data_867 ^ i_input_data[712 % IN_WIDTH];
                989 / IN_WIDTH: ping_storage_data_867 <= (fillup_transition == 1'b1) ? i_input_data[989 % IN_WIDTH] : ping_storage_data_867 ^ i_input_data[989 % IN_WIDTH];
                1083 / IN_WIDTH: ping_storage_data_867 <= (fillup_transition == 1'b1) ? i_input_data[1083 % IN_WIDTH] : ping_storage_data_867 ^ i_input_data[1083 % IN_WIDTH];
                default: ping_storage_data_867 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_867;
                endcase
            end else begin
                case (input_count)
                485 / IN_WIDTH: pong_storage_data_867 <= (fillup_transition == 1'b1) ? i_input_data[485 % IN_WIDTH] : pong_storage_data_867 ^ i_input_data[485 % IN_WIDTH];
                712 / IN_WIDTH: pong_storage_data_867 <= (fillup_transition == 1'b1) ? i_input_data[712 % IN_WIDTH] : pong_storage_data_867 ^ i_input_data[712 % IN_WIDTH];
                989 / IN_WIDTH: pong_storage_data_867 <= (fillup_transition == 1'b1) ? i_input_data[989 % IN_WIDTH] : pong_storage_data_867 ^ i_input_data[989 % IN_WIDTH];
                1083 / IN_WIDTH: pong_storage_data_867 <= (fillup_transition == 1'b1) ? i_input_data[1083 % IN_WIDTH] : pong_storage_data_867 ^ i_input_data[1083 % IN_WIDTH];
                default: pong_storage_data_867 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_867;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_867 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_867;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_867 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_867;
            end
        end
    end
end

logic ping_storage_data_868;
logic pong_storage_data_868;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_868 <= 1'b0;
        pong_storage_data_868 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                486 / IN_WIDTH: ping_storage_data_868 <= (fillup_transition == 1'b1) ? i_input_data[486 % IN_WIDTH] : ping_storage_data_868 ^ i_input_data[486 % IN_WIDTH];
                713 / IN_WIDTH: ping_storage_data_868 <= (fillup_transition == 1'b1) ? i_input_data[713 % IN_WIDTH] : ping_storage_data_868 ^ i_input_data[713 % IN_WIDTH];
                990 / IN_WIDTH: ping_storage_data_868 <= (fillup_transition == 1'b1) ? i_input_data[990 % IN_WIDTH] : ping_storage_data_868 ^ i_input_data[990 % IN_WIDTH];
                1084 / IN_WIDTH: ping_storage_data_868 <= (fillup_transition == 1'b1) ? i_input_data[1084 % IN_WIDTH] : ping_storage_data_868 ^ i_input_data[1084 % IN_WIDTH];
                default: ping_storage_data_868 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_868;
                endcase
            end else begin
                case (input_count)
                486 / IN_WIDTH: pong_storage_data_868 <= (fillup_transition == 1'b1) ? i_input_data[486 % IN_WIDTH] : pong_storage_data_868 ^ i_input_data[486 % IN_WIDTH];
                713 / IN_WIDTH: pong_storage_data_868 <= (fillup_transition == 1'b1) ? i_input_data[713 % IN_WIDTH] : pong_storage_data_868 ^ i_input_data[713 % IN_WIDTH];
                990 / IN_WIDTH: pong_storage_data_868 <= (fillup_transition == 1'b1) ? i_input_data[990 % IN_WIDTH] : pong_storage_data_868 ^ i_input_data[990 % IN_WIDTH];
                1084 / IN_WIDTH: pong_storage_data_868 <= (fillup_transition == 1'b1) ? i_input_data[1084 % IN_WIDTH] : pong_storage_data_868 ^ i_input_data[1084 % IN_WIDTH];
                default: pong_storage_data_868 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_868;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_868 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_868;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_868 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_868;
            end
        end
    end
end

logic ping_storage_data_869;
logic pong_storage_data_869;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_869 <= 1'b0;
        pong_storage_data_869 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                487 / IN_WIDTH: ping_storage_data_869 <= (fillup_transition == 1'b1) ? i_input_data[487 % IN_WIDTH] : ping_storage_data_869 ^ i_input_data[487 % IN_WIDTH];
                714 / IN_WIDTH: ping_storage_data_869 <= (fillup_transition == 1'b1) ? i_input_data[714 % IN_WIDTH] : ping_storage_data_869 ^ i_input_data[714 % IN_WIDTH];
                991 / IN_WIDTH: ping_storage_data_869 <= (fillup_transition == 1'b1) ? i_input_data[991 % IN_WIDTH] : ping_storage_data_869 ^ i_input_data[991 % IN_WIDTH];
                1085 / IN_WIDTH: ping_storage_data_869 <= (fillup_transition == 1'b1) ? i_input_data[1085 % IN_WIDTH] : ping_storage_data_869 ^ i_input_data[1085 % IN_WIDTH];
                default: ping_storage_data_869 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_869;
                endcase
            end else begin
                case (input_count)
                487 / IN_WIDTH: pong_storage_data_869 <= (fillup_transition == 1'b1) ? i_input_data[487 % IN_WIDTH] : pong_storage_data_869 ^ i_input_data[487 % IN_WIDTH];
                714 / IN_WIDTH: pong_storage_data_869 <= (fillup_transition == 1'b1) ? i_input_data[714 % IN_WIDTH] : pong_storage_data_869 ^ i_input_data[714 % IN_WIDTH];
                991 / IN_WIDTH: pong_storage_data_869 <= (fillup_transition == 1'b1) ? i_input_data[991 % IN_WIDTH] : pong_storage_data_869 ^ i_input_data[991 % IN_WIDTH];
                1085 / IN_WIDTH: pong_storage_data_869 <= (fillup_transition == 1'b1) ? i_input_data[1085 % IN_WIDTH] : pong_storage_data_869 ^ i_input_data[1085 % IN_WIDTH];
                default: pong_storage_data_869 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_869;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_869 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_869;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_869 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_869;
            end
        end
    end
end

logic ping_storage_data_870;
logic pong_storage_data_870;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_870 <= 1'b0;
        pong_storage_data_870 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                488 / IN_WIDTH: ping_storage_data_870 <= (fillup_transition == 1'b1) ? i_input_data[488 % IN_WIDTH] : ping_storage_data_870 ^ i_input_data[488 % IN_WIDTH];
                715 / IN_WIDTH: ping_storage_data_870 <= (fillup_transition == 1'b1) ? i_input_data[715 % IN_WIDTH] : ping_storage_data_870 ^ i_input_data[715 % IN_WIDTH];
                992 / IN_WIDTH: ping_storage_data_870 <= (fillup_transition == 1'b1) ? i_input_data[992 % IN_WIDTH] : ping_storage_data_870 ^ i_input_data[992 % IN_WIDTH];
                1086 / IN_WIDTH: ping_storage_data_870 <= (fillup_transition == 1'b1) ? i_input_data[1086 % IN_WIDTH] : ping_storage_data_870 ^ i_input_data[1086 % IN_WIDTH];
                default: ping_storage_data_870 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_870;
                endcase
            end else begin
                case (input_count)
                488 / IN_WIDTH: pong_storage_data_870 <= (fillup_transition == 1'b1) ? i_input_data[488 % IN_WIDTH] : pong_storage_data_870 ^ i_input_data[488 % IN_WIDTH];
                715 / IN_WIDTH: pong_storage_data_870 <= (fillup_transition == 1'b1) ? i_input_data[715 % IN_WIDTH] : pong_storage_data_870 ^ i_input_data[715 % IN_WIDTH];
                992 / IN_WIDTH: pong_storage_data_870 <= (fillup_transition == 1'b1) ? i_input_data[992 % IN_WIDTH] : pong_storage_data_870 ^ i_input_data[992 % IN_WIDTH];
                1086 / IN_WIDTH: pong_storage_data_870 <= (fillup_transition == 1'b1) ? i_input_data[1086 % IN_WIDTH] : pong_storage_data_870 ^ i_input_data[1086 % IN_WIDTH];
                default: pong_storage_data_870 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_870;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_870 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_870;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_870 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_870;
            end
        end
    end
end

logic ping_storage_data_871;
logic pong_storage_data_871;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_871 <= 1'b0;
        pong_storage_data_871 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                489 / IN_WIDTH: ping_storage_data_871 <= (fillup_transition == 1'b1) ? i_input_data[489 % IN_WIDTH] : ping_storage_data_871 ^ i_input_data[489 % IN_WIDTH];
                716 / IN_WIDTH: ping_storage_data_871 <= (fillup_transition == 1'b1) ? i_input_data[716 % IN_WIDTH] : ping_storage_data_871 ^ i_input_data[716 % IN_WIDTH];
                993 / IN_WIDTH: ping_storage_data_871 <= (fillup_transition == 1'b1) ? i_input_data[993 % IN_WIDTH] : ping_storage_data_871 ^ i_input_data[993 % IN_WIDTH];
                1087 / IN_WIDTH: ping_storage_data_871 <= (fillup_transition == 1'b1) ? i_input_data[1087 % IN_WIDTH] : ping_storage_data_871 ^ i_input_data[1087 % IN_WIDTH];
                default: ping_storage_data_871 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_871;
                endcase
            end else begin
                case (input_count)
                489 / IN_WIDTH: pong_storage_data_871 <= (fillup_transition == 1'b1) ? i_input_data[489 % IN_WIDTH] : pong_storage_data_871 ^ i_input_data[489 % IN_WIDTH];
                716 / IN_WIDTH: pong_storage_data_871 <= (fillup_transition == 1'b1) ? i_input_data[716 % IN_WIDTH] : pong_storage_data_871 ^ i_input_data[716 % IN_WIDTH];
                993 / IN_WIDTH: pong_storage_data_871 <= (fillup_transition == 1'b1) ? i_input_data[993 % IN_WIDTH] : pong_storage_data_871 ^ i_input_data[993 % IN_WIDTH];
                1087 / IN_WIDTH: pong_storage_data_871 <= (fillup_transition == 1'b1) ? i_input_data[1087 % IN_WIDTH] : pong_storage_data_871 ^ i_input_data[1087 % IN_WIDTH];
                default: pong_storage_data_871 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_871;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_871 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_871;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_871 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_871;
            end
        end
    end
end

logic ping_storage_data_872;
logic pong_storage_data_872;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_872 <= 1'b0;
        pong_storage_data_872 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                490 / IN_WIDTH: ping_storage_data_872 <= (fillup_transition == 1'b1) ? i_input_data[490 % IN_WIDTH] : ping_storage_data_872 ^ i_input_data[490 % IN_WIDTH];
                717 / IN_WIDTH: ping_storage_data_872 <= (fillup_transition == 1'b1) ? i_input_data[717 % IN_WIDTH] : ping_storage_data_872 ^ i_input_data[717 % IN_WIDTH];
                994 / IN_WIDTH: ping_storage_data_872 <= (fillup_transition == 1'b1) ? i_input_data[994 % IN_WIDTH] : ping_storage_data_872 ^ i_input_data[994 % IN_WIDTH];
                1088 / IN_WIDTH: ping_storage_data_872 <= (fillup_transition == 1'b1) ? i_input_data[1088 % IN_WIDTH] : ping_storage_data_872 ^ i_input_data[1088 % IN_WIDTH];
                default: ping_storage_data_872 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_872;
                endcase
            end else begin
                case (input_count)
                490 / IN_WIDTH: pong_storage_data_872 <= (fillup_transition == 1'b1) ? i_input_data[490 % IN_WIDTH] : pong_storage_data_872 ^ i_input_data[490 % IN_WIDTH];
                717 / IN_WIDTH: pong_storage_data_872 <= (fillup_transition == 1'b1) ? i_input_data[717 % IN_WIDTH] : pong_storage_data_872 ^ i_input_data[717 % IN_WIDTH];
                994 / IN_WIDTH: pong_storage_data_872 <= (fillup_transition == 1'b1) ? i_input_data[994 % IN_WIDTH] : pong_storage_data_872 ^ i_input_data[994 % IN_WIDTH];
                1088 / IN_WIDTH: pong_storage_data_872 <= (fillup_transition == 1'b1) ? i_input_data[1088 % IN_WIDTH] : pong_storage_data_872 ^ i_input_data[1088 % IN_WIDTH];
                default: pong_storage_data_872 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_872;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_872 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_872;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_872 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_872;
            end
        end
    end
end

logic ping_storage_data_873;
logic pong_storage_data_873;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_873 <= 1'b0;
        pong_storage_data_873 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                491 / IN_WIDTH: ping_storage_data_873 <= (fillup_transition == 1'b1) ? i_input_data[491 % IN_WIDTH] : ping_storage_data_873 ^ i_input_data[491 % IN_WIDTH];
                718 / IN_WIDTH: ping_storage_data_873 <= (fillup_transition == 1'b1) ? i_input_data[718 % IN_WIDTH] : ping_storage_data_873 ^ i_input_data[718 % IN_WIDTH];
                995 / IN_WIDTH: ping_storage_data_873 <= (fillup_transition == 1'b1) ? i_input_data[995 % IN_WIDTH] : ping_storage_data_873 ^ i_input_data[995 % IN_WIDTH];
                1089 / IN_WIDTH: ping_storage_data_873 <= (fillup_transition == 1'b1) ? i_input_data[1089 % IN_WIDTH] : ping_storage_data_873 ^ i_input_data[1089 % IN_WIDTH];
                default: ping_storage_data_873 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_873;
                endcase
            end else begin
                case (input_count)
                491 / IN_WIDTH: pong_storage_data_873 <= (fillup_transition == 1'b1) ? i_input_data[491 % IN_WIDTH] : pong_storage_data_873 ^ i_input_data[491 % IN_WIDTH];
                718 / IN_WIDTH: pong_storage_data_873 <= (fillup_transition == 1'b1) ? i_input_data[718 % IN_WIDTH] : pong_storage_data_873 ^ i_input_data[718 % IN_WIDTH];
                995 / IN_WIDTH: pong_storage_data_873 <= (fillup_transition == 1'b1) ? i_input_data[995 % IN_WIDTH] : pong_storage_data_873 ^ i_input_data[995 % IN_WIDTH];
                1089 / IN_WIDTH: pong_storage_data_873 <= (fillup_transition == 1'b1) ? i_input_data[1089 % IN_WIDTH] : pong_storage_data_873 ^ i_input_data[1089 % IN_WIDTH];
                default: pong_storage_data_873 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_873;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_873 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_873;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_873 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_873;
            end
        end
    end
end

logic ping_storage_data_874;
logic pong_storage_data_874;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_874 <= 1'b0;
        pong_storage_data_874 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                492 / IN_WIDTH: ping_storage_data_874 <= (fillup_transition == 1'b1) ? i_input_data[492 % IN_WIDTH] : ping_storage_data_874 ^ i_input_data[492 % IN_WIDTH];
                719 / IN_WIDTH: ping_storage_data_874 <= (fillup_transition == 1'b1) ? i_input_data[719 % IN_WIDTH] : ping_storage_data_874 ^ i_input_data[719 % IN_WIDTH];
                996 / IN_WIDTH: ping_storage_data_874 <= (fillup_transition == 1'b1) ? i_input_data[996 % IN_WIDTH] : ping_storage_data_874 ^ i_input_data[996 % IN_WIDTH];
                1090 / IN_WIDTH: ping_storage_data_874 <= (fillup_transition == 1'b1) ? i_input_data[1090 % IN_WIDTH] : ping_storage_data_874 ^ i_input_data[1090 % IN_WIDTH];
                default: ping_storage_data_874 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_874;
                endcase
            end else begin
                case (input_count)
                492 / IN_WIDTH: pong_storage_data_874 <= (fillup_transition == 1'b1) ? i_input_data[492 % IN_WIDTH] : pong_storage_data_874 ^ i_input_data[492 % IN_WIDTH];
                719 / IN_WIDTH: pong_storage_data_874 <= (fillup_transition == 1'b1) ? i_input_data[719 % IN_WIDTH] : pong_storage_data_874 ^ i_input_data[719 % IN_WIDTH];
                996 / IN_WIDTH: pong_storage_data_874 <= (fillup_transition == 1'b1) ? i_input_data[996 % IN_WIDTH] : pong_storage_data_874 ^ i_input_data[996 % IN_WIDTH];
                1090 / IN_WIDTH: pong_storage_data_874 <= (fillup_transition == 1'b1) ? i_input_data[1090 % IN_WIDTH] : pong_storage_data_874 ^ i_input_data[1090 % IN_WIDTH];
                default: pong_storage_data_874 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_874;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_874 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_874;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_874 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_874;
            end
        end
    end
end

logic ping_storage_data_875;
logic pong_storage_data_875;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_875 <= 1'b0;
        pong_storage_data_875 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                493 / IN_WIDTH: ping_storage_data_875 <= (fillup_transition == 1'b1) ? i_input_data[493 % IN_WIDTH] : ping_storage_data_875 ^ i_input_data[493 % IN_WIDTH];
                720 / IN_WIDTH: ping_storage_data_875 <= (fillup_transition == 1'b1) ? i_input_data[720 % IN_WIDTH] : ping_storage_data_875 ^ i_input_data[720 % IN_WIDTH];
                997 / IN_WIDTH: ping_storage_data_875 <= (fillup_transition == 1'b1) ? i_input_data[997 % IN_WIDTH] : ping_storage_data_875 ^ i_input_data[997 % IN_WIDTH];
                1091 / IN_WIDTH: ping_storage_data_875 <= (fillup_transition == 1'b1) ? i_input_data[1091 % IN_WIDTH] : ping_storage_data_875 ^ i_input_data[1091 % IN_WIDTH];
                default: ping_storage_data_875 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_875;
                endcase
            end else begin
                case (input_count)
                493 / IN_WIDTH: pong_storage_data_875 <= (fillup_transition == 1'b1) ? i_input_data[493 % IN_WIDTH] : pong_storage_data_875 ^ i_input_data[493 % IN_WIDTH];
                720 / IN_WIDTH: pong_storage_data_875 <= (fillup_transition == 1'b1) ? i_input_data[720 % IN_WIDTH] : pong_storage_data_875 ^ i_input_data[720 % IN_WIDTH];
                997 / IN_WIDTH: pong_storage_data_875 <= (fillup_transition == 1'b1) ? i_input_data[997 % IN_WIDTH] : pong_storage_data_875 ^ i_input_data[997 % IN_WIDTH];
                1091 / IN_WIDTH: pong_storage_data_875 <= (fillup_transition == 1'b1) ? i_input_data[1091 % IN_WIDTH] : pong_storage_data_875 ^ i_input_data[1091 % IN_WIDTH];
                default: pong_storage_data_875 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_875;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_875 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_875;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_875 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_875;
            end
        end
    end
end

logic ping_storage_data_876;
logic pong_storage_data_876;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_876 <= 1'b0;
        pong_storage_data_876 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                494 / IN_WIDTH: ping_storage_data_876 <= (fillup_transition == 1'b1) ? i_input_data[494 % IN_WIDTH] : ping_storage_data_876 ^ i_input_data[494 % IN_WIDTH];
                721 / IN_WIDTH: ping_storage_data_876 <= (fillup_transition == 1'b1) ? i_input_data[721 % IN_WIDTH] : ping_storage_data_876 ^ i_input_data[721 % IN_WIDTH];
                998 / IN_WIDTH: ping_storage_data_876 <= (fillup_transition == 1'b1) ? i_input_data[998 % IN_WIDTH] : ping_storage_data_876 ^ i_input_data[998 % IN_WIDTH];
                1092 / IN_WIDTH: ping_storage_data_876 <= (fillup_transition == 1'b1) ? i_input_data[1092 % IN_WIDTH] : ping_storage_data_876 ^ i_input_data[1092 % IN_WIDTH];
                default: ping_storage_data_876 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_876;
                endcase
            end else begin
                case (input_count)
                494 / IN_WIDTH: pong_storage_data_876 <= (fillup_transition == 1'b1) ? i_input_data[494 % IN_WIDTH] : pong_storage_data_876 ^ i_input_data[494 % IN_WIDTH];
                721 / IN_WIDTH: pong_storage_data_876 <= (fillup_transition == 1'b1) ? i_input_data[721 % IN_WIDTH] : pong_storage_data_876 ^ i_input_data[721 % IN_WIDTH];
                998 / IN_WIDTH: pong_storage_data_876 <= (fillup_transition == 1'b1) ? i_input_data[998 % IN_WIDTH] : pong_storage_data_876 ^ i_input_data[998 % IN_WIDTH];
                1092 / IN_WIDTH: pong_storage_data_876 <= (fillup_transition == 1'b1) ? i_input_data[1092 % IN_WIDTH] : pong_storage_data_876 ^ i_input_data[1092 % IN_WIDTH];
                default: pong_storage_data_876 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_876;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_876 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_876;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_876 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_876;
            end
        end
    end
end

logic ping_storage_data_877;
logic pong_storage_data_877;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_877 <= 1'b0;
        pong_storage_data_877 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                495 / IN_WIDTH: ping_storage_data_877 <= (fillup_transition == 1'b1) ? i_input_data[495 % IN_WIDTH] : ping_storage_data_877 ^ i_input_data[495 % IN_WIDTH];
                722 / IN_WIDTH: ping_storage_data_877 <= (fillup_transition == 1'b1) ? i_input_data[722 % IN_WIDTH] : ping_storage_data_877 ^ i_input_data[722 % IN_WIDTH];
                999 / IN_WIDTH: ping_storage_data_877 <= (fillup_transition == 1'b1) ? i_input_data[999 % IN_WIDTH] : ping_storage_data_877 ^ i_input_data[999 % IN_WIDTH];
                1093 / IN_WIDTH: ping_storage_data_877 <= (fillup_transition == 1'b1) ? i_input_data[1093 % IN_WIDTH] : ping_storage_data_877 ^ i_input_data[1093 % IN_WIDTH];
                default: ping_storage_data_877 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_877;
                endcase
            end else begin
                case (input_count)
                495 / IN_WIDTH: pong_storage_data_877 <= (fillup_transition == 1'b1) ? i_input_data[495 % IN_WIDTH] : pong_storage_data_877 ^ i_input_data[495 % IN_WIDTH];
                722 / IN_WIDTH: pong_storage_data_877 <= (fillup_transition == 1'b1) ? i_input_data[722 % IN_WIDTH] : pong_storage_data_877 ^ i_input_data[722 % IN_WIDTH];
                999 / IN_WIDTH: pong_storage_data_877 <= (fillup_transition == 1'b1) ? i_input_data[999 % IN_WIDTH] : pong_storage_data_877 ^ i_input_data[999 % IN_WIDTH];
                1093 / IN_WIDTH: pong_storage_data_877 <= (fillup_transition == 1'b1) ? i_input_data[1093 % IN_WIDTH] : pong_storage_data_877 ^ i_input_data[1093 % IN_WIDTH];
                default: pong_storage_data_877 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_877;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_877 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_877;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_877 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_877;
            end
        end
    end
end

logic ping_storage_data_878;
logic pong_storage_data_878;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_878 <= 1'b0;
        pong_storage_data_878 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                496 / IN_WIDTH: ping_storage_data_878 <= (fillup_transition == 1'b1) ? i_input_data[496 % IN_WIDTH] : ping_storage_data_878 ^ i_input_data[496 % IN_WIDTH];
                723 / IN_WIDTH: ping_storage_data_878 <= (fillup_transition == 1'b1) ? i_input_data[723 % IN_WIDTH] : ping_storage_data_878 ^ i_input_data[723 % IN_WIDTH];
                1000 / IN_WIDTH: ping_storage_data_878 <= (fillup_transition == 1'b1) ? i_input_data[1000 % IN_WIDTH] : ping_storage_data_878 ^ i_input_data[1000 % IN_WIDTH];
                1094 / IN_WIDTH: ping_storage_data_878 <= (fillup_transition == 1'b1) ? i_input_data[1094 % IN_WIDTH] : ping_storage_data_878 ^ i_input_data[1094 % IN_WIDTH];
                default: ping_storage_data_878 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_878;
                endcase
            end else begin
                case (input_count)
                496 / IN_WIDTH: pong_storage_data_878 <= (fillup_transition == 1'b1) ? i_input_data[496 % IN_WIDTH] : pong_storage_data_878 ^ i_input_data[496 % IN_WIDTH];
                723 / IN_WIDTH: pong_storage_data_878 <= (fillup_transition == 1'b1) ? i_input_data[723 % IN_WIDTH] : pong_storage_data_878 ^ i_input_data[723 % IN_WIDTH];
                1000 / IN_WIDTH: pong_storage_data_878 <= (fillup_transition == 1'b1) ? i_input_data[1000 % IN_WIDTH] : pong_storage_data_878 ^ i_input_data[1000 % IN_WIDTH];
                1094 / IN_WIDTH: pong_storage_data_878 <= (fillup_transition == 1'b1) ? i_input_data[1094 % IN_WIDTH] : pong_storage_data_878 ^ i_input_data[1094 % IN_WIDTH];
                default: pong_storage_data_878 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_878;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_878 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_878;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_878 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_878;
            end
        end
    end
end

logic ping_storage_data_879;
logic pong_storage_data_879;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_879 <= 1'b0;
        pong_storage_data_879 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                497 / IN_WIDTH: ping_storage_data_879 <= (fillup_transition == 1'b1) ? i_input_data[497 % IN_WIDTH] : ping_storage_data_879 ^ i_input_data[497 % IN_WIDTH];
                724 / IN_WIDTH: ping_storage_data_879 <= (fillup_transition == 1'b1) ? i_input_data[724 % IN_WIDTH] : ping_storage_data_879 ^ i_input_data[724 % IN_WIDTH];
                1001 / IN_WIDTH: ping_storage_data_879 <= (fillup_transition == 1'b1) ? i_input_data[1001 % IN_WIDTH] : ping_storage_data_879 ^ i_input_data[1001 % IN_WIDTH];
                1095 / IN_WIDTH: ping_storage_data_879 <= (fillup_transition == 1'b1) ? i_input_data[1095 % IN_WIDTH] : ping_storage_data_879 ^ i_input_data[1095 % IN_WIDTH];
                default: ping_storage_data_879 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_879;
                endcase
            end else begin
                case (input_count)
                497 / IN_WIDTH: pong_storage_data_879 <= (fillup_transition == 1'b1) ? i_input_data[497 % IN_WIDTH] : pong_storage_data_879 ^ i_input_data[497 % IN_WIDTH];
                724 / IN_WIDTH: pong_storage_data_879 <= (fillup_transition == 1'b1) ? i_input_data[724 % IN_WIDTH] : pong_storage_data_879 ^ i_input_data[724 % IN_WIDTH];
                1001 / IN_WIDTH: pong_storage_data_879 <= (fillup_transition == 1'b1) ? i_input_data[1001 % IN_WIDTH] : pong_storage_data_879 ^ i_input_data[1001 % IN_WIDTH];
                1095 / IN_WIDTH: pong_storage_data_879 <= (fillup_transition == 1'b1) ? i_input_data[1095 % IN_WIDTH] : pong_storage_data_879 ^ i_input_data[1095 % IN_WIDTH];
                default: pong_storage_data_879 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_879;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_879 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_879;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_879 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_879;
            end
        end
    end
end

logic ping_storage_data_880;
logic pong_storage_data_880;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_880 <= 1'b0;
        pong_storage_data_880 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                498 / IN_WIDTH: ping_storage_data_880 <= (fillup_transition == 1'b1) ? i_input_data[498 % IN_WIDTH] : ping_storage_data_880 ^ i_input_data[498 % IN_WIDTH];
                725 / IN_WIDTH: ping_storage_data_880 <= (fillup_transition == 1'b1) ? i_input_data[725 % IN_WIDTH] : ping_storage_data_880 ^ i_input_data[725 % IN_WIDTH];
                1002 / IN_WIDTH: ping_storage_data_880 <= (fillup_transition == 1'b1) ? i_input_data[1002 % IN_WIDTH] : ping_storage_data_880 ^ i_input_data[1002 % IN_WIDTH];
                1096 / IN_WIDTH: ping_storage_data_880 <= (fillup_transition == 1'b1) ? i_input_data[1096 % IN_WIDTH] : ping_storage_data_880 ^ i_input_data[1096 % IN_WIDTH];
                default: ping_storage_data_880 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_880;
                endcase
            end else begin
                case (input_count)
                498 / IN_WIDTH: pong_storage_data_880 <= (fillup_transition == 1'b1) ? i_input_data[498 % IN_WIDTH] : pong_storage_data_880 ^ i_input_data[498 % IN_WIDTH];
                725 / IN_WIDTH: pong_storage_data_880 <= (fillup_transition == 1'b1) ? i_input_data[725 % IN_WIDTH] : pong_storage_data_880 ^ i_input_data[725 % IN_WIDTH];
                1002 / IN_WIDTH: pong_storage_data_880 <= (fillup_transition == 1'b1) ? i_input_data[1002 % IN_WIDTH] : pong_storage_data_880 ^ i_input_data[1002 % IN_WIDTH];
                1096 / IN_WIDTH: pong_storage_data_880 <= (fillup_transition == 1'b1) ? i_input_data[1096 % IN_WIDTH] : pong_storage_data_880 ^ i_input_data[1096 % IN_WIDTH];
                default: pong_storage_data_880 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_880;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_880 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_880;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_880 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_880;
            end
        end
    end
end

logic ping_storage_data_881;
logic pong_storage_data_881;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_881 <= 1'b0;
        pong_storage_data_881 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                499 / IN_WIDTH: ping_storage_data_881 <= (fillup_transition == 1'b1) ? i_input_data[499 % IN_WIDTH] : ping_storage_data_881 ^ i_input_data[499 % IN_WIDTH];
                726 / IN_WIDTH: ping_storage_data_881 <= (fillup_transition == 1'b1) ? i_input_data[726 % IN_WIDTH] : ping_storage_data_881 ^ i_input_data[726 % IN_WIDTH];
                1003 / IN_WIDTH: ping_storage_data_881 <= (fillup_transition == 1'b1) ? i_input_data[1003 % IN_WIDTH] : ping_storage_data_881 ^ i_input_data[1003 % IN_WIDTH];
                1097 / IN_WIDTH: ping_storage_data_881 <= (fillup_transition == 1'b1) ? i_input_data[1097 % IN_WIDTH] : ping_storage_data_881 ^ i_input_data[1097 % IN_WIDTH];
                default: ping_storage_data_881 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_881;
                endcase
            end else begin
                case (input_count)
                499 / IN_WIDTH: pong_storage_data_881 <= (fillup_transition == 1'b1) ? i_input_data[499 % IN_WIDTH] : pong_storage_data_881 ^ i_input_data[499 % IN_WIDTH];
                726 / IN_WIDTH: pong_storage_data_881 <= (fillup_transition == 1'b1) ? i_input_data[726 % IN_WIDTH] : pong_storage_data_881 ^ i_input_data[726 % IN_WIDTH];
                1003 / IN_WIDTH: pong_storage_data_881 <= (fillup_transition == 1'b1) ? i_input_data[1003 % IN_WIDTH] : pong_storage_data_881 ^ i_input_data[1003 % IN_WIDTH];
                1097 / IN_WIDTH: pong_storage_data_881 <= (fillup_transition == 1'b1) ? i_input_data[1097 % IN_WIDTH] : pong_storage_data_881 ^ i_input_data[1097 % IN_WIDTH];
                default: pong_storage_data_881 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_881;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_881 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_881;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_881 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_881;
            end
        end
    end
end

logic ping_storage_data_882;
logic pong_storage_data_882;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_882 <= 1'b0;
        pong_storage_data_882 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                500 / IN_WIDTH: ping_storage_data_882 <= (fillup_transition == 1'b1) ? i_input_data[500 % IN_WIDTH] : ping_storage_data_882 ^ i_input_data[500 % IN_WIDTH];
                727 / IN_WIDTH: ping_storage_data_882 <= (fillup_transition == 1'b1) ? i_input_data[727 % IN_WIDTH] : ping_storage_data_882 ^ i_input_data[727 % IN_WIDTH];
                1004 / IN_WIDTH: ping_storage_data_882 <= (fillup_transition == 1'b1) ? i_input_data[1004 % IN_WIDTH] : ping_storage_data_882 ^ i_input_data[1004 % IN_WIDTH];
                1098 / IN_WIDTH: ping_storage_data_882 <= (fillup_transition == 1'b1) ? i_input_data[1098 % IN_WIDTH] : ping_storage_data_882 ^ i_input_data[1098 % IN_WIDTH];
                default: ping_storage_data_882 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_882;
                endcase
            end else begin
                case (input_count)
                500 / IN_WIDTH: pong_storage_data_882 <= (fillup_transition == 1'b1) ? i_input_data[500 % IN_WIDTH] : pong_storage_data_882 ^ i_input_data[500 % IN_WIDTH];
                727 / IN_WIDTH: pong_storage_data_882 <= (fillup_transition == 1'b1) ? i_input_data[727 % IN_WIDTH] : pong_storage_data_882 ^ i_input_data[727 % IN_WIDTH];
                1004 / IN_WIDTH: pong_storage_data_882 <= (fillup_transition == 1'b1) ? i_input_data[1004 % IN_WIDTH] : pong_storage_data_882 ^ i_input_data[1004 % IN_WIDTH];
                1098 / IN_WIDTH: pong_storage_data_882 <= (fillup_transition == 1'b1) ? i_input_data[1098 % IN_WIDTH] : pong_storage_data_882 ^ i_input_data[1098 % IN_WIDTH];
                default: pong_storage_data_882 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_882;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_882 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_882;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_882 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_882;
            end
        end
    end
end

logic ping_storage_data_883;
logic pong_storage_data_883;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_883 <= 1'b0;
        pong_storage_data_883 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                501 / IN_WIDTH: ping_storage_data_883 <= (fillup_transition == 1'b1) ? i_input_data[501 % IN_WIDTH] : ping_storage_data_883 ^ i_input_data[501 % IN_WIDTH];
                728 / IN_WIDTH: ping_storage_data_883 <= (fillup_transition == 1'b1) ? i_input_data[728 % IN_WIDTH] : ping_storage_data_883 ^ i_input_data[728 % IN_WIDTH];
                1005 / IN_WIDTH: ping_storage_data_883 <= (fillup_transition == 1'b1) ? i_input_data[1005 % IN_WIDTH] : ping_storage_data_883 ^ i_input_data[1005 % IN_WIDTH];
                1099 / IN_WIDTH: ping_storage_data_883 <= (fillup_transition == 1'b1) ? i_input_data[1099 % IN_WIDTH] : ping_storage_data_883 ^ i_input_data[1099 % IN_WIDTH];
                default: ping_storage_data_883 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_883;
                endcase
            end else begin
                case (input_count)
                501 / IN_WIDTH: pong_storage_data_883 <= (fillup_transition == 1'b1) ? i_input_data[501 % IN_WIDTH] : pong_storage_data_883 ^ i_input_data[501 % IN_WIDTH];
                728 / IN_WIDTH: pong_storage_data_883 <= (fillup_transition == 1'b1) ? i_input_data[728 % IN_WIDTH] : pong_storage_data_883 ^ i_input_data[728 % IN_WIDTH];
                1005 / IN_WIDTH: pong_storage_data_883 <= (fillup_transition == 1'b1) ? i_input_data[1005 % IN_WIDTH] : pong_storage_data_883 ^ i_input_data[1005 % IN_WIDTH];
                1099 / IN_WIDTH: pong_storage_data_883 <= (fillup_transition == 1'b1) ? i_input_data[1099 % IN_WIDTH] : pong_storage_data_883 ^ i_input_data[1099 % IN_WIDTH];
                default: pong_storage_data_883 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_883;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_883 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_883;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_883 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_883;
            end
        end
    end
end

logic ping_storage_data_884;
logic pong_storage_data_884;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_884 <= 1'b0;
        pong_storage_data_884 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                502 / IN_WIDTH: ping_storage_data_884 <= (fillup_transition == 1'b1) ? i_input_data[502 % IN_WIDTH] : ping_storage_data_884 ^ i_input_data[502 % IN_WIDTH];
                729 / IN_WIDTH: ping_storage_data_884 <= (fillup_transition == 1'b1) ? i_input_data[729 % IN_WIDTH] : ping_storage_data_884 ^ i_input_data[729 % IN_WIDTH];
                1006 / IN_WIDTH: ping_storage_data_884 <= (fillup_transition == 1'b1) ? i_input_data[1006 % IN_WIDTH] : ping_storage_data_884 ^ i_input_data[1006 % IN_WIDTH];
                1100 / IN_WIDTH: ping_storage_data_884 <= (fillup_transition == 1'b1) ? i_input_data[1100 % IN_WIDTH] : ping_storage_data_884 ^ i_input_data[1100 % IN_WIDTH];
                default: ping_storage_data_884 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_884;
                endcase
            end else begin
                case (input_count)
                502 / IN_WIDTH: pong_storage_data_884 <= (fillup_transition == 1'b1) ? i_input_data[502 % IN_WIDTH] : pong_storage_data_884 ^ i_input_data[502 % IN_WIDTH];
                729 / IN_WIDTH: pong_storage_data_884 <= (fillup_transition == 1'b1) ? i_input_data[729 % IN_WIDTH] : pong_storage_data_884 ^ i_input_data[729 % IN_WIDTH];
                1006 / IN_WIDTH: pong_storage_data_884 <= (fillup_transition == 1'b1) ? i_input_data[1006 % IN_WIDTH] : pong_storage_data_884 ^ i_input_data[1006 % IN_WIDTH];
                1100 / IN_WIDTH: pong_storage_data_884 <= (fillup_transition == 1'b1) ? i_input_data[1100 % IN_WIDTH] : pong_storage_data_884 ^ i_input_data[1100 % IN_WIDTH];
                default: pong_storage_data_884 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_884;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_884 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_884;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_884 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_884;
            end
        end
    end
end

logic ping_storage_data_885;
logic pong_storage_data_885;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_885 <= 1'b0;
        pong_storage_data_885 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                503 / IN_WIDTH: ping_storage_data_885 <= (fillup_transition == 1'b1) ? i_input_data[503 % IN_WIDTH] : ping_storage_data_885 ^ i_input_data[503 % IN_WIDTH];
                730 / IN_WIDTH: ping_storage_data_885 <= (fillup_transition == 1'b1) ? i_input_data[730 % IN_WIDTH] : ping_storage_data_885 ^ i_input_data[730 % IN_WIDTH];
                1007 / IN_WIDTH: ping_storage_data_885 <= (fillup_transition == 1'b1) ? i_input_data[1007 % IN_WIDTH] : ping_storage_data_885 ^ i_input_data[1007 % IN_WIDTH];
                1101 / IN_WIDTH: ping_storage_data_885 <= (fillup_transition == 1'b1) ? i_input_data[1101 % IN_WIDTH] : ping_storage_data_885 ^ i_input_data[1101 % IN_WIDTH];
                default: ping_storage_data_885 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_885;
                endcase
            end else begin
                case (input_count)
                503 / IN_WIDTH: pong_storage_data_885 <= (fillup_transition == 1'b1) ? i_input_data[503 % IN_WIDTH] : pong_storage_data_885 ^ i_input_data[503 % IN_WIDTH];
                730 / IN_WIDTH: pong_storage_data_885 <= (fillup_transition == 1'b1) ? i_input_data[730 % IN_WIDTH] : pong_storage_data_885 ^ i_input_data[730 % IN_WIDTH];
                1007 / IN_WIDTH: pong_storage_data_885 <= (fillup_transition == 1'b1) ? i_input_data[1007 % IN_WIDTH] : pong_storage_data_885 ^ i_input_data[1007 % IN_WIDTH];
                1101 / IN_WIDTH: pong_storage_data_885 <= (fillup_transition == 1'b1) ? i_input_data[1101 % IN_WIDTH] : pong_storage_data_885 ^ i_input_data[1101 % IN_WIDTH];
                default: pong_storage_data_885 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_885;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_885 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_885;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_885 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_885;
            end
        end
    end
end

logic ping_storage_data_886;
logic pong_storage_data_886;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_886 <= 1'b0;
        pong_storage_data_886 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                504 / IN_WIDTH: ping_storage_data_886 <= (fillup_transition == 1'b1) ? i_input_data[504 % IN_WIDTH] : ping_storage_data_886 ^ i_input_data[504 % IN_WIDTH];
                731 / IN_WIDTH: ping_storage_data_886 <= (fillup_transition == 1'b1) ? i_input_data[731 % IN_WIDTH] : ping_storage_data_886 ^ i_input_data[731 % IN_WIDTH];
                1008 / IN_WIDTH: ping_storage_data_886 <= (fillup_transition == 1'b1) ? i_input_data[1008 % IN_WIDTH] : ping_storage_data_886 ^ i_input_data[1008 % IN_WIDTH];
                1102 / IN_WIDTH: ping_storage_data_886 <= (fillup_transition == 1'b1) ? i_input_data[1102 % IN_WIDTH] : ping_storage_data_886 ^ i_input_data[1102 % IN_WIDTH];
                default: ping_storage_data_886 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_886;
                endcase
            end else begin
                case (input_count)
                504 / IN_WIDTH: pong_storage_data_886 <= (fillup_transition == 1'b1) ? i_input_data[504 % IN_WIDTH] : pong_storage_data_886 ^ i_input_data[504 % IN_WIDTH];
                731 / IN_WIDTH: pong_storage_data_886 <= (fillup_transition == 1'b1) ? i_input_data[731 % IN_WIDTH] : pong_storage_data_886 ^ i_input_data[731 % IN_WIDTH];
                1008 / IN_WIDTH: pong_storage_data_886 <= (fillup_transition == 1'b1) ? i_input_data[1008 % IN_WIDTH] : pong_storage_data_886 ^ i_input_data[1008 % IN_WIDTH];
                1102 / IN_WIDTH: pong_storage_data_886 <= (fillup_transition == 1'b1) ? i_input_data[1102 % IN_WIDTH] : pong_storage_data_886 ^ i_input_data[1102 % IN_WIDTH];
                default: pong_storage_data_886 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_886;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_886 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_886;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_886 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_886;
            end
        end
    end
end

logic ping_storage_data_887;
logic pong_storage_data_887;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_887 <= 1'b0;
        pong_storage_data_887 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                505 / IN_WIDTH: ping_storage_data_887 <= (fillup_transition == 1'b1) ? i_input_data[505 % IN_WIDTH] : ping_storage_data_887 ^ i_input_data[505 % IN_WIDTH];
                732 / IN_WIDTH: ping_storage_data_887 <= (fillup_transition == 1'b1) ? i_input_data[732 % IN_WIDTH] : ping_storage_data_887 ^ i_input_data[732 % IN_WIDTH];
                1009 / IN_WIDTH: ping_storage_data_887 <= (fillup_transition == 1'b1) ? i_input_data[1009 % IN_WIDTH] : ping_storage_data_887 ^ i_input_data[1009 % IN_WIDTH];
                1103 / IN_WIDTH: ping_storage_data_887 <= (fillup_transition == 1'b1) ? i_input_data[1103 % IN_WIDTH] : ping_storage_data_887 ^ i_input_data[1103 % IN_WIDTH];
                default: ping_storage_data_887 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_887;
                endcase
            end else begin
                case (input_count)
                505 / IN_WIDTH: pong_storage_data_887 <= (fillup_transition == 1'b1) ? i_input_data[505 % IN_WIDTH] : pong_storage_data_887 ^ i_input_data[505 % IN_WIDTH];
                732 / IN_WIDTH: pong_storage_data_887 <= (fillup_transition == 1'b1) ? i_input_data[732 % IN_WIDTH] : pong_storage_data_887 ^ i_input_data[732 % IN_WIDTH];
                1009 / IN_WIDTH: pong_storage_data_887 <= (fillup_transition == 1'b1) ? i_input_data[1009 % IN_WIDTH] : pong_storage_data_887 ^ i_input_data[1009 % IN_WIDTH];
                1103 / IN_WIDTH: pong_storage_data_887 <= (fillup_transition == 1'b1) ? i_input_data[1103 % IN_WIDTH] : pong_storage_data_887 ^ i_input_data[1103 % IN_WIDTH];
                default: pong_storage_data_887 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_887;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_887 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_887;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_887 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_887;
            end
        end
    end
end

logic ping_storage_data_888;
logic pong_storage_data_888;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_888 <= 1'b0;
        pong_storage_data_888 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                506 / IN_WIDTH: ping_storage_data_888 <= (fillup_transition == 1'b1) ? i_input_data[506 % IN_WIDTH] : ping_storage_data_888 ^ i_input_data[506 % IN_WIDTH];
                733 / IN_WIDTH: ping_storage_data_888 <= (fillup_transition == 1'b1) ? i_input_data[733 % IN_WIDTH] : ping_storage_data_888 ^ i_input_data[733 % IN_WIDTH];
                1010 / IN_WIDTH: ping_storage_data_888 <= (fillup_transition == 1'b1) ? i_input_data[1010 % IN_WIDTH] : ping_storage_data_888 ^ i_input_data[1010 % IN_WIDTH];
                1104 / IN_WIDTH: ping_storage_data_888 <= (fillup_transition == 1'b1) ? i_input_data[1104 % IN_WIDTH] : ping_storage_data_888 ^ i_input_data[1104 % IN_WIDTH];
                default: ping_storage_data_888 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_888;
                endcase
            end else begin
                case (input_count)
                506 / IN_WIDTH: pong_storage_data_888 <= (fillup_transition == 1'b1) ? i_input_data[506 % IN_WIDTH] : pong_storage_data_888 ^ i_input_data[506 % IN_WIDTH];
                733 / IN_WIDTH: pong_storage_data_888 <= (fillup_transition == 1'b1) ? i_input_data[733 % IN_WIDTH] : pong_storage_data_888 ^ i_input_data[733 % IN_WIDTH];
                1010 / IN_WIDTH: pong_storage_data_888 <= (fillup_transition == 1'b1) ? i_input_data[1010 % IN_WIDTH] : pong_storage_data_888 ^ i_input_data[1010 % IN_WIDTH];
                1104 / IN_WIDTH: pong_storage_data_888 <= (fillup_transition == 1'b1) ? i_input_data[1104 % IN_WIDTH] : pong_storage_data_888 ^ i_input_data[1104 % IN_WIDTH];
                default: pong_storage_data_888 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_888;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_888 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_888;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_888 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_888;
            end
        end
    end
end

logic ping_storage_data_889;
logic pong_storage_data_889;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_889 <= 1'b0;
        pong_storage_data_889 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                507 / IN_WIDTH: ping_storage_data_889 <= (fillup_transition == 1'b1) ? i_input_data[507 % IN_WIDTH] : ping_storage_data_889 ^ i_input_data[507 % IN_WIDTH];
                734 / IN_WIDTH: ping_storage_data_889 <= (fillup_transition == 1'b1) ? i_input_data[734 % IN_WIDTH] : ping_storage_data_889 ^ i_input_data[734 % IN_WIDTH];
                1011 / IN_WIDTH: ping_storage_data_889 <= (fillup_transition == 1'b1) ? i_input_data[1011 % IN_WIDTH] : ping_storage_data_889 ^ i_input_data[1011 % IN_WIDTH];
                1105 / IN_WIDTH: ping_storage_data_889 <= (fillup_transition == 1'b1) ? i_input_data[1105 % IN_WIDTH] : ping_storage_data_889 ^ i_input_data[1105 % IN_WIDTH];
                default: ping_storage_data_889 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_889;
                endcase
            end else begin
                case (input_count)
                507 / IN_WIDTH: pong_storage_data_889 <= (fillup_transition == 1'b1) ? i_input_data[507 % IN_WIDTH] : pong_storage_data_889 ^ i_input_data[507 % IN_WIDTH];
                734 / IN_WIDTH: pong_storage_data_889 <= (fillup_transition == 1'b1) ? i_input_data[734 % IN_WIDTH] : pong_storage_data_889 ^ i_input_data[734 % IN_WIDTH];
                1011 / IN_WIDTH: pong_storage_data_889 <= (fillup_transition == 1'b1) ? i_input_data[1011 % IN_WIDTH] : pong_storage_data_889 ^ i_input_data[1011 % IN_WIDTH];
                1105 / IN_WIDTH: pong_storage_data_889 <= (fillup_transition == 1'b1) ? i_input_data[1105 % IN_WIDTH] : pong_storage_data_889 ^ i_input_data[1105 % IN_WIDTH];
                default: pong_storage_data_889 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_889;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_889 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_889;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_889 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_889;
            end
        end
    end
end

logic ping_storage_data_890;
logic pong_storage_data_890;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_890 <= 1'b0;
        pong_storage_data_890 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                508 / IN_WIDTH: ping_storage_data_890 <= (fillup_transition == 1'b1) ? i_input_data[508 % IN_WIDTH] : ping_storage_data_890 ^ i_input_data[508 % IN_WIDTH];
                735 / IN_WIDTH: ping_storage_data_890 <= (fillup_transition == 1'b1) ? i_input_data[735 % IN_WIDTH] : ping_storage_data_890 ^ i_input_data[735 % IN_WIDTH];
                1012 / IN_WIDTH: ping_storage_data_890 <= (fillup_transition == 1'b1) ? i_input_data[1012 % IN_WIDTH] : ping_storage_data_890 ^ i_input_data[1012 % IN_WIDTH];
                1106 / IN_WIDTH: ping_storage_data_890 <= (fillup_transition == 1'b1) ? i_input_data[1106 % IN_WIDTH] : ping_storage_data_890 ^ i_input_data[1106 % IN_WIDTH];
                default: ping_storage_data_890 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_890;
                endcase
            end else begin
                case (input_count)
                508 / IN_WIDTH: pong_storage_data_890 <= (fillup_transition == 1'b1) ? i_input_data[508 % IN_WIDTH] : pong_storage_data_890 ^ i_input_data[508 % IN_WIDTH];
                735 / IN_WIDTH: pong_storage_data_890 <= (fillup_transition == 1'b1) ? i_input_data[735 % IN_WIDTH] : pong_storage_data_890 ^ i_input_data[735 % IN_WIDTH];
                1012 / IN_WIDTH: pong_storage_data_890 <= (fillup_transition == 1'b1) ? i_input_data[1012 % IN_WIDTH] : pong_storage_data_890 ^ i_input_data[1012 % IN_WIDTH];
                1106 / IN_WIDTH: pong_storage_data_890 <= (fillup_transition == 1'b1) ? i_input_data[1106 % IN_WIDTH] : pong_storage_data_890 ^ i_input_data[1106 % IN_WIDTH];
                default: pong_storage_data_890 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_890;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_890 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_890;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_890 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_890;
            end
        end
    end
end

logic ping_storage_data_891;
logic pong_storage_data_891;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_891 <= 1'b0;
        pong_storage_data_891 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                509 / IN_WIDTH: ping_storage_data_891 <= (fillup_transition == 1'b1) ? i_input_data[509 % IN_WIDTH] : ping_storage_data_891 ^ i_input_data[509 % IN_WIDTH];
                736 / IN_WIDTH: ping_storage_data_891 <= (fillup_transition == 1'b1) ? i_input_data[736 % IN_WIDTH] : ping_storage_data_891 ^ i_input_data[736 % IN_WIDTH];
                1013 / IN_WIDTH: ping_storage_data_891 <= (fillup_transition == 1'b1) ? i_input_data[1013 % IN_WIDTH] : ping_storage_data_891 ^ i_input_data[1013 % IN_WIDTH];
                1107 / IN_WIDTH: ping_storage_data_891 <= (fillup_transition == 1'b1) ? i_input_data[1107 % IN_WIDTH] : ping_storage_data_891 ^ i_input_data[1107 % IN_WIDTH];
                default: ping_storage_data_891 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_891;
                endcase
            end else begin
                case (input_count)
                509 / IN_WIDTH: pong_storage_data_891 <= (fillup_transition == 1'b1) ? i_input_data[509 % IN_WIDTH] : pong_storage_data_891 ^ i_input_data[509 % IN_WIDTH];
                736 / IN_WIDTH: pong_storage_data_891 <= (fillup_transition == 1'b1) ? i_input_data[736 % IN_WIDTH] : pong_storage_data_891 ^ i_input_data[736 % IN_WIDTH];
                1013 / IN_WIDTH: pong_storage_data_891 <= (fillup_transition == 1'b1) ? i_input_data[1013 % IN_WIDTH] : pong_storage_data_891 ^ i_input_data[1013 % IN_WIDTH];
                1107 / IN_WIDTH: pong_storage_data_891 <= (fillup_transition == 1'b1) ? i_input_data[1107 % IN_WIDTH] : pong_storage_data_891 ^ i_input_data[1107 % IN_WIDTH];
                default: pong_storage_data_891 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_891;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_891 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_891;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_891 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_891;
            end
        end
    end
end

logic ping_storage_data_892;
logic pong_storage_data_892;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_892 <= 1'b0;
        pong_storage_data_892 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                510 / IN_WIDTH: ping_storage_data_892 <= (fillup_transition == 1'b1) ? i_input_data[510 % IN_WIDTH] : ping_storage_data_892 ^ i_input_data[510 % IN_WIDTH];
                737 / IN_WIDTH: ping_storage_data_892 <= (fillup_transition == 1'b1) ? i_input_data[737 % IN_WIDTH] : ping_storage_data_892 ^ i_input_data[737 % IN_WIDTH];
                1014 / IN_WIDTH: ping_storage_data_892 <= (fillup_transition == 1'b1) ? i_input_data[1014 % IN_WIDTH] : ping_storage_data_892 ^ i_input_data[1014 % IN_WIDTH];
                1108 / IN_WIDTH: ping_storage_data_892 <= (fillup_transition == 1'b1) ? i_input_data[1108 % IN_WIDTH] : ping_storage_data_892 ^ i_input_data[1108 % IN_WIDTH];
                default: ping_storage_data_892 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_892;
                endcase
            end else begin
                case (input_count)
                510 / IN_WIDTH: pong_storage_data_892 <= (fillup_transition == 1'b1) ? i_input_data[510 % IN_WIDTH] : pong_storage_data_892 ^ i_input_data[510 % IN_WIDTH];
                737 / IN_WIDTH: pong_storage_data_892 <= (fillup_transition == 1'b1) ? i_input_data[737 % IN_WIDTH] : pong_storage_data_892 ^ i_input_data[737 % IN_WIDTH];
                1014 / IN_WIDTH: pong_storage_data_892 <= (fillup_transition == 1'b1) ? i_input_data[1014 % IN_WIDTH] : pong_storage_data_892 ^ i_input_data[1014 % IN_WIDTH];
                1108 / IN_WIDTH: pong_storage_data_892 <= (fillup_transition == 1'b1) ? i_input_data[1108 % IN_WIDTH] : pong_storage_data_892 ^ i_input_data[1108 % IN_WIDTH];
                default: pong_storage_data_892 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_892;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_892 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_892;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_892 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_892;
            end
        end
    end
end

logic ping_storage_data_893;
logic pong_storage_data_893;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_893 <= 1'b0;
        pong_storage_data_893 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                511 / IN_WIDTH: ping_storage_data_893 <= (fillup_transition == 1'b1) ? i_input_data[511 % IN_WIDTH] : ping_storage_data_893 ^ i_input_data[511 % IN_WIDTH];
                738 / IN_WIDTH: ping_storage_data_893 <= (fillup_transition == 1'b1) ? i_input_data[738 % IN_WIDTH] : ping_storage_data_893 ^ i_input_data[738 % IN_WIDTH];
                1015 / IN_WIDTH: ping_storage_data_893 <= (fillup_transition == 1'b1) ? i_input_data[1015 % IN_WIDTH] : ping_storage_data_893 ^ i_input_data[1015 % IN_WIDTH];
                1109 / IN_WIDTH: ping_storage_data_893 <= (fillup_transition == 1'b1) ? i_input_data[1109 % IN_WIDTH] : ping_storage_data_893 ^ i_input_data[1109 % IN_WIDTH];
                default: ping_storage_data_893 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_893;
                endcase
            end else begin
                case (input_count)
                511 / IN_WIDTH: pong_storage_data_893 <= (fillup_transition == 1'b1) ? i_input_data[511 % IN_WIDTH] : pong_storage_data_893 ^ i_input_data[511 % IN_WIDTH];
                738 / IN_WIDTH: pong_storage_data_893 <= (fillup_transition == 1'b1) ? i_input_data[738 % IN_WIDTH] : pong_storage_data_893 ^ i_input_data[738 % IN_WIDTH];
                1015 / IN_WIDTH: pong_storage_data_893 <= (fillup_transition == 1'b1) ? i_input_data[1015 % IN_WIDTH] : pong_storage_data_893 ^ i_input_data[1015 % IN_WIDTH];
                1109 / IN_WIDTH: pong_storage_data_893 <= (fillup_transition == 1'b1) ? i_input_data[1109 % IN_WIDTH] : pong_storage_data_893 ^ i_input_data[1109 % IN_WIDTH];
                default: pong_storage_data_893 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_893;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_893 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_893;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_893 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_893;
            end
        end
    end
end

logic ping_storage_data_894;
logic pong_storage_data_894;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_894 <= 1'b0;
        pong_storage_data_894 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                512 / IN_WIDTH: ping_storage_data_894 <= (fillup_transition == 1'b1) ? i_input_data[512 % IN_WIDTH] : ping_storage_data_894 ^ i_input_data[512 % IN_WIDTH];
                739 / IN_WIDTH: ping_storage_data_894 <= (fillup_transition == 1'b1) ? i_input_data[739 % IN_WIDTH] : ping_storage_data_894 ^ i_input_data[739 % IN_WIDTH];
                1016 / IN_WIDTH: ping_storage_data_894 <= (fillup_transition == 1'b1) ? i_input_data[1016 % IN_WIDTH] : ping_storage_data_894 ^ i_input_data[1016 % IN_WIDTH];
                1110 / IN_WIDTH: ping_storage_data_894 <= (fillup_transition == 1'b1) ? i_input_data[1110 % IN_WIDTH] : ping_storage_data_894 ^ i_input_data[1110 % IN_WIDTH];
                default: ping_storage_data_894 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_894;
                endcase
            end else begin
                case (input_count)
                512 / IN_WIDTH: pong_storage_data_894 <= (fillup_transition == 1'b1) ? i_input_data[512 % IN_WIDTH] : pong_storage_data_894 ^ i_input_data[512 % IN_WIDTH];
                739 / IN_WIDTH: pong_storage_data_894 <= (fillup_transition == 1'b1) ? i_input_data[739 % IN_WIDTH] : pong_storage_data_894 ^ i_input_data[739 % IN_WIDTH];
                1016 / IN_WIDTH: pong_storage_data_894 <= (fillup_transition == 1'b1) ? i_input_data[1016 % IN_WIDTH] : pong_storage_data_894 ^ i_input_data[1016 % IN_WIDTH];
                1110 / IN_WIDTH: pong_storage_data_894 <= (fillup_transition == 1'b1) ? i_input_data[1110 % IN_WIDTH] : pong_storage_data_894 ^ i_input_data[1110 % IN_WIDTH];
                default: pong_storage_data_894 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_894;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_894 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_894;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_894 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_894;
            end
        end
    end
end

logic ping_storage_data_895;
logic pong_storage_data_895;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_895 <= 1'b0;
        pong_storage_data_895 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                513 / IN_WIDTH: ping_storage_data_895 <= (fillup_transition == 1'b1) ? i_input_data[513 % IN_WIDTH] : ping_storage_data_895 ^ i_input_data[513 % IN_WIDTH];
                740 / IN_WIDTH: ping_storage_data_895 <= (fillup_transition == 1'b1) ? i_input_data[740 % IN_WIDTH] : ping_storage_data_895 ^ i_input_data[740 % IN_WIDTH];
                1017 / IN_WIDTH: ping_storage_data_895 <= (fillup_transition == 1'b1) ? i_input_data[1017 % IN_WIDTH] : ping_storage_data_895 ^ i_input_data[1017 % IN_WIDTH];
                1111 / IN_WIDTH: ping_storage_data_895 <= (fillup_transition == 1'b1) ? i_input_data[1111 % IN_WIDTH] : ping_storage_data_895 ^ i_input_data[1111 % IN_WIDTH];
                default: ping_storage_data_895 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_895;
                endcase
            end else begin
                case (input_count)
                513 / IN_WIDTH: pong_storage_data_895 <= (fillup_transition == 1'b1) ? i_input_data[513 % IN_WIDTH] : pong_storage_data_895 ^ i_input_data[513 % IN_WIDTH];
                740 / IN_WIDTH: pong_storage_data_895 <= (fillup_transition == 1'b1) ? i_input_data[740 % IN_WIDTH] : pong_storage_data_895 ^ i_input_data[740 % IN_WIDTH];
                1017 / IN_WIDTH: pong_storage_data_895 <= (fillup_transition == 1'b1) ? i_input_data[1017 % IN_WIDTH] : pong_storage_data_895 ^ i_input_data[1017 % IN_WIDTH];
                1111 / IN_WIDTH: pong_storage_data_895 <= (fillup_transition == 1'b1) ? i_input_data[1111 % IN_WIDTH] : pong_storage_data_895 ^ i_input_data[1111 % IN_WIDTH];
                default: pong_storage_data_895 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_895;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_895 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_895;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_895 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_895;
            end
        end
    end
end

logic ping_storage_data_896;
logic pong_storage_data_896;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_896 <= 1'b0;
        pong_storage_data_896 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                514 / IN_WIDTH: ping_storage_data_896 <= (fillup_transition == 1'b1) ? i_input_data[514 % IN_WIDTH] : ping_storage_data_896 ^ i_input_data[514 % IN_WIDTH];
                741 / IN_WIDTH: ping_storage_data_896 <= (fillup_transition == 1'b1) ? i_input_data[741 % IN_WIDTH] : ping_storage_data_896 ^ i_input_data[741 % IN_WIDTH];
                1018 / IN_WIDTH: ping_storage_data_896 <= (fillup_transition == 1'b1) ? i_input_data[1018 % IN_WIDTH] : ping_storage_data_896 ^ i_input_data[1018 % IN_WIDTH];
                1112 / IN_WIDTH: ping_storage_data_896 <= (fillup_transition == 1'b1) ? i_input_data[1112 % IN_WIDTH] : ping_storage_data_896 ^ i_input_data[1112 % IN_WIDTH];
                default: ping_storage_data_896 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_896;
                endcase
            end else begin
                case (input_count)
                514 / IN_WIDTH: pong_storage_data_896 <= (fillup_transition == 1'b1) ? i_input_data[514 % IN_WIDTH] : pong_storage_data_896 ^ i_input_data[514 % IN_WIDTH];
                741 / IN_WIDTH: pong_storage_data_896 <= (fillup_transition == 1'b1) ? i_input_data[741 % IN_WIDTH] : pong_storage_data_896 ^ i_input_data[741 % IN_WIDTH];
                1018 / IN_WIDTH: pong_storage_data_896 <= (fillup_transition == 1'b1) ? i_input_data[1018 % IN_WIDTH] : pong_storage_data_896 ^ i_input_data[1018 % IN_WIDTH];
                1112 / IN_WIDTH: pong_storage_data_896 <= (fillup_transition == 1'b1) ? i_input_data[1112 % IN_WIDTH] : pong_storage_data_896 ^ i_input_data[1112 % IN_WIDTH];
                default: pong_storage_data_896 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_896;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_896 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_896;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_896 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_896;
            end
        end
    end
end

logic ping_storage_data_897;
logic pong_storage_data_897;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_897 <= 1'b0;
        pong_storage_data_897 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                515 / IN_WIDTH: ping_storage_data_897 <= (fillup_transition == 1'b1) ? i_input_data[515 % IN_WIDTH] : ping_storage_data_897 ^ i_input_data[515 % IN_WIDTH];
                742 / IN_WIDTH: ping_storage_data_897 <= (fillup_transition == 1'b1) ? i_input_data[742 % IN_WIDTH] : ping_storage_data_897 ^ i_input_data[742 % IN_WIDTH];
                1019 / IN_WIDTH: ping_storage_data_897 <= (fillup_transition == 1'b1) ? i_input_data[1019 % IN_WIDTH] : ping_storage_data_897 ^ i_input_data[1019 % IN_WIDTH];
                1113 / IN_WIDTH: ping_storage_data_897 <= (fillup_transition == 1'b1) ? i_input_data[1113 % IN_WIDTH] : ping_storage_data_897 ^ i_input_data[1113 % IN_WIDTH];
                default: ping_storage_data_897 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_897;
                endcase
            end else begin
                case (input_count)
                515 / IN_WIDTH: pong_storage_data_897 <= (fillup_transition == 1'b1) ? i_input_data[515 % IN_WIDTH] : pong_storage_data_897 ^ i_input_data[515 % IN_WIDTH];
                742 / IN_WIDTH: pong_storage_data_897 <= (fillup_transition == 1'b1) ? i_input_data[742 % IN_WIDTH] : pong_storage_data_897 ^ i_input_data[742 % IN_WIDTH];
                1019 / IN_WIDTH: pong_storage_data_897 <= (fillup_transition == 1'b1) ? i_input_data[1019 % IN_WIDTH] : pong_storage_data_897 ^ i_input_data[1019 % IN_WIDTH];
                1113 / IN_WIDTH: pong_storage_data_897 <= (fillup_transition == 1'b1) ? i_input_data[1113 % IN_WIDTH] : pong_storage_data_897 ^ i_input_data[1113 % IN_WIDTH];
                default: pong_storage_data_897 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_897;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_897 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_897;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_897 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_897;
            end
        end
    end
end

logic ping_storage_data_898;
logic pong_storage_data_898;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_898 <= 1'b0;
        pong_storage_data_898 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                516 / IN_WIDTH: ping_storage_data_898 <= (fillup_transition == 1'b1) ? i_input_data[516 % IN_WIDTH] : ping_storage_data_898 ^ i_input_data[516 % IN_WIDTH];
                743 / IN_WIDTH: ping_storage_data_898 <= (fillup_transition == 1'b1) ? i_input_data[743 % IN_WIDTH] : ping_storage_data_898 ^ i_input_data[743 % IN_WIDTH];
                1020 / IN_WIDTH: ping_storage_data_898 <= (fillup_transition == 1'b1) ? i_input_data[1020 % IN_WIDTH] : ping_storage_data_898 ^ i_input_data[1020 % IN_WIDTH];
                1114 / IN_WIDTH: ping_storage_data_898 <= (fillup_transition == 1'b1) ? i_input_data[1114 % IN_WIDTH] : ping_storage_data_898 ^ i_input_data[1114 % IN_WIDTH];
                default: ping_storage_data_898 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_898;
                endcase
            end else begin
                case (input_count)
                516 / IN_WIDTH: pong_storage_data_898 <= (fillup_transition == 1'b1) ? i_input_data[516 % IN_WIDTH] : pong_storage_data_898 ^ i_input_data[516 % IN_WIDTH];
                743 / IN_WIDTH: pong_storage_data_898 <= (fillup_transition == 1'b1) ? i_input_data[743 % IN_WIDTH] : pong_storage_data_898 ^ i_input_data[743 % IN_WIDTH];
                1020 / IN_WIDTH: pong_storage_data_898 <= (fillup_transition == 1'b1) ? i_input_data[1020 % IN_WIDTH] : pong_storage_data_898 ^ i_input_data[1020 % IN_WIDTH];
                1114 / IN_WIDTH: pong_storage_data_898 <= (fillup_transition == 1'b1) ? i_input_data[1114 % IN_WIDTH] : pong_storage_data_898 ^ i_input_data[1114 % IN_WIDTH];
                default: pong_storage_data_898 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_898;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_898 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_898;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_898 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_898;
            end
        end
    end
end

logic ping_storage_data_899;
logic pong_storage_data_899;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_899 <= 1'b0;
        pong_storage_data_899 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                517 / IN_WIDTH: ping_storage_data_899 <= (fillup_transition == 1'b1) ? i_input_data[517 % IN_WIDTH] : ping_storage_data_899 ^ i_input_data[517 % IN_WIDTH];
                744 / IN_WIDTH: ping_storage_data_899 <= (fillup_transition == 1'b1) ? i_input_data[744 % IN_WIDTH] : ping_storage_data_899 ^ i_input_data[744 % IN_WIDTH];
                1021 / IN_WIDTH: ping_storage_data_899 <= (fillup_transition == 1'b1) ? i_input_data[1021 % IN_WIDTH] : ping_storage_data_899 ^ i_input_data[1021 % IN_WIDTH];
                1115 / IN_WIDTH: ping_storage_data_899 <= (fillup_transition == 1'b1) ? i_input_data[1115 % IN_WIDTH] : ping_storage_data_899 ^ i_input_data[1115 % IN_WIDTH];
                default: ping_storage_data_899 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_899;
                endcase
            end else begin
                case (input_count)
                517 / IN_WIDTH: pong_storage_data_899 <= (fillup_transition == 1'b1) ? i_input_data[517 % IN_WIDTH] : pong_storage_data_899 ^ i_input_data[517 % IN_WIDTH];
                744 / IN_WIDTH: pong_storage_data_899 <= (fillup_transition == 1'b1) ? i_input_data[744 % IN_WIDTH] : pong_storage_data_899 ^ i_input_data[744 % IN_WIDTH];
                1021 / IN_WIDTH: pong_storage_data_899 <= (fillup_transition == 1'b1) ? i_input_data[1021 % IN_WIDTH] : pong_storage_data_899 ^ i_input_data[1021 % IN_WIDTH];
                1115 / IN_WIDTH: pong_storage_data_899 <= (fillup_transition == 1'b1) ? i_input_data[1115 % IN_WIDTH] : pong_storage_data_899 ^ i_input_data[1115 % IN_WIDTH];
                default: pong_storage_data_899 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_899;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_899 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_899;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_899 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_899;
            end
        end
    end
end

logic ping_storage_data_900;
logic pong_storage_data_900;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_900 <= 1'b0;
        pong_storage_data_900 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                518 / IN_WIDTH: ping_storage_data_900 <= (fillup_transition == 1'b1) ? i_input_data[518 % IN_WIDTH] : ping_storage_data_900 ^ i_input_data[518 % IN_WIDTH];
                745 / IN_WIDTH: ping_storage_data_900 <= (fillup_transition == 1'b1) ? i_input_data[745 % IN_WIDTH] : ping_storage_data_900 ^ i_input_data[745 % IN_WIDTH];
                1022 / IN_WIDTH: ping_storage_data_900 <= (fillup_transition == 1'b1) ? i_input_data[1022 % IN_WIDTH] : ping_storage_data_900 ^ i_input_data[1022 % IN_WIDTH];
                1116 / IN_WIDTH: ping_storage_data_900 <= (fillup_transition == 1'b1) ? i_input_data[1116 % IN_WIDTH] : ping_storage_data_900 ^ i_input_data[1116 % IN_WIDTH];
                default: ping_storage_data_900 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_900;
                endcase
            end else begin
                case (input_count)
                518 / IN_WIDTH: pong_storage_data_900 <= (fillup_transition == 1'b1) ? i_input_data[518 % IN_WIDTH] : pong_storage_data_900 ^ i_input_data[518 % IN_WIDTH];
                745 / IN_WIDTH: pong_storage_data_900 <= (fillup_transition == 1'b1) ? i_input_data[745 % IN_WIDTH] : pong_storage_data_900 ^ i_input_data[745 % IN_WIDTH];
                1022 / IN_WIDTH: pong_storage_data_900 <= (fillup_transition == 1'b1) ? i_input_data[1022 % IN_WIDTH] : pong_storage_data_900 ^ i_input_data[1022 % IN_WIDTH];
                1116 / IN_WIDTH: pong_storage_data_900 <= (fillup_transition == 1'b1) ? i_input_data[1116 % IN_WIDTH] : pong_storage_data_900 ^ i_input_data[1116 % IN_WIDTH];
                default: pong_storage_data_900 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_900;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_900 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_900;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_900 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_900;
            end
        end
    end
end

logic ping_storage_data_901;
logic pong_storage_data_901;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_901 <= 1'b0;
        pong_storage_data_901 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                519 / IN_WIDTH: ping_storage_data_901 <= (fillup_transition == 1'b1) ? i_input_data[519 % IN_WIDTH] : ping_storage_data_901 ^ i_input_data[519 % IN_WIDTH];
                746 / IN_WIDTH: ping_storage_data_901 <= (fillup_transition == 1'b1) ? i_input_data[746 % IN_WIDTH] : ping_storage_data_901 ^ i_input_data[746 % IN_WIDTH];
                1023 / IN_WIDTH: ping_storage_data_901 <= (fillup_transition == 1'b1) ? i_input_data[1023 % IN_WIDTH] : ping_storage_data_901 ^ i_input_data[1023 % IN_WIDTH];
                1117 / IN_WIDTH: ping_storage_data_901 <= (fillup_transition == 1'b1) ? i_input_data[1117 % IN_WIDTH] : ping_storage_data_901 ^ i_input_data[1117 % IN_WIDTH];
                default: ping_storage_data_901 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_901;
                endcase
            end else begin
                case (input_count)
                519 / IN_WIDTH: pong_storage_data_901 <= (fillup_transition == 1'b1) ? i_input_data[519 % IN_WIDTH] : pong_storage_data_901 ^ i_input_data[519 % IN_WIDTH];
                746 / IN_WIDTH: pong_storage_data_901 <= (fillup_transition == 1'b1) ? i_input_data[746 % IN_WIDTH] : pong_storage_data_901 ^ i_input_data[746 % IN_WIDTH];
                1023 / IN_WIDTH: pong_storage_data_901 <= (fillup_transition == 1'b1) ? i_input_data[1023 % IN_WIDTH] : pong_storage_data_901 ^ i_input_data[1023 % IN_WIDTH];
                1117 / IN_WIDTH: pong_storage_data_901 <= (fillup_transition == 1'b1) ? i_input_data[1117 % IN_WIDTH] : pong_storage_data_901 ^ i_input_data[1117 % IN_WIDTH];
                default: pong_storage_data_901 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_901;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_901 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_901;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_901 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_901;
            end
        end
    end
end

logic ping_storage_data_902;
logic pong_storage_data_902;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_902 <= 1'b0;
        pong_storage_data_902 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                520 / IN_WIDTH: ping_storage_data_902 <= (fillup_transition == 1'b1) ? i_input_data[520 % IN_WIDTH] : ping_storage_data_902 ^ i_input_data[520 % IN_WIDTH];
                747 / IN_WIDTH: ping_storage_data_902 <= (fillup_transition == 1'b1) ? i_input_data[747 % IN_WIDTH] : ping_storage_data_902 ^ i_input_data[747 % IN_WIDTH];
                1024 / IN_WIDTH: ping_storage_data_902 <= (fillup_transition == 1'b1) ? i_input_data[1024 % IN_WIDTH] : ping_storage_data_902 ^ i_input_data[1024 % IN_WIDTH];
                1118 / IN_WIDTH: ping_storage_data_902 <= (fillup_transition == 1'b1) ? i_input_data[1118 % IN_WIDTH] : ping_storage_data_902 ^ i_input_data[1118 % IN_WIDTH];
                default: ping_storage_data_902 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_902;
                endcase
            end else begin
                case (input_count)
                520 / IN_WIDTH: pong_storage_data_902 <= (fillup_transition == 1'b1) ? i_input_data[520 % IN_WIDTH] : pong_storage_data_902 ^ i_input_data[520 % IN_WIDTH];
                747 / IN_WIDTH: pong_storage_data_902 <= (fillup_transition == 1'b1) ? i_input_data[747 % IN_WIDTH] : pong_storage_data_902 ^ i_input_data[747 % IN_WIDTH];
                1024 / IN_WIDTH: pong_storage_data_902 <= (fillup_transition == 1'b1) ? i_input_data[1024 % IN_WIDTH] : pong_storage_data_902 ^ i_input_data[1024 % IN_WIDTH];
                1118 / IN_WIDTH: pong_storage_data_902 <= (fillup_transition == 1'b1) ? i_input_data[1118 % IN_WIDTH] : pong_storage_data_902 ^ i_input_data[1118 % IN_WIDTH];
                default: pong_storage_data_902 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_902;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_902 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_902;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_902 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_902;
            end
        end
    end
end

logic ping_storage_data_903;
logic pong_storage_data_903;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_903 <= 1'b0;
        pong_storage_data_903 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                521 / IN_WIDTH: ping_storage_data_903 <= (fillup_transition == 1'b1) ? i_input_data[521 % IN_WIDTH] : ping_storage_data_903 ^ i_input_data[521 % IN_WIDTH];
                748 / IN_WIDTH: ping_storage_data_903 <= (fillup_transition == 1'b1) ? i_input_data[748 % IN_WIDTH] : ping_storage_data_903 ^ i_input_data[748 % IN_WIDTH];
                1025 / IN_WIDTH: ping_storage_data_903 <= (fillup_transition == 1'b1) ? i_input_data[1025 % IN_WIDTH] : ping_storage_data_903 ^ i_input_data[1025 % IN_WIDTH];
                1119 / IN_WIDTH: ping_storage_data_903 <= (fillup_transition == 1'b1) ? i_input_data[1119 % IN_WIDTH] : ping_storage_data_903 ^ i_input_data[1119 % IN_WIDTH];
                default: ping_storage_data_903 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_903;
                endcase
            end else begin
                case (input_count)
                521 / IN_WIDTH: pong_storage_data_903 <= (fillup_transition == 1'b1) ? i_input_data[521 % IN_WIDTH] : pong_storage_data_903 ^ i_input_data[521 % IN_WIDTH];
                748 / IN_WIDTH: pong_storage_data_903 <= (fillup_transition == 1'b1) ? i_input_data[748 % IN_WIDTH] : pong_storage_data_903 ^ i_input_data[748 % IN_WIDTH];
                1025 / IN_WIDTH: pong_storage_data_903 <= (fillup_transition == 1'b1) ? i_input_data[1025 % IN_WIDTH] : pong_storage_data_903 ^ i_input_data[1025 % IN_WIDTH];
                1119 / IN_WIDTH: pong_storage_data_903 <= (fillup_transition == 1'b1) ? i_input_data[1119 % IN_WIDTH] : pong_storage_data_903 ^ i_input_data[1119 % IN_WIDTH];
                default: pong_storage_data_903 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_903;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_903 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_903;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_903 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_903;
            end
        end
    end
end

logic ping_storage_data_904;
logic pong_storage_data_904;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_904 <= 1'b0;
        pong_storage_data_904 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                522 / IN_WIDTH: ping_storage_data_904 <= (fillup_transition == 1'b1) ? i_input_data[522 % IN_WIDTH] : ping_storage_data_904 ^ i_input_data[522 % IN_WIDTH];
                749 / IN_WIDTH: ping_storage_data_904 <= (fillup_transition == 1'b1) ? i_input_data[749 % IN_WIDTH] : ping_storage_data_904 ^ i_input_data[749 % IN_WIDTH];
                1026 / IN_WIDTH: ping_storage_data_904 <= (fillup_transition == 1'b1) ? i_input_data[1026 % IN_WIDTH] : ping_storage_data_904 ^ i_input_data[1026 % IN_WIDTH];
                1120 / IN_WIDTH: ping_storage_data_904 <= (fillup_transition == 1'b1) ? i_input_data[1120 % IN_WIDTH] : ping_storage_data_904 ^ i_input_data[1120 % IN_WIDTH];
                default: ping_storage_data_904 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_904;
                endcase
            end else begin
                case (input_count)
                522 / IN_WIDTH: pong_storage_data_904 <= (fillup_transition == 1'b1) ? i_input_data[522 % IN_WIDTH] : pong_storage_data_904 ^ i_input_data[522 % IN_WIDTH];
                749 / IN_WIDTH: pong_storage_data_904 <= (fillup_transition == 1'b1) ? i_input_data[749 % IN_WIDTH] : pong_storage_data_904 ^ i_input_data[749 % IN_WIDTH];
                1026 / IN_WIDTH: pong_storage_data_904 <= (fillup_transition == 1'b1) ? i_input_data[1026 % IN_WIDTH] : pong_storage_data_904 ^ i_input_data[1026 % IN_WIDTH];
                1120 / IN_WIDTH: pong_storage_data_904 <= (fillup_transition == 1'b1) ? i_input_data[1120 % IN_WIDTH] : pong_storage_data_904 ^ i_input_data[1120 % IN_WIDTH];
                default: pong_storage_data_904 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_904;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_904 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_904;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_904 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_904;
            end
        end
    end
end

logic ping_storage_data_905;
logic pong_storage_data_905;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_905 <= 1'b0;
        pong_storage_data_905 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                523 / IN_WIDTH: ping_storage_data_905 <= (fillup_transition == 1'b1) ? i_input_data[523 % IN_WIDTH] : ping_storage_data_905 ^ i_input_data[523 % IN_WIDTH];
                750 / IN_WIDTH: ping_storage_data_905 <= (fillup_transition == 1'b1) ? i_input_data[750 % IN_WIDTH] : ping_storage_data_905 ^ i_input_data[750 % IN_WIDTH];
                1027 / IN_WIDTH: ping_storage_data_905 <= (fillup_transition == 1'b1) ? i_input_data[1027 % IN_WIDTH] : ping_storage_data_905 ^ i_input_data[1027 % IN_WIDTH];
                1121 / IN_WIDTH: ping_storage_data_905 <= (fillup_transition == 1'b1) ? i_input_data[1121 % IN_WIDTH] : ping_storage_data_905 ^ i_input_data[1121 % IN_WIDTH];
                default: ping_storage_data_905 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_905;
                endcase
            end else begin
                case (input_count)
                523 / IN_WIDTH: pong_storage_data_905 <= (fillup_transition == 1'b1) ? i_input_data[523 % IN_WIDTH] : pong_storage_data_905 ^ i_input_data[523 % IN_WIDTH];
                750 / IN_WIDTH: pong_storage_data_905 <= (fillup_transition == 1'b1) ? i_input_data[750 % IN_WIDTH] : pong_storage_data_905 ^ i_input_data[750 % IN_WIDTH];
                1027 / IN_WIDTH: pong_storage_data_905 <= (fillup_transition == 1'b1) ? i_input_data[1027 % IN_WIDTH] : pong_storage_data_905 ^ i_input_data[1027 % IN_WIDTH];
                1121 / IN_WIDTH: pong_storage_data_905 <= (fillup_transition == 1'b1) ? i_input_data[1121 % IN_WIDTH] : pong_storage_data_905 ^ i_input_data[1121 % IN_WIDTH];
                default: pong_storage_data_905 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_905;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_905 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_905;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_905 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_905;
            end
        end
    end
end

logic ping_storage_data_906;
logic pong_storage_data_906;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_906 <= 1'b0;
        pong_storage_data_906 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                524 / IN_WIDTH: ping_storage_data_906 <= (fillup_transition == 1'b1) ? i_input_data[524 % IN_WIDTH] : ping_storage_data_906 ^ i_input_data[524 % IN_WIDTH];
                751 / IN_WIDTH: ping_storage_data_906 <= (fillup_transition == 1'b1) ? i_input_data[751 % IN_WIDTH] : ping_storage_data_906 ^ i_input_data[751 % IN_WIDTH];
                1028 / IN_WIDTH: ping_storage_data_906 <= (fillup_transition == 1'b1) ? i_input_data[1028 % IN_WIDTH] : ping_storage_data_906 ^ i_input_data[1028 % IN_WIDTH];
                1122 / IN_WIDTH: ping_storage_data_906 <= (fillup_transition == 1'b1) ? i_input_data[1122 % IN_WIDTH] : ping_storage_data_906 ^ i_input_data[1122 % IN_WIDTH];
                default: ping_storage_data_906 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_906;
                endcase
            end else begin
                case (input_count)
                524 / IN_WIDTH: pong_storage_data_906 <= (fillup_transition == 1'b1) ? i_input_data[524 % IN_WIDTH] : pong_storage_data_906 ^ i_input_data[524 % IN_WIDTH];
                751 / IN_WIDTH: pong_storage_data_906 <= (fillup_transition == 1'b1) ? i_input_data[751 % IN_WIDTH] : pong_storage_data_906 ^ i_input_data[751 % IN_WIDTH];
                1028 / IN_WIDTH: pong_storage_data_906 <= (fillup_transition == 1'b1) ? i_input_data[1028 % IN_WIDTH] : pong_storage_data_906 ^ i_input_data[1028 % IN_WIDTH];
                1122 / IN_WIDTH: pong_storage_data_906 <= (fillup_transition == 1'b1) ? i_input_data[1122 % IN_WIDTH] : pong_storage_data_906 ^ i_input_data[1122 % IN_WIDTH];
                default: pong_storage_data_906 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_906;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_906 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_906;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_906 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_906;
            end
        end
    end
end

logic ping_storage_data_907;
logic pong_storage_data_907;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_907 <= 1'b0;
        pong_storage_data_907 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                525 / IN_WIDTH: ping_storage_data_907 <= (fillup_transition == 1'b1) ? i_input_data[525 % IN_WIDTH] : ping_storage_data_907 ^ i_input_data[525 % IN_WIDTH];
                752 / IN_WIDTH: ping_storage_data_907 <= (fillup_transition == 1'b1) ? i_input_data[752 % IN_WIDTH] : ping_storage_data_907 ^ i_input_data[752 % IN_WIDTH];
                1029 / IN_WIDTH: ping_storage_data_907 <= (fillup_transition == 1'b1) ? i_input_data[1029 % IN_WIDTH] : ping_storage_data_907 ^ i_input_data[1029 % IN_WIDTH];
                1123 / IN_WIDTH: ping_storage_data_907 <= (fillup_transition == 1'b1) ? i_input_data[1123 % IN_WIDTH] : ping_storage_data_907 ^ i_input_data[1123 % IN_WIDTH];
                default: ping_storage_data_907 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_907;
                endcase
            end else begin
                case (input_count)
                525 / IN_WIDTH: pong_storage_data_907 <= (fillup_transition == 1'b1) ? i_input_data[525 % IN_WIDTH] : pong_storage_data_907 ^ i_input_data[525 % IN_WIDTH];
                752 / IN_WIDTH: pong_storage_data_907 <= (fillup_transition == 1'b1) ? i_input_data[752 % IN_WIDTH] : pong_storage_data_907 ^ i_input_data[752 % IN_WIDTH];
                1029 / IN_WIDTH: pong_storage_data_907 <= (fillup_transition == 1'b1) ? i_input_data[1029 % IN_WIDTH] : pong_storage_data_907 ^ i_input_data[1029 % IN_WIDTH];
                1123 / IN_WIDTH: pong_storage_data_907 <= (fillup_transition == 1'b1) ? i_input_data[1123 % IN_WIDTH] : pong_storage_data_907 ^ i_input_data[1123 % IN_WIDTH];
                default: pong_storage_data_907 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_907;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_907 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_907;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_907 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_907;
            end
        end
    end
end

logic ping_storage_data_908;
logic pong_storage_data_908;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_908 <= 1'b0;
        pong_storage_data_908 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                526 / IN_WIDTH: ping_storage_data_908 <= (fillup_transition == 1'b1) ? i_input_data[526 % IN_WIDTH] : ping_storage_data_908 ^ i_input_data[526 % IN_WIDTH];
                753 / IN_WIDTH: ping_storage_data_908 <= (fillup_transition == 1'b1) ? i_input_data[753 % IN_WIDTH] : ping_storage_data_908 ^ i_input_data[753 % IN_WIDTH];
                1030 / IN_WIDTH: ping_storage_data_908 <= (fillup_transition == 1'b1) ? i_input_data[1030 % IN_WIDTH] : ping_storage_data_908 ^ i_input_data[1030 % IN_WIDTH];
                1124 / IN_WIDTH: ping_storage_data_908 <= (fillup_transition == 1'b1) ? i_input_data[1124 % IN_WIDTH] : ping_storage_data_908 ^ i_input_data[1124 % IN_WIDTH];
                default: ping_storage_data_908 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_908;
                endcase
            end else begin
                case (input_count)
                526 / IN_WIDTH: pong_storage_data_908 <= (fillup_transition == 1'b1) ? i_input_data[526 % IN_WIDTH] : pong_storage_data_908 ^ i_input_data[526 % IN_WIDTH];
                753 / IN_WIDTH: pong_storage_data_908 <= (fillup_transition == 1'b1) ? i_input_data[753 % IN_WIDTH] : pong_storage_data_908 ^ i_input_data[753 % IN_WIDTH];
                1030 / IN_WIDTH: pong_storage_data_908 <= (fillup_transition == 1'b1) ? i_input_data[1030 % IN_WIDTH] : pong_storage_data_908 ^ i_input_data[1030 % IN_WIDTH];
                1124 / IN_WIDTH: pong_storage_data_908 <= (fillup_transition == 1'b1) ? i_input_data[1124 % IN_WIDTH] : pong_storage_data_908 ^ i_input_data[1124 % IN_WIDTH];
                default: pong_storage_data_908 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_908;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_908 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_908;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_908 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_908;
            end
        end
    end
end

logic ping_storage_data_909;
logic pong_storage_data_909;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_909 <= 1'b0;
        pong_storage_data_909 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                527 / IN_WIDTH: ping_storage_data_909 <= (fillup_transition == 1'b1) ? i_input_data[527 % IN_WIDTH] : ping_storage_data_909 ^ i_input_data[527 % IN_WIDTH];
                754 / IN_WIDTH: ping_storage_data_909 <= (fillup_transition == 1'b1) ? i_input_data[754 % IN_WIDTH] : ping_storage_data_909 ^ i_input_data[754 % IN_WIDTH];
                1031 / IN_WIDTH: ping_storage_data_909 <= (fillup_transition == 1'b1) ? i_input_data[1031 % IN_WIDTH] : ping_storage_data_909 ^ i_input_data[1031 % IN_WIDTH];
                1125 / IN_WIDTH: ping_storage_data_909 <= (fillup_transition == 1'b1) ? i_input_data[1125 % IN_WIDTH] : ping_storage_data_909 ^ i_input_data[1125 % IN_WIDTH];
                default: ping_storage_data_909 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_909;
                endcase
            end else begin
                case (input_count)
                527 / IN_WIDTH: pong_storage_data_909 <= (fillup_transition == 1'b1) ? i_input_data[527 % IN_WIDTH] : pong_storage_data_909 ^ i_input_data[527 % IN_WIDTH];
                754 / IN_WIDTH: pong_storage_data_909 <= (fillup_transition == 1'b1) ? i_input_data[754 % IN_WIDTH] : pong_storage_data_909 ^ i_input_data[754 % IN_WIDTH];
                1031 / IN_WIDTH: pong_storage_data_909 <= (fillup_transition == 1'b1) ? i_input_data[1031 % IN_WIDTH] : pong_storage_data_909 ^ i_input_data[1031 % IN_WIDTH];
                1125 / IN_WIDTH: pong_storage_data_909 <= (fillup_transition == 1'b1) ? i_input_data[1125 % IN_WIDTH] : pong_storage_data_909 ^ i_input_data[1125 % IN_WIDTH];
                default: pong_storage_data_909 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_909;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_909 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_909;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_909 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_909;
            end
        end
    end
end

logic ping_storage_data_910;
logic pong_storage_data_910;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_910 <= 1'b0;
        pong_storage_data_910 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                528 / IN_WIDTH: ping_storage_data_910 <= (fillup_transition == 1'b1) ? i_input_data[528 % IN_WIDTH] : ping_storage_data_910 ^ i_input_data[528 % IN_WIDTH];
                755 / IN_WIDTH: ping_storage_data_910 <= (fillup_transition == 1'b1) ? i_input_data[755 % IN_WIDTH] : ping_storage_data_910 ^ i_input_data[755 % IN_WIDTH];
                1032 / IN_WIDTH: ping_storage_data_910 <= (fillup_transition == 1'b1) ? i_input_data[1032 % IN_WIDTH] : ping_storage_data_910 ^ i_input_data[1032 % IN_WIDTH];
                1126 / IN_WIDTH: ping_storage_data_910 <= (fillup_transition == 1'b1) ? i_input_data[1126 % IN_WIDTH] : ping_storage_data_910 ^ i_input_data[1126 % IN_WIDTH];
                default: ping_storage_data_910 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_910;
                endcase
            end else begin
                case (input_count)
                528 / IN_WIDTH: pong_storage_data_910 <= (fillup_transition == 1'b1) ? i_input_data[528 % IN_WIDTH] : pong_storage_data_910 ^ i_input_data[528 % IN_WIDTH];
                755 / IN_WIDTH: pong_storage_data_910 <= (fillup_transition == 1'b1) ? i_input_data[755 % IN_WIDTH] : pong_storage_data_910 ^ i_input_data[755 % IN_WIDTH];
                1032 / IN_WIDTH: pong_storage_data_910 <= (fillup_transition == 1'b1) ? i_input_data[1032 % IN_WIDTH] : pong_storage_data_910 ^ i_input_data[1032 % IN_WIDTH];
                1126 / IN_WIDTH: pong_storage_data_910 <= (fillup_transition == 1'b1) ? i_input_data[1126 % IN_WIDTH] : pong_storage_data_910 ^ i_input_data[1126 % IN_WIDTH];
                default: pong_storage_data_910 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_910;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_910 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_910;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_910 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_910;
            end
        end
    end
end

logic ping_storage_data_911;
logic pong_storage_data_911;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_911 <= 1'b0;
        pong_storage_data_911 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                529 / IN_WIDTH: ping_storage_data_911 <= (fillup_transition == 1'b1) ? i_input_data[529 % IN_WIDTH] : ping_storage_data_911 ^ i_input_data[529 % IN_WIDTH];
                756 / IN_WIDTH: ping_storage_data_911 <= (fillup_transition == 1'b1) ? i_input_data[756 % IN_WIDTH] : ping_storage_data_911 ^ i_input_data[756 % IN_WIDTH];
                1033 / IN_WIDTH: ping_storage_data_911 <= (fillup_transition == 1'b1) ? i_input_data[1033 % IN_WIDTH] : ping_storage_data_911 ^ i_input_data[1033 % IN_WIDTH];
                1127 / IN_WIDTH: ping_storage_data_911 <= (fillup_transition == 1'b1) ? i_input_data[1127 % IN_WIDTH] : ping_storage_data_911 ^ i_input_data[1127 % IN_WIDTH];
                default: ping_storage_data_911 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_911;
                endcase
            end else begin
                case (input_count)
                529 / IN_WIDTH: pong_storage_data_911 <= (fillup_transition == 1'b1) ? i_input_data[529 % IN_WIDTH] : pong_storage_data_911 ^ i_input_data[529 % IN_WIDTH];
                756 / IN_WIDTH: pong_storage_data_911 <= (fillup_transition == 1'b1) ? i_input_data[756 % IN_WIDTH] : pong_storage_data_911 ^ i_input_data[756 % IN_WIDTH];
                1033 / IN_WIDTH: pong_storage_data_911 <= (fillup_transition == 1'b1) ? i_input_data[1033 % IN_WIDTH] : pong_storage_data_911 ^ i_input_data[1033 % IN_WIDTH];
                1127 / IN_WIDTH: pong_storage_data_911 <= (fillup_transition == 1'b1) ? i_input_data[1127 % IN_WIDTH] : pong_storage_data_911 ^ i_input_data[1127 % IN_WIDTH];
                default: pong_storage_data_911 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_911;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_911 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_911;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_911 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_911;
            end
        end
    end
end

logic ping_storage_data_912;
logic pong_storage_data_912;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_912 <= 1'b0;
        pong_storage_data_912 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                530 / IN_WIDTH: ping_storage_data_912 <= (fillup_transition == 1'b1) ? i_input_data[530 % IN_WIDTH] : ping_storage_data_912 ^ i_input_data[530 % IN_WIDTH];
                757 / IN_WIDTH: ping_storage_data_912 <= (fillup_transition == 1'b1) ? i_input_data[757 % IN_WIDTH] : ping_storage_data_912 ^ i_input_data[757 % IN_WIDTH];
                1034 / IN_WIDTH: ping_storage_data_912 <= (fillup_transition == 1'b1) ? i_input_data[1034 % IN_WIDTH] : ping_storage_data_912 ^ i_input_data[1034 % IN_WIDTH];
                1128 / IN_WIDTH: ping_storage_data_912 <= (fillup_transition == 1'b1) ? i_input_data[1128 % IN_WIDTH] : ping_storage_data_912 ^ i_input_data[1128 % IN_WIDTH];
                default: ping_storage_data_912 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_912;
                endcase
            end else begin
                case (input_count)
                530 / IN_WIDTH: pong_storage_data_912 <= (fillup_transition == 1'b1) ? i_input_data[530 % IN_WIDTH] : pong_storage_data_912 ^ i_input_data[530 % IN_WIDTH];
                757 / IN_WIDTH: pong_storage_data_912 <= (fillup_transition == 1'b1) ? i_input_data[757 % IN_WIDTH] : pong_storage_data_912 ^ i_input_data[757 % IN_WIDTH];
                1034 / IN_WIDTH: pong_storage_data_912 <= (fillup_transition == 1'b1) ? i_input_data[1034 % IN_WIDTH] : pong_storage_data_912 ^ i_input_data[1034 % IN_WIDTH];
                1128 / IN_WIDTH: pong_storage_data_912 <= (fillup_transition == 1'b1) ? i_input_data[1128 % IN_WIDTH] : pong_storage_data_912 ^ i_input_data[1128 % IN_WIDTH];
                default: pong_storage_data_912 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_912;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_912 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_912;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_912 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_912;
            end
        end
    end
end

logic ping_storage_data_913;
logic pong_storage_data_913;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_913 <= 1'b0;
        pong_storage_data_913 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                531 / IN_WIDTH: ping_storage_data_913 <= (fillup_transition == 1'b1) ? i_input_data[531 % IN_WIDTH] : ping_storage_data_913 ^ i_input_data[531 % IN_WIDTH];
                758 / IN_WIDTH: ping_storage_data_913 <= (fillup_transition == 1'b1) ? i_input_data[758 % IN_WIDTH] : ping_storage_data_913 ^ i_input_data[758 % IN_WIDTH];
                1035 / IN_WIDTH: ping_storage_data_913 <= (fillup_transition == 1'b1) ? i_input_data[1035 % IN_WIDTH] : ping_storage_data_913 ^ i_input_data[1035 % IN_WIDTH];
                1129 / IN_WIDTH: ping_storage_data_913 <= (fillup_transition == 1'b1) ? i_input_data[1129 % IN_WIDTH] : ping_storage_data_913 ^ i_input_data[1129 % IN_WIDTH];
                default: ping_storage_data_913 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_913;
                endcase
            end else begin
                case (input_count)
                531 / IN_WIDTH: pong_storage_data_913 <= (fillup_transition == 1'b1) ? i_input_data[531 % IN_WIDTH] : pong_storage_data_913 ^ i_input_data[531 % IN_WIDTH];
                758 / IN_WIDTH: pong_storage_data_913 <= (fillup_transition == 1'b1) ? i_input_data[758 % IN_WIDTH] : pong_storage_data_913 ^ i_input_data[758 % IN_WIDTH];
                1035 / IN_WIDTH: pong_storage_data_913 <= (fillup_transition == 1'b1) ? i_input_data[1035 % IN_WIDTH] : pong_storage_data_913 ^ i_input_data[1035 % IN_WIDTH];
                1129 / IN_WIDTH: pong_storage_data_913 <= (fillup_transition == 1'b1) ? i_input_data[1129 % IN_WIDTH] : pong_storage_data_913 ^ i_input_data[1129 % IN_WIDTH];
                default: pong_storage_data_913 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_913;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_913 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_913;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_913 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_913;
            end
        end
    end
end

logic ping_storage_data_914;
logic pong_storage_data_914;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_914 <= 1'b0;
        pong_storage_data_914 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                532 / IN_WIDTH: ping_storage_data_914 <= (fillup_transition == 1'b1) ? i_input_data[532 % IN_WIDTH] : ping_storage_data_914 ^ i_input_data[532 % IN_WIDTH];
                759 / IN_WIDTH: ping_storage_data_914 <= (fillup_transition == 1'b1) ? i_input_data[759 % IN_WIDTH] : ping_storage_data_914 ^ i_input_data[759 % IN_WIDTH];
                1036 / IN_WIDTH: ping_storage_data_914 <= (fillup_transition == 1'b1) ? i_input_data[1036 % IN_WIDTH] : ping_storage_data_914 ^ i_input_data[1036 % IN_WIDTH];
                1130 / IN_WIDTH: ping_storage_data_914 <= (fillup_transition == 1'b1) ? i_input_data[1130 % IN_WIDTH] : ping_storage_data_914 ^ i_input_data[1130 % IN_WIDTH];
                default: ping_storage_data_914 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_914;
                endcase
            end else begin
                case (input_count)
                532 / IN_WIDTH: pong_storage_data_914 <= (fillup_transition == 1'b1) ? i_input_data[532 % IN_WIDTH] : pong_storage_data_914 ^ i_input_data[532 % IN_WIDTH];
                759 / IN_WIDTH: pong_storage_data_914 <= (fillup_transition == 1'b1) ? i_input_data[759 % IN_WIDTH] : pong_storage_data_914 ^ i_input_data[759 % IN_WIDTH];
                1036 / IN_WIDTH: pong_storage_data_914 <= (fillup_transition == 1'b1) ? i_input_data[1036 % IN_WIDTH] : pong_storage_data_914 ^ i_input_data[1036 % IN_WIDTH];
                1130 / IN_WIDTH: pong_storage_data_914 <= (fillup_transition == 1'b1) ? i_input_data[1130 % IN_WIDTH] : pong_storage_data_914 ^ i_input_data[1130 % IN_WIDTH];
                default: pong_storage_data_914 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_914;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_914 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_914;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_914 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_914;
            end
        end
    end
end

logic ping_storage_data_915;
logic pong_storage_data_915;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_915 <= 1'b0;
        pong_storage_data_915 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                533 / IN_WIDTH: ping_storage_data_915 <= (fillup_transition == 1'b1) ? i_input_data[533 % IN_WIDTH] : ping_storage_data_915 ^ i_input_data[533 % IN_WIDTH];
                760 / IN_WIDTH: ping_storage_data_915 <= (fillup_transition == 1'b1) ? i_input_data[760 % IN_WIDTH] : ping_storage_data_915 ^ i_input_data[760 % IN_WIDTH];
                1037 / IN_WIDTH: ping_storage_data_915 <= (fillup_transition == 1'b1) ? i_input_data[1037 % IN_WIDTH] : ping_storage_data_915 ^ i_input_data[1037 % IN_WIDTH];
                1131 / IN_WIDTH: ping_storage_data_915 <= (fillup_transition == 1'b1) ? i_input_data[1131 % IN_WIDTH] : ping_storage_data_915 ^ i_input_data[1131 % IN_WIDTH];
                default: ping_storage_data_915 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_915;
                endcase
            end else begin
                case (input_count)
                533 / IN_WIDTH: pong_storage_data_915 <= (fillup_transition == 1'b1) ? i_input_data[533 % IN_WIDTH] : pong_storage_data_915 ^ i_input_data[533 % IN_WIDTH];
                760 / IN_WIDTH: pong_storage_data_915 <= (fillup_transition == 1'b1) ? i_input_data[760 % IN_WIDTH] : pong_storage_data_915 ^ i_input_data[760 % IN_WIDTH];
                1037 / IN_WIDTH: pong_storage_data_915 <= (fillup_transition == 1'b1) ? i_input_data[1037 % IN_WIDTH] : pong_storage_data_915 ^ i_input_data[1037 % IN_WIDTH];
                1131 / IN_WIDTH: pong_storage_data_915 <= (fillup_transition == 1'b1) ? i_input_data[1131 % IN_WIDTH] : pong_storage_data_915 ^ i_input_data[1131 % IN_WIDTH];
                default: pong_storage_data_915 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_915;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_915 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_915;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_915 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_915;
            end
        end
    end
end

logic ping_storage_data_916;
logic pong_storage_data_916;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_916 <= 1'b0;
        pong_storage_data_916 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                534 / IN_WIDTH: ping_storage_data_916 <= (fillup_transition == 1'b1) ? i_input_data[534 % IN_WIDTH] : ping_storage_data_916 ^ i_input_data[534 % IN_WIDTH];
                761 / IN_WIDTH: ping_storage_data_916 <= (fillup_transition == 1'b1) ? i_input_data[761 % IN_WIDTH] : ping_storage_data_916 ^ i_input_data[761 % IN_WIDTH];
                1038 / IN_WIDTH: ping_storage_data_916 <= (fillup_transition == 1'b1) ? i_input_data[1038 % IN_WIDTH] : ping_storage_data_916 ^ i_input_data[1038 % IN_WIDTH];
                1132 / IN_WIDTH: ping_storage_data_916 <= (fillup_transition == 1'b1) ? i_input_data[1132 % IN_WIDTH] : ping_storage_data_916 ^ i_input_data[1132 % IN_WIDTH];
                default: ping_storage_data_916 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_916;
                endcase
            end else begin
                case (input_count)
                534 / IN_WIDTH: pong_storage_data_916 <= (fillup_transition == 1'b1) ? i_input_data[534 % IN_WIDTH] : pong_storage_data_916 ^ i_input_data[534 % IN_WIDTH];
                761 / IN_WIDTH: pong_storage_data_916 <= (fillup_transition == 1'b1) ? i_input_data[761 % IN_WIDTH] : pong_storage_data_916 ^ i_input_data[761 % IN_WIDTH];
                1038 / IN_WIDTH: pong_storage_data_916 <= (fillup_transition == 1'b1) ? i_input_data[1038 % IN_WIDTH] : pong_storage_data_916 ^ i_input_data[1038 % IN_WIDTH];
                1132 / IN_WIDTH: pong_storage_data_916 <= (fillup_transition == 1'b1) ? i_input_data[1132 % IN_WIDTH] : pong_storage_data_916 ^ i_input_data[1132 % IN_WIDTH];
                default: pong_storage_data_916 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_916;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_916 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_916;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_916 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_916;
            end
        end
    end
end

logic ping_storage_data_917;
logic pong_storage_data_917;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_917 <= 1'b0;
        pong_storage_data_917 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                535 / IN_WIDTH: ping_storage_data_917 <= (fillup_transition == 1'b1) ? i_input_data[535 % IN_WIDTH] : ping_storage_data_917 ^ i_input_data[535 % IN_WIDTH];
                762 / IN_WIDTH: ping_storage_data_917 <= (fillup_transition == 1'b1) ? i_input_data[762 % IN_WIDTH] : ping_storage_data_917 ^ i_input_data[762 % IN_WIDTH];
                1039 / IN_WIDTH: ping_storage_data_917 <= (fillup_transition == 1'b1) ? i_input_data[1039 % IN_WIDTH] : ping_storage_data_917 ^ i_input_data[1039 % IN_WIDTH];
                1133 / IN_WIDTH: ping_storage_data_917 <= (fillup_transition == 1'b1) ? i_input_data[1133 % IN_WIDTH] : ping_storage_data_917 ^ i_input_data[1133 % IN_WIDTH];
                default: ping_storage_data_917 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_917;
                endcase
            end else begin
                case (input_count)
                535 / IN_WIDTH: pong_storage_data_917 <= (fillup_transition == 1'b1) ? i_input_data[535 % IN_WIDTH] : pong_storage_data_917 ^ i_input_data[535 % IN_WIDTH];
                762 / IN_WIDTH: pong_storage_data_917 <= (fillup_transition == 1'b1) ? i_input_data[762 % IN_WIDTH] : pong_storage_data_917 ^ i_input_data[762 % IN_WIDTH];
                1039 / IN_WIDTH: pong_storage_data_917 <= (fillup_transition == 1'b1) ? i_input_data[1039 % IN_WIDTH] : pong_storage_data_917 ^ i_input_data[1039 % IN_WIDTH];
                1133 / IN_WIDTH: pong_storage_data_917 <= (fillup_transition == 1'b1) ? i_input_data[1133 % IN_WIDTH] : pong_storage_data_917 ^ i_input_data[1133 % IN_WIDTH];
                default: pong_storage_data_917 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_917;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_917 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_917;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_917 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_917;
            end
        end
    end
end

logic ping_storage_data_918;
logic pong_storage_data_918;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_918 <= 1'b0;
        pong_storage_data_918 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                536 / IN_WIDTH: ping_storage_data_918 <= (fillup_transition == 1'b1) ? i_input_data[536 % IN_WIDTH] : ping_storage_data_918 ^ i_input_data[536 % IN_WIDTH];
                763 / IN_WIDTH: ping_storage_data_918 <= (fillup_transition == 1'b1) ? i_input_data[763 % IN_WIDTH] : ping_storage_data_918 ^ i_input_data[763 % IN_WIDTH];
                1040 / IN_WIDTH: ping_storage_data_918 <= (fillup_transition == 1'b1) ? i_input_data[1040 % IN_WIDTH] : ping_storage_data_918 ^ i_input_data[1040 % IN_WIDTH];
                1134 / IN_WIDTH: ping_storage_data_918 <= (fillup_transition == 1'b1) ? i_input_data[1134 % IN_WIDTH] : ping_storage_data_918 ^ i_input_data[1134 % IN_WIDTH];
                default: ping_storage_data_918 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_918;
                endcase
            end else begin
                case (input_count)
                536 / IN_WIDTH: pong_storage_data_918 <= (fillup_transition == 1'b1) ? i_input_data[536 % IN_WIDTH] : pong_storage_data_918 ^ i_input_data[536 % IN_WIDTH];
                763 / IN_WIDTH: pong_storage_data_918 <= (fillup_transition == 1'b1) ? i_input_data[763 % IN_WIDTH] : pong_storage_data_918 ^ i_input_data[763 % IN_WIDTH];
                1040 / IN_WIDTH: pong_storage_data_918 <= (fillup_transition == 1'b1) ? i_input_data[1040 % IN_WIDTH] : pong_storage_data_918 ^ i_input_data[1040 % IN_WIDTH];
                1134 / IN_WIDTH: pong_storage_data_918 <= (fillup_transition == 1'b1) ? i_input_data[1134 % IN_WIDTH] : pong_storage_data_918 ^ i_input_data[1134 % IN_WIDTH];
                default: pong_storage_data_918 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_918;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_918 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_918;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_918 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_918;
            end
        end
    end
end

logic ping_storage_data_919;
logic pong_storage_data_919;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_919 <= 1'b0;
        pong_storage_data_919 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                537 / IN_WIDTH: ping_storage_data_919 <= (fillup_transition == 1'b1) ? i_input_data[537 % IN_WIDTH] : ping_storage_data_919 ^ i_input_data[537 % IN_WIDTH];
                764 / IN_WIDTH: ping_storage_data_919 <= (fillup_transition == 1'b1) ? i_input_data[764 % IN_WIDTH] : ping_storage_data_919 ^ i_input_data[764 % IN_WIDTH];
                1041 / IN_WIDTH: ping_storage_data_919 <= (fillup_transition == 1'b1) ? i_input_data[1041 % IN_WIDTH] : ping_storage_data_919 ^ i_input_data[1041 % IN_WIDTH];
                1135 / IN_WIDTH: ping_storage_data_919 <= (fillup_transition == 1'b1) ? i_input_data[1135 % IN_WIDTH] : ping_storage_data_919 ^ i_input_data[1135 % IN_WIDTH];
                default: ping_storage_data_919 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_919;
                endcase
            end else begin
                case (input_count)
                537 / IN_WIDTH: pong_storage_data_919 <= (fillup_transition == 1'b1) ? i_input_data[537 % IN_WIDTH] : pong_storage_data_919 ^ i_input_data[537 % IN_WIDTH];
                764 / IN_WIDTH: pong_storage_data_919 <= (fillup_transition == 1'b1) ? i_input_data[764 % IN_WIDTH] : pong_storage_data_919 ^ i_input_data[764 % IN_WIDTH];
                1041 / IN_WIDTH: pong_storage_data_919 <= (fillup_transition == 1'b1) ? i_input_data[1041 % IN_WIDTH] : pong_storage_data_919 ^ i_input_data[1041 % IN_WIDTH];
                1135 / IN_WIDTH: pong_storage_data_919 <= (fillup_transition == 1'b1) ? i_input_data[1135 % IN_WIDTH] : pong_storage_data_919 ^ i_input_data[1135 % IN_WIDTH];
                default: pong_storage_data_919 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_919;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_919 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_919;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_919 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_919;
            end
        end
    end
end

logic ping_storage_data_920;
logic pong_storage_data_920;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_920 <= 1'b0;
        pong_storage_data_920 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                538 / IN_WIDTH: ping_storage_data_920 <= (fillup_transition == 1'b1) ? i_input_data[538 % IN_WIDTH] : ping_storage_data_920 ^ i_input_data[538 % IN_WIDTH];
                765 / IN_WIDTH: ping_storage_data_920 <= (fillup_transition == 1'b1) ? i_input_data[765 % IN_WIDTH] : ping_storage_data_920 ^ i_input_data[765 % IN_WIDTH];
                1042 / IN_WIDTH: ping_storage_data_920 <= (fillup_transition == 1'b1) ? i_input_data[1042 % IN_WIDTH] : ping_storage_data_920 ^ i_input_data[1042 % IN_WIDTH];
                1136 / IN_WIDTH: ping_storage_data_920 <= (fillup_transition == 1'b1) ? i_input_data[1136 % IN_WIDTH] : ping_storage_data_920 ^ i_input_data[1136 % IN_WIDTH];
                default: ping_storage_data_920 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_920;
                endcase
            end else begin
                case (input_count)
                538 / IN_WIDTH: pong_storage_data_920 <= (fillup_transition == 1'b1) ? i_input_data[538 % IN_WIDTH] : pong_storage_data_920 ^ i_input_data[538 % IN_WIDTH];
                765 / IN_WIDTH: pong_storage_data_920 <= (fillup_transition == 1'b1) ? i_input_data[765 % IN_WIDTH] : pong_storage_data_920 ^ i_input_data[765 % IN_WIDTH];
                1042 / IN_WIDTH: pong_storage_data_920 <= (fillup_transition == 1'b1) ? i_input_data[1042 % IN_WIDTH] : pong_storage_data_920 ^ i_input_data[1042 % IN_WIDTH];
                1136 / IN_WIDTH: pong_storage_data_920 <= (fillup_transition == 1'b1) ? i_input_data[1136 % IN_WIDTH] : pong_storage_data_920 ^ i_input_data[1136 % IN_WIDTH];
                default: pong_storage_data_920 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_920;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_920 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_920;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_920 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_920;
            end
        end
    end
end

logic ping_storage_data_921;
logic pong_storage_data_921;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_921 <= 1'b0;
        pong_storage_data_921 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                539 / IN_WIDTH: ping_storage_data_921 <= (fillup_transition == 1'b1) ? i_input_data[539 % IN_WIDTH] : ping_storage_data_921 ^ i_input_data[539 % IN_WIDTH];
                766 / IN_WIDTH: ping_storage_data_921 <= (fillup_transition == 1'b1) ? i_input_data[766 % IN_WIDTH] : ping_storage_data_921 ^ i_input_data[766 % IN_WIDTH];
                1043 / IN_WIDTH: ping_storage_data_921 <= (fillup_transition == 1'b1) ? i_input_data[1043 % IN_WIDTH] : ping_storage_data_921 ^ i_input_data[1043 % IN_WIDTH];
                1137 / IN_WIDTH: ping_storage_data_921 <= (fillup_transition == 1'b1) ? i_input_data[1137 % IN_WIDTH] : ping_storage_data_921 ^ i_input_data[1137 % IN_WIDTH];
                default: ping_storage_data_921 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_921;
                endcase
            end else begin
                case (input_count)
                539 / IN_WIDTH: pong_storage_data_921 <= (fillup_transition == 1'b1) ? i_input_data[539 % IN_WIDTH] : pong_storage_data_921 ^ i_input_data[539 % IN_WIDTH];
                766 / IN_WIDTH: pong_storage_data_921 <= (fillup_transition == 1'b1) ? i_input_data[766 % IN_WIDTH] : pong_storage_data_921 ^ i_input_data[766 % IN_WIDTH];
                1043 / IN_WIDTH: pong_storage_data_921 <= (fillup_transition == 1'b1) ? i_input_data[1043 % IN_WIDTH] : pong_storage_data_921 ^ i_input_data[1043 % IN_WIDTH];
                1137 / IN_WIDTH: pong_storage_data_921 <= (fillup_transition == 1'b1) ? i_input_data[1137 % IN_WIDTH] : pong_storage_data_921 ^ i_input_data[1137 % IN_WIDTH];
                default: pong_storage_data_921 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_921;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_921 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_921;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_921 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_921;
            end
        end
    end
end

logic ping_storage_data_922;
logic pong_storage_data_922;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_922 <= 1'b0;
        pong_storage_data_922 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                540 / IN_WIDTH: ping_storage_data_922 <= (fillup_transition == 1'b1) ? i_input_data[540 % IN_WIDTH] : ping_storage_data_922 ^ i_input_data[540 % IN_WIDTH];
                767 / IN_WIDTH: ping_storage_data_922 <= (fillup_transition == 1'b1) ? i_input_data[767 % IN_WIDTH] : ping_storage_data_922 ^ i_input_data[767 % IN_WIDTH];
                1044 / IN_WIDTH: ping_storage_data_922 <= (fillup_transition == 1'b1) ? i_input_data[1044 % IN_WIDTH] : ping_storage_data_922 ^ i_input_data[1044 % IN_WIDTH];
                1138 / IN_WIDTH: ping_storage_data_922 <= (fillup_transition == 1'b1) ? i_input_data[1138 % IN_WIDTH] : ping_storage_data_922 ^ i_input_data[1138 % IN_WIDTH];
                default: ping_storage_data_922 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_922;
                endcase
            end else begin
                case (input_count)
                540 / IN_WIDTH: pong_storage_data_922 <= (fillup_transition == 1'b1) ? i_input_data[540 % IN_WIDTH] : pong_storage_data_922 ^ i_input_data[540 % IN_WIDTH];
                767 / IN_WIDTH: pong_storage_data_922 <= (fillup_transition == 1'b1) ? i_input_data[767 % IN_WIDTH] : pong_storage_data_922 ^ i_input_data[767 % IN_WIDTH];
                1044 / IN_WIDTH: pong_storage_data_922 <= (fillup_transition == 1'b1) ? i_input_data[1044 % IN_WIDTH] : pong_storage_data_922 ^ i_input_data[1044 % IN_WIDTH];
                1138 / IN_WIDTH: pong_storage_data_922 <= (fillup_transition == 1'b1) ? i_input_data[1138 % IN_WIDTH] : pong_storage_data_922 ^ i_input_data[1138 % IN_WIDTH];
                default: pong_storage_data_922 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_922;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_922 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_922;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_922 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_922;
            end
        end
    end
end

logic ping_storage_data_923;
logic pong_storage_data_923;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_923 <= 1'b0;
        pong_storage_data_923 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                541 / IN_WIDTH: ping_storage_data_923 <= (fillup_transition == 1'b1) ? i_input_data[541 % IN_WIDTH] : ping_storage_data_923 ^ i_input_data[541 % IN_WIDTH];
                672 / IN_WIDTH: ping_storage_data_923 <= (fillup_transition == 1'b1) ? i_input_data[672 % IN_WIDTH] : ping_storage_data_923 ^ i_input_data[672 % IN_WIDTH];
                1045 / IN_WIDTH: ping_storage_data_923 <= (fillup_transition == 1'b1) ? i_input_data[1045 % IN_WIDTH] : ping_storage_data_923 ^ i_input_data[1045 % IN_WIDTH];
                1139 / IN_WIDTH: ping_storage_data_923 <= (fillup_transition == 1'b1) ? i_input_data[1139 % IN_WIDTH] : ping_storage_data_923 ^ i_input_data[1139 % IN_WIDTH];
                default: ping_storage_data_923 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_923;
                endcase
            end else begin
                case (input_count)
                541 / IN_WIDTH: pong_storage_data_923 <= (fillup_transition == 1'b1) ? i_input_data[541 % IN_WIDTH] : pong_storage_data_923 ^ i_input_data[541 % IN_WIDTH];
                672 / IN_WIDTH: pong_storage_data_923 <= (fillup_transition == 1'b1) ? i_input_data[672 % IN_WIDTH] : pong_storage_data_923 ^ i_input_data[672 % IN_WIDTH];
                1045 / IN_WIDTH: pong_storage_data_923 <= (fillup_transition == 1'b1) ? i_input_data[1045 % IN_WIDTH] : pong_storage_data_923 ^ i_input_data[1045 % IN_WIDTH];
                1139 / IN_WIDTH: pong_storage_data_923 <= (fillup_transition == 1'b1) ? i_input_data[1139 % IN_WIDTH] : pong_storage_data_923 ^ i_input_data[1139 % IN_WIDTH];
                default: pong_storage_data_923 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_923;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_923 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_923;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_923 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_923;
            end
        end
    end
end

logic ping_storage_data_924;
logic pong_storage_data_924;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_924 <= 1'b0;
        pong_storage_data_924 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                542 / IN_WIDTH: ping_storage_data_924 <= (fillup_transition == 1'b1) ? i_input_data[542 % IN_WIDTH] : ping_storage_data_924 ^ i_input_data[542 % IN_WIDTH];
                673 / IN_WIDTH: ping_storage_data_924 <= (fillup_transition == 1'b1) ? i_input_data[673 % IN_WIDTH] : ping_storage_data_924 ^ i_input_data[673 % IN_WIDTH];
                1046 / IN_WIDTH: ping_storage_data_924 <= (fillup_transition == 1'b1) ? i_input_data[1046 % IN_WIDTH] : ping_storage_data_924 ^ i_input_data[1046 % IN_WIDTH];
                1140 / IN_WIDTH: ping_storage_data_924 <= (fillup_transition == 1'b1) ? i_input_data[1140 % IN_WIDTH] : ping_storage_data_924 ^ i_input_data[1140 % IN_WIDTH];
                default: ping_storage_data_924 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_924;
                endcase
            end else begin
                case (input_count)
                542 / IN_WIDTH: pong_storage_data_924 <= (fillup_transition == 1'b1) ? i_input_data[542 % IN_WIDTH] : pong_storage_data_924 ^ i_input_data[542 % IN_WIDTH];
                673 / IN_WIDTH: pong_storage_data_924 <= (fillup_transition == 1'b1) ? i_input_data[673 % IN_WIDTH] : pong_storage_data_924 ^ i_input_data[673 % IN_WIDTH];
                1046 / IN_WIDTH: pong_storage_data_924 <= (fillup_transition == 1'b1) ? i_input_data[1046 % IN_WIDTH] : pong_storage_data_924 ^ i_input_data[1046 % IN_WIDTH];
                1140 / IN_WIDTH: pong_storage_data_924 <= (fillup_transition == 1'b1) ? i_input_data[1140 % IN_WIDTH] : pong_storage_data_924 ^ i_input_data[1140 % IN_WIDTH];
                default: pong_storage_data_924 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_924;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_924 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_924;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_924 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_924;
            end
        end
    end
end

logic ping_storage_data_925;
logic pong_storage_data_925;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_925 <= 1'b0;
        pong_storage_data_925 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                543 / IN_WIDTH: ping_storage_data_925 <= (fillup_transition == 1'b1) ? i_input_data[543 % IN_WIDTH] : ping_storage_data_925 ^ i_input_data[543 % IN_WIDTH];
                674 / IN_WIDTH: ping_storage_data_925 <= (fillup_transition == 1'b1) ? i_input_data[674 % IN_WIDTH] : ping_storage_data_925 ^ i_input_data[674 % IN_WIDTH];
                1047 / IN_WIDTH: ping_storage_data_925 <= (fillup_transition == 1'b1) ? i_input_data[1047 % IN_WIDTH] : ping_storage_data_925 ^ i_input_data[1047 % IN_WIDTH];
                1141 / IN_WIDTH: ping_storage_data_925 <= (fillup_transition == 1'b1) ? i_input_data[1141 % IN_WIDTH] : ping_storage_data_925 ^ i_input_data[1141 % IN_WIDTH];
                default: ping_storage_data_925 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_925;
                endcase
            end else begin
                case (input_count)
                543 / IN_WIDTH: pong_storage_data_925 <= (fillup_transition == 1'b1) ? i_input_data[543 % IN_WIDTH] : pong_storage_data_925 ^ i_input_data[543 % IN_WIDTH];
                674 / IN_WIDTH: pong_storage_data_925 <= (fillup_transition == 1'b1) ? i_input_data[674 % IN_WIDTH] : pong_storage_data_925 ^ i_input_data[674 % IN_WIDTH];
                1047 / IN_WIDTH: pong_storage_data_925 <= (fillup_transition == 1'b1) ? i_input_data[1047 % IN_WIDTH] : pong_storage_data_925 ^ i_input_data[1047 % IN_WIDTH];
                1141 / IN_WIDTH: pong_storage_data_925 <= (fillup_transition == 1'b1) ? i_input_data[1141 % IN_WIDTH] : pong_storage_data_925 ^ i_input_data[1141 % IN_WIDTH];
                default: pong_storage_data_925 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_925;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_925 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_925;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_925 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_925;
            end
        end
    end
end

logic ping_storage_data_926;
logic pong_storage_data_926;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_926 <= 1'b0;
        pong_storage_data_926 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                544 / IN_WIDTH: ping_storage_data_926 <= (fillup_transition == 1'b1) ? i_input_data[544 % IN_WIDTH] : ping_storage_data_926 ^ i_input_data[544 % IN_WIDTH];
                675 / IN_WIDTH: ping_storage_data_926 <= (fillup_transition == 1'b1) ? i_input_data[675 % IN_WIDTH] : ping_storage_data_926 ^ i_input_data[675 % IN_WIDTH];
                1048 / IN_WIDTH: ping_storage_data_926 <= (fillup_transition == 1'b1) ? i_input_data[1048 % IN_WIDTH] : ping_storage_data_926 ^ i_input_data[1048 % IN_WIDTH];
                1142 / IN_WIDTH: ping_storage_data_926 <= (fillup_transition == 1'b1) ? i_input_data[1142 % IN_WIDTH] : ping_storage_data_926 ^ i_input_data[1142 % IN_WIDTH];
                default: ping_storage_data_926 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_926;
                endcase
            end else begin
                case (input_count)
                544 / IN_WIDTH: pong_storage_data_926 <= (fillup_transition == 1'b1) ? i_input_data[544 % IN_WIDTH] : pong_storage_data_926 ^ i_input_data[544 % IN_WIDTH];
                675 / IN_WIDTH: pong_storage_data_926 <= (fillup_transition == 1'b1) ? i_input_data[675 % IN_WIDTH] : pong_storage_data_926 ^ i_input_data[675 % IN_WIDTH];
                1048 / IN_WIDTH: pong_storage_data_926 <= (fillup_transition == 1'b1) ? i_input_data[1048 % IN_WIDTH] : pong_storage_data_926 ^ i_input_data[1048 % IN_WIDTH];
                1142 / IN_WIDTH: pong_storage_data_926 <= (fillup_transition == 1'b1) ? i_input_data[1142 % IN_WIDTH] : pong_storage_data_926 ^ i_input_data[1142 % IN_WIDTH];
                default: pong_storage_data_926 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_926;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_926 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_926;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_926 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_926;
            end
        end
    end
end

logic ping_storage_data_927;
logic pong_storage_data_927;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_927 <= 1'b0;
        pong_storage_data_927 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                545 / IN_WIDTH: ping_storage_data_927 <= (fillup_transition == 1'b1) ? i_input_data[545 % IN_WIDTH] : ping_storage_data_927 ^ i_input_data[545 % IN_WIDTH];
                676 / IN_WIDTH: ping_storage_data_927 <= (fillup_transition == 1'b1) ? i_input_data[676 % IN_WIDTH] : ping_storage_data_927 ^ i_input_data[676 % IN_WIDTH];
                1049 / IN_WIDTH: ping_storage_data_927 <= (fillup_transition == 1'b1) ? i_input_data[1049 % IN_WIDTH] : ping_storage_data_927 ^ i_input_data[1049 % IN_WIDTH];
                1143 / IN_WIDTH: ping_storage_data_927 <= (fillup_transition == 1'b1) ? i_input_data[1143 % IN_WIDTH] : ping_storage_data_927 ^ i_input_data[1143 % IN_WIDTH];
                default: ping_storage_data_927 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_927;
                endcase
            end else begin
                case (input_count)
                545 / IN_WIDTH: pong_storage_data_927 <= (fillup_transition == 1'b1) ? i_input_data[545 % IN_WIDTH] : pong_storage_data_927 ^ i_input_data[545 % IN_WIDTH];
                676 / IN_WIDTH: pong_storage_data_927 <= (fillup_transition == 1'b1) ? i_input_data[676 % IN_WIDTH] : pong_storage_data_927 ^ i_input_data[676 % IN_WIDTH];
                1049 / IN_WIDTH: pong_storage_data_927 <= (fillup_transition == 1'b1) ? i_input_data[1049 % IN_WIDTH] : pong_storage_data_927 ^ i_input_data[1049 % IN_WIDTH];
                1143 / IN_WIDTH: pong_storage_data_927 <= (fillup_transition == 1'b1) ? i_input_data[1143 % IN_WIDTH] : pong_storage_data_927 ^ i_input_data[1143 % IN_WIDTH];
                default: pong_storage_data_927 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_927;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_927 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_927;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_927 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_927;
            end
        end
    end
end

logic ping_storage_data_928;
logic pong_storage_data_928;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_928 <= 1'b0;
        pong_storage_data_928 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                546 / IN_WIDTH: ping_storage_data_928 <= (fillup_transition == 1'b1) ? i_input_data[546 % IN_WIDTH] : ping_storage_data_928 ^ i_input_data[546 % IN_WIDTH];
                677 / IN_WIDTH: ping_storage_data_928 <= (fillup_transition == 1'b1) ? i_input_data[677 % IN_WIDTH] : ping_storage_data_928 ^ i_input_data[677 % IN_WIDTH];
                1050 / IN_WIDTH: ping_storage_data_928 <= (fillup_transition == 1'b1) ? i_input_data[1050 % IN_WIDTH] : ping_storage_data_928 ^ i_input_data[1050 % IN_WIDTH];
                1144 / IN_WIDTH: ping_storage_data_928 <= (fillup_transition == 1'b1) ? i_input_data[1144 % IN_WIDTH] : ping_storage_data_928 ^ i_input_data[1144 % IN_WIDTH];
                default: ping_storage_data_928 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_928;
                endcase
            end else begin
                case (input_count)
                546 / IN_WIDTH: pong_storage_data_928 <= (fillup_transition == 1'b1) ? i_input_data[546 % IN_WIDTH] : pong_storage_data_928 ^ i_input_data[546 % IN_WIDTH];
                677 / IN_WIDTH: pong_storage_data_928 <= (fillup_transition == 1'b1) ? i_input_data[677 % IN_WIDTH] : pong_storage_data_928 ^ i_input_data[677 % IN_WIDTH];
                1050 / IN_WIDTH: pong_storage_data_928 <= (fillup_transition == 1'b1) ? i_input_data[1050 % IN_WIDTH] : pong_storage_data_928 ^ i_input_data[1050 % IN_WIDTH];
                1144 / IN_WIDTH: pong_storage_data_928 <= (fillup_transition == 1'b1) ? i_input_data[1144 % IN_WIDTH] : pong_storage_data_928 ^ i_input_data[1144 % IN_WIDTH];
                default: pong_storage_data_928 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_928;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_928 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_928;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_928 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_928;
            end
        end
    end
end

logic ping_storage_data_929;
logic pong_storage_data_929;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_929 <= 1'b0;
        pong_storage_data_929 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                547 / IN_WIDTH: ping_storage_data_929 <= (fillup_transition == 1'b1) ? i_input_data[547 % IN_WIDTH] : ping_storage_data_929 ^ i_input_data[547 % IN_WIDTH];
                678 / IN_WIDTH: ping_storage_data_929 <= (fillup_transition == 1'b1) ? i_input_data[678 % IN_WIDTH] : ping_storage_data_929 ^ i_input_data[678 % IN_WIDTH];
                1051 / IN_WIDTH: ping_storage_data_929 <= (fillup_transition == 1'b1) ? i_input_data[1051 % IN_WIDTH] : ping_storage_data_929 ^ i_input_data[1051 % IN_WIDTH];
                1145 / IN_WIDTH: ping_storage_data_929 <= (fillup_transition == 1'b1) ? i_input_data[1145 % IN_WIDTH] : ping_storage_data_929 ^ i_input_data[1145 % IN_WIDTH];
                default: ping_storage_data_929 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_929;
                endcase
            end else begin
                case (input_count)
                547 / IN_WIDTH: pong_storage_data_929 <= (fillup_transition == 1'b1) ? i_input_data[547 % IN_WIDTH] : pong_storage_data_929 ^ i_input_data[547 % IN_WIDTH];
                678 / IN_WIDTH: pong_storage_data_929 <= (fillup_transition == 1'b1) ? i_input_data[678 % IN_WIDTH] : pong_storage_data_929 ^ i_input_data[678 % IN_WIDTH];
                1051 / IN_WIDTH: pong_storage_data_929 <= (fillup_transition == 1'b1) ? i_input_data[1051 % IN_WIDTH] : pong_storage_data_929 ^ i_input_data[1051 % IN_WIDTH];
                1145 / IN_WIDTH: pong_storage_data_929 <= (fillup_transition == 1'b1) ? i_input_data[1145 % IN_WIDTH] : pong_storage_data_929 ^ i_input_data[1145 % IN_WIDTH];
                default: pong_storage_data_929 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_929;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_929 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_929;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_929 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_929;
            end
        end
    end
end

logic ping_storage_data_930;
logic pong_storage_data_930;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_930 <= 1'b0;
        pong_storage_data_930 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                548 / IN_WIDTH: ping_storage_data_930 <= (fillup_transition == 1'b1) ? i_input_data[548 % IN_WIDTH] : ping_storage_data_930 ^ i_input_data[548 % IN_WIDTH];
                679 / IN_WIDTH: ping_storage_data_930 <= (fillup_transition == 1'b1) ? i_input_data[679 % IN_WIDTH] : ping_storage_data_930 ^ i_input_data[679 % IN_WIDTH];
                1052 / IN_WIDTH: ping_storage_data_930 <= (fillup_transition == 1'b1) ? i_input_data[1052 % IN_WIDTH] : ping_storage_data_930 ^ i_input_data[1052 % IN_WIDTH];
                1146 / IN_WIDTH: ping_storage_data_930 <= (fillup_transition == 1'b1) ? i_input_data[1146 % IN_WIDTH] : ping_storage_data_930 ^ i_input_data[1146 % IN_WIDTH];
                default: ping_storage_data_930 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_930;
                endcase
            end else begin
                case (input_count)
                548 / IN_WIDTH: pong_storage_data_930 <= (fillup_transition == 1'b1) ? i_input_data[548 % IN_WIDTH] : pong_storage_data_930 ^ i_input_data[548 % IN_WIDTH];
                679 / IN_WIDTH: pong_storage_data_930 <= (fillup_transition == 1'b1) ? i_input_data[679 % IN_WIDTH] : pong_storage_data_930 ^ i_input_data[679 % IN_WIDTH];
                1052 / IN_WIDTH: pong_storage_data_930 <= (fillup_transition == 1'b1) ? i_input_data[1052 % IN_WIDTH] : pong_storage_data_930 ^ i_input_data[1052 % IN_WIDTH];
                1146 / IN_WIDTH: pong_storage_data_930 <= (fillup_transition == 1'b1) ? i_input_data[1146 % IN_WIDTH] : pong_storage_data_930 ^ i_input_data[1146 % IN_WIDTH];
                default: pong_storage_data_930 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_930;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_930 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_930;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_930 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_930;
            end
        end
    end
end

logic ping_storage_data_931;
logic pong_storage_data_931;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_931 <= 1'b0;
        pong_storage_data_931 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                549 / IN_WIDTH: ping_storage_data_931 <= (fillup_transition == 1'b1) ? i_input_data[549 % IN_WIDTH] : ping_storage_data_931 ^ i_input_data[549 % IN_WIDTH];
                680 / IN_WIDTH: ping_storage_data_931 <= (fillup_transition == 1'b1) ? i_input_data[680 % IN_WIDTH] : ping_storage_data_931 ^ i_input_data[680 % IN_WIDTH];
                1053 / IN_WIDTH: ping_storage_data_931 <= (fillup_transition == 1'b1) ? i_input_data[1053 % IN_WIDTH] : ping_storage_data_931 ^ i_input_data[1053 % IN_WIDTH];
                1147 / IN_WIDTH: ping_storage_data_931 <= (fillup_transition == 1'b1) ? i_input_data[1147 % IN_WIDTH] : ping_storage_data_931 ^ i_input_data[1147 % IN_WIDTH];
                default: ping_storage_data_931 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_931;
                endcase
            end else begin
                case (input_count)
                549 / IN_WIDTH: pong_storage_data_931 <= (fillup_transition == 1'b1) ? i_input_data[549 % IN_WIDTH] : pong_storage_data_931 ^ i_input_data[549 % IN_WIDTH];
                680 / IN_WIDTH: pong_storage_data_931 <= (fillup_transition == 1'b1) ? i_input_data[680 % IN_WIDTH] : pong_storage_data_931 ^ i_input_data[680 % IN_WIDTH];
                1053 / IN_WIDTH: pong_storage_data_931 <= (fillup_transition == 1'b1) ? i_input_data[1053 % IN_WIDTH] : pong_storage_data_931 ^ i_input_data[1053 % IN_WIDTH];
                1147 / IN_WIDTH: pong_storage_data_931 <= (fillup_transition == 1'b1) ? i_input_data[1147 % IN_WIDTH] : pong_storage_data_931 ^ i_input_data[1147 % IN_WIDTH];
                default: pong_storage_data_931 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_931;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_931 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_931;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_931 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_931;
            end
        end
    end
end

logic ping_storage_data_932;
logic pong_storage_data_932;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_932 <= 1'b0;
        pong_storage_data_932 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                550 / IN_WIDTH: ping_storage_data_932 <= (fillup_transition == 1'b1) ? i_input_data[550 % IN_WIDTH] : ping_storage_data_932 ^ i_input_data[550 % IN_WIDTH];
                681 / IN_WIDTH: ping_storage_data_932 <= (fillup_transition == 1'b1) ? i_input_data[681 % IN_WIDTH] : ping_storage_data_932 ^ i_input_data[681 % IN_WIDTH];
                1054 / IN_WIDTH: ping_storage_data_932 <= (fillup_transition == 1'b1) ? i_input_data[1054 % IN_WIDTH] : ping_storage_data_932 ^ i_input_data[1054 % IN_WIDTH];
                1148 / IN_WIDTH: ping_storage_data_932 <= (fillup_transition == 1'b1) ? i_input_data[1148 % IN_WIDTH] : ping_storage_data_932 ^ i_input_data[1148 % IN_WIDTH];
                default: ping_storage_data_932 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_932;
                endcase
            end else begin
                case (input_count)
                550 / IN_WIDTH: pong_storage_data_932 <= (fillup_transition == 1'b1) ? i_input_data[550 % IN_WIDTH] : pong_storage_data_932 ^ i_input_data[550 % IN_WIDTH];
                681 / IN_WIDTH: pong_storage_data_932 <= (fillup_transition == 1'b1) ? i_input_data[681 % IN_WIDTH] : pong_storage_data_932 ^ i_input_data[681 % IN_WIDTH];
                1054 / IN_WIDTH: pong_storage_data_932 <= (fillup_transition == 1'b1) ? i_input_data[1054 % IN_WIDTH] : pong_storage_data_932 ^ i_input_data[1054 % IN_WIDTH];
                1148 / IN_WIDTH: pong_storage_data_932 <= (fillup_transition == 1'b1) ? i_input_data[1148 % IN_WIDTH] : pong_storage_data_932 ^ i_input_data[1148 % IN_WIDTH];
                default: pong_storage_data_932 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_932;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_932 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_932;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_932 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_932;
            end
        end
    end
end

logic ping_storage_data_933;
logic pong_storage_data_933;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_933 <= 1'b0;
        pong_storage_data_933 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                551 / IN_WIDTH: ping_storage_data_933 <= (fillup_transition == 1'b1) ? i_input_data[551 % IN_WIDTH] : ping_storage_data_933 ^ i_input_data[551 % IN_WIDTH];
                682 / IN_WIDTH: ping_storage_data_933 <= (fillup_transition == 1'b1) ? i_input_data[682 % IN_WIDTH] : ping_storage_data_933 ^ i_input_data[682 % IN_WIDTH];
                1055 / IN_WIDTH: ping_storage_data_933 <= (fillup_transition == 1'b1) ? i_input_data[1055 % IN_WIDTH] : ping_storage_data_933 ^ i_input_data[1055 % IN_WIDTH];
                1149 / IN_WIDTH: ping_storage_data_933 <= (fillup_transition == 1'b1) ? i_input_data[1149 % IN_WIDTH] : ping_storage_data_933 ^ i_input_data[1149 % IN_WIDTH];
                default: ping_storage_data_933 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_933;
                endcase
            end else begin
                case (input_count)
                551 / IN_WIDTH: pong_storage_data_933 <= (fillup_transition == 1'b1) ? i_input_data[551 % IN_WIDTH] : pong_storage_data_933 ^ i_input_data[551 % IN_WIDTH];
                682 / IN_WIDTH: pong_storage_data_933 <= (fillup_transition == 1'b1) ? i_input_data[682 % IN_WIDTH] : pong_storage_data_933 ^ i_input_data[682 % IN_WIDTH];
                1055 / IN_WIDTH: pong_storage_data_933 <= (fillup_transition == 1'b1) ? i_input_data[1055 % IN_WIDTH] : pong_storage_data_933 ^ i_input_data[1055 % IN_WIDTH];
                1149 / IN_WIDTH: pong_storage_data_933 <= (fillup_transition == 1'b1) ? i_input_data[1149 % IN_WIDTH] : pong_storage_data_933 ^ i_input_data[1149 % IN_WIDTH];
                default: pong_storage_data_933 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_933;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_933 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_933;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_933 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_933;
            end
        end
    end
end

logic ping_storage_data_934;
logic pong_storage_data_934;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_934 <= 1'b0;
        pong_storage_data_934 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                552 / IN_WIDTH: ping_storage_data_934 <= (fillup_transition == 1'b1) ? i_input_data[552 % IN_WIDTH] : ping_storage_data_934 ^ i_input_data[552 % IN_WIDTH];
                683 / IN_WIDTH: ping_storage_data_934 <= (fillup_transition == 1'b1) ? i_input_data[683 % IN_WIDTH] : ping_storage_data_934 ^ i_input_data[683 % IN_WIDTH];
                960 / IN_WIDTH: ping_storage_data_934 <= (fillup_transition == 1'b1) ? i_input_data[960 % IN_WIDTH] : ping_storage_data_934 ^ i_input_data[960 % IN_WIDTH];
                1150 / IN_WIDTH: ping_storage_data_934 <= (fillup_transition == 1'b1) ? i_input_data[1150 % IN_WIDTH] : ping_storage_data_934 ^ i_input_data[1150 % IN_WIDTH];
                default: ping_storage_data_934 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_934;
                endcase
            end else begin
                case (input_count)
                552 / IN_WIDTH: pong_storage_data_934 <= (fillup_transition == 1'b1) ? i_input_data[552 % IN_WIDTH] : pong_storage_data_934 ^ i_input_data[552 % IN_WIDTH];
                683 / IN_WIDTH: pong_storage_data_934 <= (fillup_transition == 1'b1) ? i_input_data[683 % IN_WIDTH] : pong_storage_data_934 ^ i_input_data[683 % IN_WIDTH];
                960 / IN_WIDTH: pong_storage_data_934 <= (fillup_transition == 1'b1) ? i_input_data[960 % IN_WIDTH] : pong_storage_data_934 ^ i_input_data[960 % IN_WIDTH];
                1150 / IN_WIDTH: pong_storage_data_934 <= (fillup_transition == 1'b1) ? i_input_data[1150 % IN_WIDTH] : pong_storage_data_934 ^ i_input_data[1150 % IN_WIDTH];
                default: pong_storage_data_934 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_934;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_934 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_934;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_934 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_934;
            end
        end
    end
end

logic ping_storage_data_935;
logic pong_storage_data_935;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_935 <= 1'b0;
        pong_storage_data_935 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                553 / IN_WIDTH: ping_storage_data_935 <= (fillup_transition == 1'b1) ? i_input_data[553 % IN_WIDTH] : ping_storage_data_935 ^ i_input_data[553 % IN_WIDTH];
                684 / IN_WIDTH: ping_storage_data_935 <= (fillup_transition == 1'b1) ? i_input_data[684 % IN_WIDTH] : ping_storage_data_935 ^ i_input_data[684 % IN_WIDTH];
                961 / IN_WIDTH: ping_storage_data_935 <= (fillup_transition == 1'b1) ? i_input_data[961 % IN_WIDTH] : ping_storage_data_935 ^ i_input_data[961 % IN_WIDTH];
                1151 / IN_WIDTH: ping_storage_data_935 <= (fillup_transition == 1'b1) ? i_input_data[1151 % IN_WIDTH] : ping_storage_data_935 ^ i_input_data[1151 % IN_WIDTH];
                default: ping_storage_data_935 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_935;
                endcase
            end else begin
                case (input_count)
                553 / IN_WIDTH: pong_storage_data_935 <= (fillup_transition == 1'b1) ? i_input_data[553 % IN_WIDTH] : pong_storage_data_935 ^ i_input_data[553 % IN_WIDTH];
                684 / IN_WIDTH: pong_storage_data_935 <= (fillup_transition == 1'b1) ? i_input_data[684 % IN_WIDTH] : pong_storage_data_935 ^ i_input_data[684 % IN_WIDTH];
                961 / IN_WIDTH: pong_storage_data_935 <= (fillup_transition == 1'b1) ? i_input_data[961 % IN_WIDTH] : pong_storage_data_935 ^ i_input_data[961 % IN_WIDTH];
                1151 / IN_WIDTH: pong_storage_data_935 <= (fillup_transition == 1'b1) ? i_input_data[1151 % IN_WIDTH] : pong_storage_data_935 ^ i_input_data[1151 % IN_WIDTH];
                default: pong_storage_data_935 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_935;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_935 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_935;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_935 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_935;
            end
        end
    end
end

logic ping_storage_data_936;
logic pong_storage_data_936;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_936 <= 1'b0;
        pong_storage_data_936 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                554 / IN_WIDTH: ping_storage_data_936 <= (fillup_transition == 1'b1) ? i_input_data[554 % IN_WIDTH] : ping_storage_data_936 ^ i_input_data[554 % IN_WIDTH];
                685 / IN_WIDTH: ping_storage_data_936 <= (fillup_transition == 1'b1) ? i_input_data[685 % IN_WIDTH] : ping_storage_data_936 ^ i_input_data[685 % IN_WIDTH];
                962 / IN_WIDTH: ping_storage_data_936 <= (fillup_transition == 1'b1) ? i_input_data[962 % IN_WIDTH] : ping_storage_data_936 ^ i_input_data[962 % IN_WIDTH];
                1056 / IN_WIDTH: ping_storage_data_936 <= (fillup_transition == 1'b1) ? i_input_data[1056 % IN_WIDTH] : ping_storage_data_936 ^ i_input_data[1056 % IN_WIDTH];
                default: ping_storage_data_936 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_936;
                endcase
            end else begin
                case (input_count)
                554 / IN_WIDTH: pong_storage_data_936 <= (fillup_transition == 1'b1) ? i_input_data[554 % IN_WIDTH] : pong_storage_data_936 ^ i_input_data[554 % IN_WIDTH];
                685 / IN_WIDTH: pong_storage_data_936 <= (fillup_transition == 1'b1) ? i_input_data[685 % IN_WIDTH] : pong_storage_data_936 ^ i_input_data[685 % IN_WIDTH];
                962 / IN_WIDTH: pong_storage_data_936 <= (fillup_transition == 1'b1) ? i_input_data[962 % IN_WIDTH] : pong_storage_data_936 ^ i_input_data[962 % IN_WIDTH];
                1056 / IN_WIDTH: pong_storage_data_936 <= (fillup_transition == 1'b1) ? i_input_data[1056 % IN_WIDTH] : pong_storage_data_936 ^ i_input_data[1056 % IN_WIDTH];
                default: pong_storage_data_936 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_936;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_936 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_936;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_936 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_936;
            end
        end
    end
end

logic ping_storage_data_937;
logic pong_storage_data_937;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_937 <= 1'b0;
        pong_storage_data_937 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                555 / IN_WIDTH: ping_storage_data_937 <= (fillup_transition == 1'b1) ? i_input_data[555 % IN_WIDTH] : ping_storage_data_937 ^ i_input_data[555 % IN_WIDTH];
                686 / IN_WIDTH: ping_storage_data_937 <= (fillup_transition == 1'b1) ? i_input_data[686 % IN_WIDTH] : ping_storage_data_937 ^ i_input_data[686 % IN_WIDTH];
                963 / IN_WIDTH: ping_storage_data_937 <= (fillup_transition == 1'b1) ? i_input_data[963 % IN_WIDTH] : ping_storage_data_937 ^ i_input_data[963 % IN_WIDTH];
                1057 / IN_WIDTH: ping_storage_data_937 <= (fillup_transition == 1'b1) ? i_input_data[1057 % IN_WIDTH] : ping_storage_data_937 ^ i_input_data[1057 % IN_WIDTH];
                default: ping_storage_data_937 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_937;
                endcase
            end else begin
                case (input_count)
                555 / IN_WIDTH: pong_storage_data_937 <= (fillup_transition == 1'b1) ? i_input_data[555 % IN_WIDTH] : pong_storage_data_937 ^ i_input_data[555 % IN_WIDTH];
                686 / IN_WIDTH: pong_storage_data_937 <= (fillup_transition == 1'b1) ? i_input_data[686 % IN_WIDTH] : pong_storage_data_937 ^ i_input_data[686 % IN_WIDTH];
                963 / IN_WIDTH: pong_storage_data_937 <= (fillup_transition == 1'b1) ? i_input_data[963 % IN_WIDTH] : pong_storage_data_937 ^ i_input_data[963 % IN_WIDTH];
                1057 / IN_WIDTH: pong_storage_data_937 <= (fillup_transition == 1'b1) ? i_input_data[1057 % IN_WIDTH] : pong_storage_data_937 ^ i_input_data[1057 % IN_WIDTH];
                default: pong_storage_data_937 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_937;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_937 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_937;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_937 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_937;
            end
        end
    end
end

logic ping_storage_data_938;
logic pong_storage_data_938;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_938 <= 1'b0;
        pong_storage_data_938 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                556 / IN_WIDTH: ping_storage_data_938 <= (fillup_transition == 1'b1) ? i_input_data[556 % IN_WIDTH] : ping_storage_data_938 ^ i_input_data[556 % IN_WIDTH];
                687 / IN_WIDTH: ping_storage_data_938 <= (fillup_transition == 1'b1) ? i_input_data[687 % IN_WIDTH] : ping_storage_data_938 ^ i_input_data[687 % IN_WIDTH];
                964 / IN_WIDTH: ping_storage_data_938 <= (fillup_transition == 1'b1) ? i_input_data[964 % IN_WIDTH] : ping_storage_data_938 ^ i_input_data[964 % IN_WIDTH];
                1058 / IN_WIDTH: ping_storage_data_938 <= (fillup_transition == 1'b1) ? i_input_data[1058 % IN_WIDTH] : ping_storage_data_938 ^ i_input_data[1058 % IN_WIDTH];
                default: ping_storage_data_938 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_938;
                endcase
            end else begin
                case (input_count)
                556 / IN_WIDTH: pong_storage_data_938 <= (fillup_transition == 1'b1) ? i_input_data[556 % IN_WIDTH] : pong_storage_data_938 ^ i_input_data[556 % IN_WIDTH];
                687 / IN_WIDTH: pong_storage_data_938 <= (fillup_transition == 1'b1) ? i_input_data[687 % IN_WIDTH] : pong_storage_data_938 ^ i_input_data[687 % IN_WIDTH];
                964 / IN_WIDTH: pong_storage_data_938 <= (fillup_transition == 1'b1) ? i_input_data[964 % IN_WIDTH] : pong_storage_data_938 ^ i_input_data[964 % IN_WIDTH];
                1058 / IN_WIDTH: pong_storage_data_938 <= (fillup_transition == 1'b1) ? i_input_data[1058 % IN_WIDTH] : pong_storage_data_938 ^ i_input_data[1058 % IN_WIDTH];
                default: pong_storage_data_938 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_938;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_938 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_938;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_938 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_938;
            end
        end
    end
end

logic ping_storage_data_939;
logic pong_storage_data_939;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_939 <= 1'b0;
        pong_storage_data_939 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                557 / IN_WIDTH: ping_storage_data_939 <= (fillup_transition == 1'b1) ? i_input_data[557 % IN_WIDTH] : ping_storage_data_939 ^ i_input_data[557 % IN_WIDTH];
                688 / IN_WIDTH: ping_storage_data_939 <= (fillup_transition == 1'b1) ? i_input_data[688 % IN_WIDTH] : ping_storage_data_939 ^ i_input_data[688 % IN_WIDTH];
                965 / IN_WIDTH: ping_storage_data_939 <= (fillup_transition == 1'b1) ? i_input_data[965 % IN_WIDTH] : ping_storage_data_939 ^ i_input_data[965 % IN_WIDTH];
                1059 / IN_WIDTH: ping_storage_data_939 <= (fillup_transition == 1'b1) ? i_input_data[1059 % IN_WIDTH] : ping_storage_data_939 ^ i_input_data[1059 % IN_WIDTH];
                default: ping_storage_data_939 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_939;
                endcase
            end else begin
                case (input_count)
                557 / IN_WIDTH: pong_storage_data_939 <= (fillup_transition == 1'b1) ? i_input_data[557 % IN_WIDTH] : pong_storage_data_939 ^ i_input_data[557 % IN_WIDTH];
                688 / IN_WIDTH: pong_storage_data_939 <= (fillup_transition == 1'b1) ? i_input_data[688 % IN_WIDTH] : pong_storage_data_939 ^ i_input_data[688 % IN_WIDTH];
                965 / IN_WIDTH: pong_storage_data_939 <= (fillup_transition == 1'b1) ? i_input_data[965 % IN_WIDTH] : pong_storage_data_939 ^ i_input_data[965 % IN_WIDTH];
                1059 / IN_WIDTH: pong_storage_data_939 <= (fillup_transition == 1'b1) ? i_input_data[1059 % IN_WIDTH] : pong_storage_data_939 ^ i_input_data[1059 % IN_WIDTH];
                default: pong_storage_data_939 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_939;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_939 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_939;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_939 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_939;
            end
        end
    end
end

logic ping_storage_data_940;
logic pong_storage_data_940;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_940 <= 1'b0;
        pong_storage_data_940 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                558 / IN_WIDTH: ping_storage_data_940 <= (fillup_transition == 1'b1) ? i_input_data[558 % IN_WIDTH] : ping_storage_data_940 ^ i_input_data[558 % IN_WIDTH];
                689 / IN_WIDTH: ping_storage_data_940 <= (fillup_transition == 1'b1) ? i_input_data[689 % IN_WIDTH] : ping_storage_data_940 ^ i_input_data[689 % IN_WIDTH];
                966 / IN_WIDTH: ping_storage_data_940 <= (fillup_transition == 1'b1) ? i_input_data[966 % IN_WIDTH] : ping_storage_data_940 ^ i_input_data[966 % IN_WIDTH];
                1060 / IN_WIDTH: ping_storage_data_940 <= (fillup_transition == 1'b1) ? i_input_data[1060 % IN_WIDTH] : ping_storage_data_940 ^ i_input_data[1060 % IN_WIDTH];
                default: ping_storage_data_940 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_940;
                endcase
            end else begin
                case (input_count)
                558 / IN_WIDTH: pong_storage_data_940 <= (fillup_transition == 1'b1) ? i_input_data[558 % IN_WIDTH] : pong_storage_data_940 ^ i_input_data[558 % IN_WIDTH];
                689 / IN_WIDTH: pong_storage_data_940 <= (fillup_transition == 1'b1) ? i_input_data[689 % IN_WIDTH] : pong_storage_data_940 ^ i_input_data[689 % IN_WIDTH];
                966 / IN_WIDTH: pong_storage_data_940 <= (fillup_transition == 1'b1) ? i_input_data[966 % IN_WIDTH] : pong_storage_data_940 ^ i_input_data[966 % IN_WIDTH];
                1060 / IN_WIDTH: pong_storage_data_940 <= (fillup_transition == 1'b1) ? i_input_data[1060 % IN_WIDTH] : pong_storage_data_940 ^ i_input_data[1060 % IN_WIDTH];
                default: pong_storage_data_940 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_940;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_940 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_940;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_940 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_940;
            end
        end
    end
end

logic ping_storage_data_941;
logic pong_storage_data_941;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_941 <= 1'b0;
        pong_storage_data_941 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                559 / IN_WIDTH: ping_storage_data_941 <= (fillup_transition == 1'b1) ? i_input_data[559 % IN_WIDTH] : ping_storage_data_941 ^ i_input_data[559 % IN_WIDTH];
                690 / IN_WIDTH: ping_storage_data_941 <= (fillup_transition == 1'b1) ? i_input_data[690 % IN_WIDTH] : ping_storage_data_941 ^ i_input_data[690 % IN_WIDTH];
                967 / IN_WIDTH: ping_storage_data_941 <= (fillup_transition == 1'b1) ? i_input_data[967 % IN_WIDTH] : ping_storage_data_941 ^ i_input_data[967 % IN_WIDTH];
                1061 / IN_WIDTH: ping_storage_data_941 <= (fillup_transition == 1'b1) ? i_input_data[1061 % IN_WIDTH] : ping_storage_data_941 ^ i_input_data[1061 % IN_WIDTH];
                default: ping_storage_data_941 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_941;
                endcase
            end else begin
                case (input_count)
                559 / IN_WIDTH: pong_storage_data_941 <= (fillup_transition == 1'b1) ? i_input_data[559 % IN_WIDTH] : pong_storage_data_941 ^ i_input_data[559 % IN_WIDTH];
                690 / IN_WIDTH: pong_storage_data_941 <= (fillup_transition == 1'b1) ? i_input_data[690 % IN_WIDTH] : pong_storage_data_941 ^ i_input_data[690 % IN_WIDTH];
                967 / IN_WIDTH: pong_storage_data_941 <= (fillup_transition == 1'b1) ? i_input_data[967 % IN_WIDTH] : pong_storage_data_941 ^ i_input_data[967 % IN_WIDTH];
                1061 / IN_WIDTH: pong_storage_data_941 <= (fillup_transition == 1'b1) ? i_input_data[1061 % IN_WIDTH] : pong_storage_data_941 ^ i_input_data[1061 % IN_WIDTH];
                default: pong_storage_data_941 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_941;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_941 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_941;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_941 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_941;
            end
        end
    end
end

logic ping_storage_data_942;
logic pong_storage_data_942;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_942 <= 1'b0;
        pong_storage_data_942 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                560 / IN_WIDTH: ping_storage_data_942 <= (fillup_transition == 1'b1) ? i_input_data[560 % IN_WIDTH] : ping_storage_data_942 ^ i_input_data[560 % IN_WIDTH];
                691 / IN_WIDTH: ping_storage_data_942 <= (fillup_transition == 1'b1) ? i_input_data[691 % IN_WIDTH] : ping_storage_data_942 ^ i_input_data[691 % IN_WIDTH];
                968 / IN_WIDTH: ping_storage_data_942 <= (fillup_transition == 1'b1) ? i_input_data[968 % IN_WIDTH] : ping_storage_data_942 ^ i_input_data[968 % IN_WIDTH];
                1062 / IN_WIDTH: ping_storage_data_942 <= (fillup_transition == 1'b1) ? i_input_data[1062 % IN_WIDTH] : ping_storage_data_942 ^ i_input_data[1062 % IN_WIDTH];
                default: ping_storage_data_942 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_942;
                endcase
            end else begin
                case (input_count)
                560 / IN_WIDTH: pong_storage_data_942 <= (fillup_transition == 1'b1) ? i_input_data[560 % IN_WIDTH] : pong_storage_data_942 ^ i_input_data[560 % IN_WIDTH];
                691 / IN_WIDTH: pong_storage_data_942 <= (fillup_transition == 1'b1) ? i_input_data[691 % IN_WIDTH] : pong_storage_data_942 ^ i_input_data[691 % IN_WIDTH];
                968 / IN_WIDTH: pong_storage_data_942 <= (fillup_transition == 1'b1) ? i_input_data[968 % IN_WIDTH] : pong_storage_data_942 ^ i_input_data[968 % IN_WIDTH];
                1062 / IN_WIDTH: pong_storage_data_942 <= (fillup_transition == 1'b1) ? i_input_data[1062 % IN_WIDTH] : pong_storage_data_942 ^ i_input_data[1062 % IN_WIDTH];
                default: pong_storage_data_942 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_942;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_942 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_942;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_942 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_942;
            end
        end
    end
end

logic ping_storage_data_943;
logic pong_storage_data_943;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_943 <= 1'b0;
        pong_storage_data_943 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                561 / IN_WIDTH: ping_storage_data_943 <= (fillup_transition == 1'b1) ? i_input_data[561 % IN_WIDTH] : ping_storage_data_943 ^ i_input_data[561 % IN_WIDTH];
                692 / IN_WIDTH: ping_storage_data_943 <= (fillup_transition == 1'b1) ? i_input_data[692 % IN_WIDTH] : ping_storage_data_943 ^ i_input_data[692 % IN_WIDTH];
                969 / IN_WIDTH: ping_storage_data_943 <= (fillup_transition == 1'b1) ? i_input_data[969 % IN_WIDTH] : ping_storage_data_943 ^ i_input_data[969 % IN_WIDTH];
                1063 / IN_WIDTH: ping_storage_data_943 <= (fillup_transition == 1'b1) ? i_input_data[1063 % IN_WIDTH] : ping_storage_data_943 ^ i_input_data[1063 % IN_WIDTH];
                default: ping_storage_data_943 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_943;
                endcase
            end else begin
                case (input_count)
                561 / IN_WIDTH: pong_storage_data_943 <= (fillup_transition == 1'b1) ? i_input_data[561 % IN_WIDTH] : pong_storage_data_943 ^ i_input_data[561 % IN_WIDTH];
                692 / IN_WIDTH: pong_storage_data_943 <= (fillup_transition == 1'b1) ? i_input_data[692 % IN_WIDTH] : pong_storage_data_943 ^ i_input_data[692 % IN_WIDTH];
                969 / IN_WIDTH: pong_storage_data_943 <= (fillup_transition == 1'b1) ? i_input_data[969 % IN_WIDTH] : pong_storage_data_943 ^ i_input_data[969 % IN_WIDTH];
                1063 / IN_WIDTH: pong_storage_data_943 <= (fillup_transition == 1'b1) ? i_input_data[1063 % IN_WIDTH] : pong_storage_data_943 ^ i_input_data[1063 % IN_WIDTH];
                default: pong_storage_data_943 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_943;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_943 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_943;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_943 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_943;
            end
        end
    end
end

logic ping_storage_data_944;
logic pong_storage_data_944;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_944 <= 1'b0;
        pong_storage_data_944 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                562 / IN_WIDTH: ping_storage_data_944 <= (fillup_transition == 1'b1) ? i_input_data[562 % IN_WIDTH] : ping_storage_data_944 ^ i_input_data[562 % IN_WIDTH];
                693 / IN_WIDTH: ping_storage_data_944 <= (fillup_transition == 1'b1) ? i_input_data[693 % IN_WIDTH] : ping_storage_data_944 ^ i_input_data[693 % IN_WIDTH];
                970 / IN_WIDTH: ping_storage_data_944 <= (fillup_transition == 1'b1) ? i_input_data[970 % IN_WIDTH] : ping_storage_data_944 ^ i_input_data[970 % IN_WIDTH];
                1064 / IN_WIDTH: ping_storage_data_944 <= (fillup_transition == 1'b1) ? i_input_data[1064 % IN_WIDTH] : ping_storage_data_944 ^ i_input_data[1064 % IN_WIDTH];
                default: ping_storage_data_944 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_944;
                endcase
            end else begin
                case (input_count)
                562 / IN_WIDTH: pong_storage_data_944 <= (fillup_transition == 1'b1) ? i_input_data[562 % IN_WIDTH] : pong_storage_data_944 ^ i_input_data[562 % IN_WIDTH];
                693 / IN_WIDTH: pong_storage_data_944 <= (fillup_transition == 1'b1) ? i_input_data[693 % IN_WIDTH] : pong_storage_data_944 ^ i_input_data[693 % IN_WIDTH];
                970 / IN_WIDTH: pong_storage_data_944 <= (fillup_transition == 1'b1) ? i_input_data[970 % IN_WIDTH] : pong_storage_data_944 ^ i_input_data[970 % IN_WIDTH];
                1064 / IN_WIDTH: pong_storage_data_944 <= (fillup_transition == 1'b1) ? i_input_data[1064 % IN_WIDTH] : pong_storage_data_944 ^ i_input_data[1064 % IN_WIDTH];
                default: pong_storage_data_944 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_944;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_944 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_944;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_944 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_944;
            end
        end
    end
end

logic ping_storage_data_945;
logic pong_storage_data_945;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_945 <= 1'b0;
        pong_storage_data_945 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                563 / IN_WIDTH: ping_storage_data_945 <= (fillup_transition == 1'b1) ? i_input_data[563 % IN_WIDTH] : ping_storage_data_945 ^ i_input_data[563 % IN_WIDTH];
                694 / IN_WIDTH: ping_storage_data_945 <= (fillup_transition == 1'b1) ? i_input_data[694 % IN_WIDTH] : ping_storage_data_945 ^ i_input_data[694 % IN_WIDTH];
                971 / IN_WIDTH: ping_storage_data_945 <= (fillup_transition == 1'b1) ? i_input_data[971 % IN_WIDTH] : ping_storage_data_945 ^ i_input_data[971 % IN_WIDTH];
                1065 / IN_WIDTH: ping_storage_data_945 <= (fillup_transition == 1'b1) ? i_input_data[1065 % IN_WIDTH] : ping_storage_data_945 ^ i_input_data[1065 % IN_WIDTH];
                default: ping_storage_data_945 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_945;
                endcase
            end else begin
                case (input_count)
                563 / IN_WIDTH: pong_storage_data_945 <= (fillup_transition == 1'b1) ? i_input_data[563 % IN_WIDTH] : pong_storage_data_945 ^ i_input_data[563 % IN_WIDTH];
                694 / IN_WIDTH: pong_storage_data_945 <= (fillup_transition == 1'b1) ? i_input_data[694 % IN_WIDTH] : pong_storage_data_945 ^ i_input_data[694 % IN_WIDTH];
                971 / IN_WIDTH: pong_storage_data_945 <= (fillup_transition == 1'b1) ? i_input_data[971 % IN_WIDTH] : pong_storage_data_945 ^ i_input_data[971 % IN_WIDTH];
                1065 / IN_WIDTH: pong_storage_data_945 <= (fillup_transition == 1'b1) ? i_input_data[1065 % IN_WIDTH] : pong_storage_data_945 ^ i_input_data[1065 % IN_WIDTH];
                default: pong_storage_data_945 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_945;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_945 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_945;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_945 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_945;
            end
        end
    end
end

logic ping_storage_data_946;
logic pong_storage_data_946;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_946 <= 1'b0;
        pong_storage_data_946 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                564 / IN_WIDTH: ping_storage_data_946 <= (fillup_transition == 1'b1) ? i_input_data[564 % IN_WIDTH] : ping_storage_data_946 ^ i_input_data[564 % IN_WIDTH];
                695 / IN_WIDTH: ping_storage_data_946 <= (fillup_transition == 1'b1) ? i_input_data[695 % IN_WIDTH] : ping_storage_data_946 ^ i_input_data[695 % IN_WIDTH];
                972 / IN_WIDTH: ping_storage_data_946 <= (fillup_transition == 1'b1) ? i_input_data[972 % IN_WIDTH] : ping_storage_data_946 ^ i_input_data[972 % IN_WIDTH];
                1066 / IN_WIDTH: ping_storage_data_946 <= (fillup_transition == 1'b1) ? i_input_data[1066 % IN_WIDTH] : ping_storage_data_946 ^ i_input_data[1066 % IN_WIDTH];
                default: ping_storage_data_946 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_946;
                endcase
            end else begin
                case (input_count)
                564 / IN_WIDTH: pong_storage_data_946 <= (fillup_transition == 1'b1) ? i_input_data[564 % IN_WIDTH] : pong_storage_data_946 ^ i_input_data[564 % IN_WIDTH];
                695 / IN_WIDTH: pong_storage_data_946 <= (fillup_transition == 1'b1) ? i_input_data[695 % IN_WIDTH] : pong_storage_data_946 ^ i_input_data[695 % IN_WIDTH];
                972 / IN_WIDTH: pong_storage_data_946 <= (fillup_transition == 1'b1) ? i_input_data[972 % IN_WIDTH] : pong_storage_data_946 ^ i_input_data[972 % IN_WIDTH];
                1066 / IN_WIDTH: pong_storage_data_946 <= (fillup_transition == 1'b1) ? i_input_data[1066 % IN_WIDTH] : pong_storage_data_946 ^ i_input_data[1066 % IN_WIDTH];
                default: pong_storage_data_946 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_946;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_946 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_946;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_946 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_946;
            end
        end
    end
end

logic ping_storage_data_947;
logic pong_storage_data_947;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_947 <= 1'b0;
        pong_storage_data_947 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                565 / IN_WIDTH: ping_storage_data_947 <= (fillup_transition == 1'b1) ? i_input_data[565 % IN_WIDTH] : ping_storage_data_947 ^ i_input_data[565 % IN_WIDTH];
                696 / IN_WIDTH: ping_storage_data_947 <= (fillup_transition == 1'b1) ? i_input_data[696 % IN_WIDTH] : ping_storage_data_947 ^ i_input_data[696 % IN_WIDTH];
                973 / IN_WIDTH: ping_storage_data_947 <= (fillup_transition == 1'b1) ? i_input_data[973 % IN_WIDTH] : ping_storage_data_947 ^ i_input_data[973 % IN_WIDTH];
                1067 / IN_WIDTH: ping_storage_data_947 <= (fillup_transition == 1'b1) ? i_input_data[1067 % IN_WIDTH] : ping_storage_data_947 ^ i_input_data[1067 % IN_WIDTH];
                default: ping_storage_data_947 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_947;
                endcase
            end else begin
                case (input_count)
                565 / IN_WIDTH: pong_storage_data_947 <= (fillup_transition == 1'b1) ? i_input_data[565 % IN_WIDTH] : pong_storage_data_947 ^ i_input_data[565 % IN_WIDTH];
                696 / IN_WIDTH: pong_storage_data_947 <= (fillup_transition == 1'b1) ? i_input_data[696 % IN_WIDTH] : pong_storage_data_947 ^ i_input_data[696 % IN_WIDTH];
                973 / IN_WIDTH: pong_storage_data_947 <= (fillup_transition == 1'b1) ? i_input_data[973 % IN_WIDTH] : pong_storage_data_947 ^ i_input_data[973 % IN_WIDTH];
                1067 / IN_WIDTH: pong_storage_data_947 <= (fillup_transition == 1'b1) ? i_input_data[1067 % IN_WIDTH] : pong_storage_data_947 ^ i_input_data[1067 % IN_WIDTH];
                default: pong_storage_data_947 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_947;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_947 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_947;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_947 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_947;
            end
        end
    end
end

logic ping_storage_data_948;
logic pong_storage_data_948;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_948 <= 1'b0;
        pong_storage_data_948 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                566 / IN_WIDTH: ping_storage_data_948 <= (fillup_transition == 1'b1) ? i_input_data[566 % IN_WIDTH] : ping_storage_data_948 ^ i_input_data[566 % IN_WIDTH];
                697 / IN_WIDTH: ping_storage_data_948 <= (fillup_transition == 1'b1) ? i_input_data[697 % IN_WIDTH] : ping_storage_data_948 ^ i_input_data[697 % IN_WIDTH];
                974 / IN_WIDTH: ping_storage_data_948 <= (fillup_transition == 1'b1) ? i_input_data[974 % IN_WIDTH] : ping_storage_data_948 ^ i_input_data[974 % IN_WIDTH];
                1068 / IN_WIDTH: ping_storage_data_948 <= (fillup_transition == 1'b1) ? i_input_data[1068 % IN_WIDTH] : ping_storage_data_948 ^ i_input_data[1068 % IN_WIDTH];
                default: ping_storage_data_948 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_948;
                endcase
            end else begin
                case (input_count)
                566 / IN_WIDTH: pong_storage_data_948 <= (fillup_transition == 1'b1) ? i_input_data[566 % IN_WIDTH] : pong_storage_data_948 ^ i_input_data[566 % IN_WIDTH];
                697 / IN_WIDTH: pong_storage_data_948 <= (fillup_transition == 1'b1) ? i_input_data[697 % IN_WIDTH] : pong_storage_data_948 ^ i_input_data[697 % IN_WIDTH];
                974 / IN_WIDTH: pong_storage_data_948 <= (fillup_transition == 1'b1) ? i_input_data[974 % IN_WIDTH] : pong_storage_data_948 ^ i_input_data[974 % IN_WIDTH];
                1068 / IN_WIDTH: pong_storage_data_948 <= (fillup_transition == 1'b1) ? i_input_data[1068 % IN_WIDTH] : pong_storage_data_948 ^ i_input_data[1068 % IN_WIDTH];
                default: pong_storage_data_948 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_948;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_948 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_948;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_948 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_948;
            end
        end
    end
end

logic ping_storage_data_949;
logic pong_storage_data_949;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_949 <= 1'b0;
        pong_storage_data_949 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                567 / IN_WIDTH: ping_storage_data_949 <= (fillup_transition == 1'b1) ? i_input_data[567 % IN_WIDTH] : ping_storage_data_949 ^ i_input_data[567 % IN_WIDTH];
                698 / IN_WIDTH: ping_storage_data_949 <= (fillup_transition == 1'b1) ? i_input_data[698 % IN_WIDTH] : ping_storage_data_949 ^ i_input_data[698 % IN_WIDTH];
                975 / IN_WIDTH: ping_storage_data_949 <= (fillup_transition == 1'b1) ? i_input_data[975 % IN_WIDTH] : ping_storage_data_949 ^ i_input_data[975 % IN_WIDTH];
                1069 / IN_WIDTH: ping_storage_data_949 <= (fillup_transition == 1'b1) ? i_input_data[1069 % IN_WIDTH] : ping_storage_data_949 ^ i_input_data[1069 % IN_WIDTH];
                default: ping_storage_data_949 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_949;
                endcase
            end else begin
                case (input_count)
                567 / IN_WIDTH: pong_storage_data_949 <= (fillup_transition == 1'b1) ? i_input_data[567 % IN_WIDTH] : pong_storage_data_949 ^ i_input_data[567 % IN_WIDTH];
                698 / IN_WIDTH: pong_storage_data_949 <= (fillup_transition == 1'b1) ? i_input_data[698 % IN_WIDTH] : pong_storage_data_949 ^ i_input_data[698 % IN_WIDTH];
                975 / IN_WIDTH: pong_storage_data_949 <= (fillup_transition == 1'b1) ? i_input_data[975 % IN_WIDTH] : pong_storage_data_949 ^ i_input_data[975 % IN_WIDTH];
                1069 / IN_WIDTH: pong_storage_data_949 <= (fillup_transition == 1'b1) ? i_input_data[1069 % IN_WIDTH] : pong_storage_data_949 ^ i_input_data[1069 % IN_WIDTH];
                default: pong_storage_data_949 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_949;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_949 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_949;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_949 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_949;
            end
        end
    end
end

logic ping_storage_data_950;
logic pong_storage_data_950;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_950 <= 1'b0;
        pong_storage_data_950 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                568 / IN_WIDTH: ping_storage_data_950 <= (fillup_transition == 1'b1) ? i_input_data[568 % IN_WIDTH] : ping_storage_data_950 ^ i_input_data[568 % IN_WIDTH];
                699 / IN_WIDTH: ping_storage_data_950 <= (fillup_transition == 1'b1) ? i_input_data[699 % IN_WIDTH] : ping_storage_data_950 ^ i_input_data[699 % IN_WIDTH];
                976 / IN_WIDTH: ping_storage_data_950 <= (fillup_transition == 1'b1) ? i_input_data[976 % IN_WIDTH] : ping_storage_data_950 ^ i_input_data[976 % IN_WIDTH];
                1070 / IN_WIDTH: ping_storage_data_950 <= (fillup_transition == 1'b1) ? i_input_data[1070 % IN_WIDTH] : ping_storage_data_950 ^ i_input_data[1070 % IN_WIDTH];
                default: ping_storage_data_950 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_950;
                endcase
            end else begin
                case (input_count)
                568 / IN_WIDTH: pong_storage_data_950 <= (fillup_transition == 1'b1) ? i_input_data[568 % IN_WIDTH] : pong_storage_data_950 ^ i_input_data[568 % IN_WIDTH];
                699 / IN_WIDTH: pong_storage_data_950 <= (fillup_transition == 1'b1) ? i_input_data[699 % IN_WIDTH] : pong_storage_data_950 ^ i_input_data[699 % IN_WIDTH];
                976 / IN_WIDTH: pong_storage_data_950 <= (fillup_transition == 1'b1) ? i_input_data[976 % IN_WIDTH] : pong_storage_data_950 ^ i_input_data[976 % IN_WIDTH];
                1070 / IN_WIDTH: pong_storage_data_950 <= (fillup_transition == 1'b1) ? i_input_data[1070 % IN_WIDTH] : pong_storage_data_950 ^ i_input_data[1070 % IN_WIDTH];
                default: pong_storage_data_950 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_950;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_950 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_950;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_950 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_950;
            end
        end
    end
end

logic ping_storage_data_951;
logic pong_storage_data_951;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_951 <= 1'b0;
        pong_storage_data_951 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                569 / IN_WIDTH: ping_storage_data_951 <= (fillup_transition == 1'b1) ? i_input_data[569 % IN_WIDTH] : ping_storage_data_951 ^ i_input_data[569 % IN_WIDTH];
                700 / IN_WIDTH: ping_storage_data_951 <= (fillup_transition == 1'b1) ? i_input_data[700 % IN_WIDTH] : ping_storage_data_951 ^ i_input_data[700 % IN_WIDTH];
                977 / IN_WIDTH: ping_storage_data_951 <= (fillup_transition == 1'b1) ? i_input_data[977 % IN_WIDTH] : ping_storage_data_951 ^ i_input_data[977 % IN_WIDTH];
                1071 / IN_WIDTH: ping_storage_data_951 <= (fillup_transition == 1'b1) ? i_input_data[1071 % IN_WIDTH] : ping_storage_data_951 ^ i_input_data[1071 % IN_WIDTH];
                default: ping_storage_data_951 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_951;
                endcase
            end else begin
                case (input_count)
                569 / IN_WIDTH: pong_storage_data_951 <= (fillup_transition == 1'b1) ? i_input_data[569 % IN_WIDTH] : pong_storage_data_951 ^ i_input_data[569 % IN_WIDTH];
                700 / IN_WIDTH: pong_storage_data_951 <= (fillup_transition == 1'b1) ? i_input_data[700 % IN_WIDTH] : pong_storage_data_951 ^ i_input_data[700 % IN_WIDTH];
                977 / IN_WIDTH: pong_storage_data_951 <= (fillup_transition == 1'b1) ? i_input_data[977 % IN_WIDTH] : pong_storage_data_951 ^ i_input_data[977 % IN_WIDTH];
                1071 / IN_WIDTH: pong_storage_data_951 <= (fillup_transition == 1'b1) ? i_input_data[1071 % IN_WIDTH] : pong_storage_data_951 ^ i_input_data[1071 % IN_WIDTH];
                default: pong_storage_data_951 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_951;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_951 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_951;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_951 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_951;
            end
        end
    end
end

logic ping_storage_data_952;
logic pong_storage_data_952;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_952 <= 1'b0;
        pong_storage_data_952 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                570 / IN_WIDTH: ping_storage_data_952 <= (fillup_transition == 1'b1) ? i_input_data[570 % IN_WIDTH] : ping_storage_data_952 ^ i_input_data[570 % IN_WIDTH];
                701 / IN_WIDTH: ping_storage_data_952 <= (fillup_transition == 1'b1) ? i_input_data[701 % IN_WIDTH] : ping_storage_data_952 ^ i_input_data[701 % IN_WIDTH];
                978 / IN_WIDTH: ping_storage_data_952 <= (fillup_transition == 1'b1) ? i_input_data[978 % IN_WIDTH] : ping_storage_data_952 ^ i_input_data[978 % IN_WIDTH];
                1072 / IN_WIDTH: ping_storage_data_952 <= (fillup_transition == 1'b1) ? i_input_data[1072 % IN_WIDTH] : ping_storage_data_952 ^ i_input_data[1072 % IN_WIDTH];
                default: ping_storage_data_952 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_952;
                endcase
            end else begin
                case (input_count)
                570 / IN_WIDTH: pong_storage_data_952 <= (fillup_transition == 1'b1) ? i_input_data[570 % IN_WIDTH] : pong_storage_data_952 ^ i_input_data[570 % IN_WIDTH];
                701 / IN_WIDTH: pong_storage_data_952 <= (fillup_transition == 1'b1) ? i_input_data[701 % IN_WIDTH] : pong_storage_data_952 ^ i_input_data[701 % IN_WIDTH];
                978 / IN_WIDTH: pong_storage_data_952 <= (fillup_transition == 1'b1) ? i_input_data[978 % IN_WIDTH] : pong_storage_data_952 ^ i_input_data[978 % IN_WIDTH];
                1072 / IN_WIDTH: pong_storage_data_952 <= (fillup_transition == 1'b1) ? i_input_data[1072 % IN_WIDTH] : pong_storage_data_952 ^ i_input_data[1072 % IN_WIDTH];
                default: pong_storage_data_952 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_952;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_952 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_952;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_952 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_952;
            end
        end
    end
end

logic ping_storage_data_953;
logic pong_storage_data_953;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_953 <= 1'b0;
        pong_storage_data_953 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                571 / IN_WIDTH: ping_storage_data_953 <= (fillup_transition == 1'b1) ? i_input_data[571 % IN_WIDTH] : ping_storage_data_953 ^ i_input_data[571 % IN_WIDTH];
                702 / IN_WIDTH: ping_storage_data_953 <= (fillup_transition == 1'b1) ? i_input_data[702 % IN_WIDTH] : ping_storage_data_953 ^ i_input_data[702 % IN_WIDTH];
                979 / IN_WIDTH: ping_storage_data_953 <= (fillup_transition == 1'b1) ? i_input_data[979 % IN_WIDTH] : ping_storage_data_953 ^ i_input_data[979 % IN_WIDTH];
                1073 / IN_WIDTH: ping_storage_data_953 <= (fillup_transition == 1'b1) ? i_input_data[1073 % IN_WIDTH] : ping_storage_data_953 ^ i_input_data[1073 % IN_WIDTH];
                default: ping_storage_data_953 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_953;
                endcase
            end else begin
                case (input_count)
                571 / IN_WIDTH: pong_storage_data_953 <= (fillup_transition == 1'b1) ? i_input_data[571 % IN_WIDTH] : pong_storage_data_953 ^ i_input_data[571 % IN_WIDTH];
                702 / IN_WIDTH: pong_storage_data_953 <= (fillup_transition == 1'b1) ? i_input_data[702 % IN_WIDTH] : pong_storage_data_953 ^ i_input_data[702 % IN_WIDTH];
                979 / IN_WIDTH: pong_storage_data_953 <= (fillup_transition == 1'b1) ? i_input_data[979 % IN_WIDTH] : pong_storage_data_953 ^ i_input_data[979 % IN_WIDTH];
                1073 / IN_WIDTH: pong_storage_data_953 <= (fillup_transition == 1'b1) ? i_input_data[1073 % IN_WIDTH] : pong_storage_data_953 ^ i_input_data[1073 % IN_WIDTH];
                default: pong_storage_data_953 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_953;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_953 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_953;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_953 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_953;
            end
        end
    end
end

logic ping_storage_data_954;
logic pong_storage_data_954;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_954 <= 1'b0;
        pong_storage_data_954 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                572 / IN_WIDTH: ping_storage_data_954 <= (fillup_transition == 1'b1) ? i_input_data[572 % IN_WIDTH] : ping_storage_data_954 ^ i_input_data[572 % IN_WIDTH];
                703 / IN_WIDTH: ping_storage_data_954 <= (fillup_transition == 1'b1) ? i_input_data[703 % IN_WIDTH] : ping_storage_data_954 ^ i_input_data[703 % IN_WIDTH];
                980 / IN_WIDTH: ping_storage_data_954 <= (fillup_transition == 1'b1) ? i_input_data[980 % IN_WIDTH] : ping_storage_data_954 ^ i_input_data[980 % IN_WIDTH];
                1074 / IN_WIDTH: ping_storage_data_954 <= (fillup_transition == 1'b1) ? i_input_data[1074 % IN_WIDTH] : ping_storage_data_954 ^ i_input_data[1074 % IN_WIDTH];
                default: ping_storage_data_954 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_954;
                endcase
            end else begin
                case (input_count)
                572 / IN_WIDTH: pong_storage_data_954 <= (fillup_transition == 1'b1) ? i_input_data[572 % IN_WIDTH] : pong_storage_data_954 ^ i_input_data[572 % IN_WIDTH];
                703 / IN_WIDTH: pong_storage_data_954 <= (fillup_transition == 1'b1) ? i_input_data[703 % IN_WIDTH] : pong_storage_data_954 ^ i_input_data[703 % IN_WIDTH];
                980 / IN_WIDTH: pong_storage_data_954 <= (fillup_transition == 1'b1) ? i_input_data[980 % IN_WIDTH] : pong_storage_data_954 ^ i_input_data[980 % IN_WIDTH];
                1074 / IN_WIDTH: pong_storage_data_954 <= (fillup_transition == 1'b1) ? i_input_data[1074 % IN_WIDTH] : pong_storage_data_954 ^ i_input_data[1074 % IN_WIDTH];
                default: pong_storage_data_954 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_954;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_954 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_954;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_954 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_954;
            end
        end
    end
end

logic ping_storage_data_955;
logic pong_storage_data_955;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_955 <= 1'b0;
        pong_storage_data_955 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                573 / IN_WIDTH: ping_storage_data_955 <= (fillup_transition == 1'b1) ? i_input_data[573 % IN_WIDTH] : ping_storage_data_955 ^ i_input_data[573 % IN_WIDTH];
                704 / IN_WIDTH: ping_storage_data_955 <= (fillup_transition == 1'b1) ? i_input_data[704 % IN_WIDTH] : ping_storage_data_955 ^ i_input_data[704 % IN_WIDTH];
                981 / IN_WIDTH: ping_storage_data_955 <= (fillup_transition == 1'b1) ? i_input_data[981 % IN_WIDTH] : ping_storage_data_955 ^ i_input_data[981 % IN_WIDTH];
                1075 / IN_WIDTH: ping_storage_data_955 <= (fillup_transition == 1'b1) ? i_input_data[1075 % IN_WIDTH] : ping_storage_data_955 ^ i_input_data[1075 % IN_WIDTH];
                default: ping_storage_data_955 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_955;
                endcase
            end else begin
                case (input_count)
                573 / IN_WIDTH: pong_storage_data_955 <= (fillup_transition == 1'b1) ? i_input_data[573 % IN_WIDTH] : pong_storage_data_955 ^ i_input_data[573 % IN_WIDTH];
                704 / IN_WIDTH: pong_storage_data_955 <= (fillup_transition == 1'b1) ? i_input_data[704 % IN_WIDTH] : pong_storage_data_955 ^ i_input_data[704 % IN_WIDTH];
                981 / IN_WIDTH: pong_storage_data_955 <= (fillup_transition == 1'b1) ? i_input_data[981 % IN_WIDTH] : pong_storage_data_955 ^ i_input_data[981 % IN_WIDTH];
                1075 / IN_WIDTH: pong_storage_data_955 <= (fillup_transition == 1'b1) ? i_input_data[1075 % IN_WIDTH] : pong_storage_data_955 ^ i_input_data[1075 % IN_WIDTH];
                default: pong_storage_data_955 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_955;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_955 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_955;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_955 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_955;
            end
        end
    end
end

logic ping_storage_data_956;
logic pong_storage_data_956;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_956 <= 1'b0;
        pong_storage_data_956 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                574 / IN_WIDTH: ping_storage_data_956 <= (fillup_transition == 1'b1) ? i_input_data[574 % IN_WIDTH] : ping_storage_data_956 ^ i_input_data[574 % IN_WIDTH];
                705 / IN_WIDTH: ping_storage_data_956 <= (fillup_transition == 1'b1) ? i_input_data[705 % IN_WIDTH] : ping_storage_data_956 ^ i_input_data[705 % IN_WIDTH];
                982 / IN_WIDTH: ping_storage_data_956 <= (fillup_transition == 1'b1) ? i_input_data[982 % IN_WIDTH] : ping_storage_data_956 ^ i_input_data[982 % IN_WIDTH];
                1076 / IN_WIDTH: ping_storage_data_956 <= (fillup_transition == 1'b1) ? i_input_data[1076 % IN_WIDTH] : ping_storage_data_956 ^ i_input_data[1076 % IN_WIDTH];
                default: ping_storage_data_956 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_956;
                endcase
            end else begin
                case (input_count)
                574 / IN_WIDTH: pong_storage_data_956 <= (fillup_transition == 1'b1) ? i_input_data[574 % IN_WIDTH] : pong_storage_data_956 ^ i_input_data[574 % IN_WIDTH];
                705 / IN_WIDTH: pong_storage_data_956 <= (fillup_transition == 1'b1) ? i_input_data[705 % IN_WIDTH] : pong_storage_data_956 ^ i_input_data[705 % IN_WIDTH];
                982 / IN_WIDTH: pong_storage_data_956 <= (fillup_transition == 1'b1) ? i_input_data[982 % IN_WIDTH] : pong_storage_data_956 ^ i_input_data[982 % IN_WIDTH];
                1076 / IN_WIDTH: pong_storage_data_956 <= (fillup_transition == 1'b1) ? i_input_data[1076 % IN_WIDTH] : pong_storage_data_956 ^ i_input_data[1076 % IN_WIDTH];
                default: pong_storage_data_956 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_956;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_956 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_956;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_956 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_956;
            end
        end
    end
end

logic ping_storage_data_957;
logic pong_storage_data_957;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_957 <= 1'b0;
        pong_storage_data_957 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                575 / IN_WIDTH: ping_storage_data_957 <= (fillup_transition == 1'b1) ? i_input_data[575 % IN_WIDTH] : ping_storage_data_957 ^ i_input_data[575 % IN_WIDTH];
                706 / IN_WIDTH: ping_storage_data_957 <= (fillup_transition == 1'b1) ? i_input_data[706 % IN_WIDTH] : ping_storage_data_957 ^ i_input_data[706 % IN_WIDTH];
                983 / IN_WIDTH: ping_storage_data_957 <= (fillup_transition == 1'b1) ? i_input_data[983 % IN_WIDTH] : ping_storage_data_957 ^ i_input_data[983 % IN_WIDTH];
                1077 / IN_WIDTH: ping_storage_data_957 <= (fillup_transition == 1'b1) ? i_input_data[1077 % IN_WIDTH] : ping_storage_data_957 ^ i_input_data[1077 % IN_WIDTH];
                default: ping_storage_data_957 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_957;
                endcase
            end else begin
                case (input_count)
                575 / IN_WIDTH: pong_storage_data_957 <= (fillup_transition == 1'b1) ? i_input_data[575 % IN_WIDTH] : pong_storage_data_957 ^ i_input_data[575 % IN_WIDTH];
                706 / IN_WIDTH: pong_storage_data_957 <= (fillup_transition == 1'b1) ? i_input_data[706 % IN_WIDTH] : pong_storage_data_957 ^ i_input_data[706 % IN_WIDTH];
                983 / IN_WIDTH: pong_storage_data_957 <= (fillup_transition == 1'b1) ? i_input_data[983 % IN_WIDTH] : pong_storage_data_957 ^ i_input_data[983 % IN_WIDTH];
                1077 / IN_WIDTH: pong_storage_data_957 <= (fillup_transition == 1'b1) ? i_input_data[1077 % IN_WIDTH] : pong_storage_data_957 ^ i_input_data[1077 % IN_WIDTH];
                default: pong_storage_data_957 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_957;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_957 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_957;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_957 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_957;
            end
        end
    end
end

logic ping_storage_data_958;
logic pong_storage_data_958;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_958 <= 1'b0;
        pong_storage_data_958 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                480 / IN_WIDTH: ping_storage_data_958 <= (fillup_transition == 1'b1) ? i_input_data[480 % IN_WIDTH] : ping_storage_data_958 ^ i_input_data[480 % IN_WIDTH];
                707 / IN_WIDTH: ping_storage_data_958 <= (fillup_transition == 1'b1) ? i_input_data[707 % IN_WIDTH] : ping_storage_data_958 ^ i_input_data[707 % IN_WIDTH];
                984 / IN_WIDTH: ping_storage_data_958 <= (fillup_transition == 1'b1) ? i_input_data[984 % IN_WIDTH] : ping_storage_data_958 ^ i_input_data[984 % IN_WIDTH];
                1078 / IN_WIDTH: ping_storage_data_958 <= (fillup_transition == 1'b1) ? i_input_data[1078 % IN_WIDTH] : ping_storage_data_958 ^ i_input_data[1078 % IN_WIDTH];
                default: ping_storage_data_958 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_958;
                endcase
            end else begin
                case (input_count)
                480 / IN_WIDTH: pong_storage_data_958 <= (fillup_transition == 1'b1) ? i_input_data[480 % IN_WIDTH] : pong_storage_data_958 ^ i_input_data[480 % IN_WIDTH];
                707 / IN_WIDTH: pong_storage_data_958 <= (fillup_transition == 1'b1) ? i_input_data[707 % IN_WIDTH] : pong_storage_data_958 ^ i_input_data[707 % IN_WIDTH];
                984 / IN_WIDTH: pong_storage_data_958 <= (fillup_transition == 1'b1) ? i_input_data[984 % IN_WIDTH] : pong_storage_data_958 ^ i_input_data[984 % IN_WIDTH];
                1078 / IN_WIDTH: pong_storage_data_958 <= (fillup_transition == 1'b1) ? i_input_data[1078 % IN_WIDTH] : pong_storage_data_958 ^ i_input_data[1078 % IN_WIDTH];
                default: pong_storage_data_958 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_958;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_958 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_958;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_958 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_958;
            end
        end
    end
end

logic ping_storage_data_959;
logic pong_storage_data_959;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_959 <= 1'b0;
        pong_storage_data_959 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                481 / IN_WIDTH: ping_storage_data_959 <= (fillup_transition == 1'b1) ? i_input_data[481 % IN_WIDTH] : ping_storage_data_959 ^ i_input_data[481 % IN_WIDTH];
                708 / IN_WIDTH: ping_storage_data_959 <= (fillup_transition == 1'b1) ? i_input_data[708 % IN_WIDTH] : ping_storage_data_959 ^ i_input_data[708 % IN_WIDTH];
                985 / IN_WIDTH: ping_storage_data_959 <= (fillup_transition == 1'b1) ? i_input_data[985 % IN_WIDTH] : ping_storage_data_959 ^ i_input_data[985 % IN_WIDTH];
                1079 / IN_WIDTH: ping_storage_data_959 <= (fillup_transition == 1'b1) ? i_input_data[1079 % IN_WIDTH] : ping_storage_data_959 ^ i_input_data[1079 % IN_WIDTH];
                default: ping_storage_data_959 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_959;
                endcase
            end else begin
                case (input_count)
                481 / IN_WIDTH: pong_storage_data_959 <= (fillup_transition == 1'b1) ? i_input_data[481 % IN_WIDTH] : pong_storage_data_959 ^ i_input_data[481 % IN_WIDTH];
                708 / IN_WIDTH: pong_storage_data_959 <= (fillup_transition == 1'b1) ? i_input_data[708 % IN_WIDTH] : pong_storage_data_959 ^ i_input_data[708 % IN_WIDTH];
                985 / IN_WIDTH: pong_storage_data_959 <= (fillup_transition == 1'b1) ? i_input_data[985 % IN_WIDTH] : pong_storage_data_959 ^ i_input_data[985 % IN_WIDTH];
                1079 / IN_WIDTH: pong_storage_data_959 <= (fillup_transition == 1'b1) ? i_input_data[1079 % IN_WIDTH] : pong_storage_data_959 ^ i_input_data[1079 % IN_WIDTH];
                default: pong_storage_data_959 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_959;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_959 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_959;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_959 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_959;
            end
        end
    end
end

logic ping_storage_data_960;
logic pong_storage_data_960;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_960 <= 1'b0;
        pong_storage_data_960 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                281 / IN_WIDTH: ping_storage_data_960 <= (fillup_transition == 1'b1) ? i_input_data[281 % IN_WIDTH] : ping_storage_data_960 ^ i_input_data[281 % IN_WIDTH];
                319 / IN_WIDTH: ping_storage_data_960 <= (fillup_transition == 1'b1) ? i_input_data[319 % IN_WIDTH] : ping_storage_data_960 ^ i_input_data[319 % IN_WIDTH];
                825 / IN_WIDTH: ping_storage_data_960 <= (fillup_transition == 1'b1) ? i_input_data[825 % IN_WIDTH] : ping_storage_data_960 ^ i_input_data[825 % IN_WIDTH];
                911 / IN_WIDTH: ping_storage_data_960 <= (fillup_transition == 1'b1) ? i_input_data[911 % IN_WIDTH] : ping_storage_data_960 ^ i_input_data[911 % IN_WIDTH];
                default: ping_storage_data_960 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_960;
                endcase
            end else begin
                case (input_count)
                281 / IN_WIDTH: pong_storage_data_960 <= (fillup_transition == 1'b1) ? i_input_data[281 % IN_WIDTH] : pong_storage_data_960 ^ i_input_data[281 % IN_WIDTH];
                319 / IN_WIDTH: pong_storage_data_960 <= (fillup_transition == 1'b1) ? i_input_data[319 % IN_WIDTH] : pong_storage_data_960 ^ i_input_data[319 % IN_WIDTH];
                825 / IN_WIDTH: pong_storage_data_960 <= (fillup_transition == 1'b1) ? i_input_data[825 % IN_WIDTH] : pong_storage_data_960 ^ i_input_data[825 % IN_WIDTH];
                911 / IN_WIDTH: pong_storage_data_960 <= (fillup_transition == 1'b1) ? i_input_data[911 % IN_WIDTH] : pong_storage_data_960 ^ i_input_data[911 % IN_WIDTH];
                default: pong_storage_data_960 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_960;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_960 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_960;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_960 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_960;
            end
        end
    end
end

logic ping_storage_data_961;
logic pong_storage_data_961;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_961 <= 1'b0;
        pong_storage_data_961 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                282 / IN_WIDTH: ping_storage_data_961 <= (fillup_transition == 1'b1) ? i_input_data[282 % IN_WIDTH] : ping_storage_data_961 ^ i_input_data[282 % IN_WIDTH];
                320 / IN_WIDTH: ping_storage_data_961 <= (fillup_transition == 1'b1) ? i_input_data[320 % IN_WIDTH] : ping_storage_data_961 ^ i_input_data[320 % IN_WIDTH];
                826 / IN_WIDTH: ping_storage_data_961 <= (fillup_transition == 1'b1) ? i_input_data[826 % IN_WIDTH] : ping_storage_data_961 ^ i_input_data[826 % IN_WIDTH];
                912 / IN_WIDTH: ping_storage_data_961 <= (fillup_transition == 1'b1) ? i_input_data[912 % IN_WIDTH] : ping_storage_data_961 ^ i_input_data[912 % IN_WIDTH];
                default: ping_storage_data_961 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_961;
                endcase
            end else begin
                case (input_count)
                282 / IN_WIDTH: pong_storage_data_961 <= (fillup_transition == 1'b1) ? i_input_data[282 % IN_WIDTH] : pong_storage_data_961 ^ i_input_data[282 % IN_WIDTH];
                320 / IN_WIDTH: pong_storage_data_961 <= (fillup_transition == 1'b1) ? i_input_data[320 % IN_WIDTH] : pong_storage_data_961 ^ i_input_data[320 % IN_WIDTH];
                826 / IN_WIDTH: pong_storage_data_961 <= (fillup_transition == 1'b1) ? i_input_data[826 % IN_WIDTH] : pong_storage_data_961 ^ i_input_data[826 % IN_WIDTH];
                912 / IN_WIDTH: pong_storage_data_961 <= (fillup_transition == 1'b1) ? i_input_data[912 % IN_WIDTH] : pong_storage_data_961 ^ i_input_data[912 % IN_WIDTH];
                default: pong_storage_data_961 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_961;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_961 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_961;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_961 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_961;
            end
        end
    end
end

logic ping_storage_data_962;
logic pong_storage_data_962;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_962 <= 1'b0;
        pong_storage_data_962 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                283 / IN_WIDTH: ping_storage_data_962 <= (fillup_transition == 1'b1) ? i_input_data[283 % IN_WIDTH] : ping_storage_data_962 ^ i_input_data[283 % IN_WIDTH];
                321 / IN_WIDTH: ping_storage_data_962 <= (fillup_transition == 1'b1) ? i_input_data[321 % IN_WIDTH] : ping_storage_data_962 ^ i_input_data[321 % IN_WIDTH];
                827 / IN_WIDTH: ping_storage_data_962 <= (fillup_transition == 1'b1) ? i_input_data[827 % IN_WIDTH] : ping_storage_data_962 ^ i_input_data[827 % IN_WIDTH];
                913 / IN_WIDTH: ping_storage_data_962 <= (fillup_transition == 1'b1) ? i_input_data[913 % IN_WIDTH] : ping_storage_data_962 ^ i_input_data[913 % IN_WIDTH];
                default: ping_storage_data_962 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_962;
                endcase
            end else begin
                case (input_count)
                283 / IN_WIDTH: pong_storage_data_962 <= (fillup_transition == 1'b1) ? i_input_data[283 % IN_WIDTH] : pong_storage_data_962 ^ i_input_data[283 % IN_WIDTH];
                321 / IN_WIDTH: pong_storage_data_962 <= (fillup_transition == 1'b1) ? i_input_data[321 % IN_WIDTH] : pong_storage_data_962 ^ i_input_data[321 % IN_WIDTH];
                827 / IN_WIDTH: pong_storage_data_962 <= (fillup_transition == 1'b1) ? i_input_data[827 % IN_WIDTH] : pong_storage_data_962 ^ i_input_data[827 % IN_WIDTH];
                913 / IN_WIDTH: pong_storage_data_962 <= (fillup_transition == 1'b1) ? i_input_data[913 % IN_WIDTH] : pong_storage_data_962 ^ i_input_data[913 % IN_WIDTH];
                default: pong_storage_data_962 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_962;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_962 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_962;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_962 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_962;
            end
        end
    end
end

logic ping_storage_data_963;
logic pong_storage_data_963;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_963 <= 1'b0;
        pong_storage_data_963 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                284 / IN_WIDTH: ping_storage_data_963 <= (fillup_transition == 1'b1) ? i_input_data[284 % IN_WIDTH] : ping_storage_data_963 ^ i_input_data[284 % IN_WIDTH];
                322 / IN_WIDTH: ping_storage_data_963 <= (fillup_transition == 1'b1) ? i_input_data[322 % IN_WIDTH] : ping_storage_data_963 ^ i_input_data[322 % IN_WIDTH];
                828 / IN_WIDTH: ping_storage_data_963 <= (fillup_transition == 1'b1) ? i_input_data[828 % IN_WIDTH] : ping_storage_data_963 ^ i_input_data[828 % IN_WIDTH];
                914 / IN_WIDTH: ping_storage_data_963 <= (fillup_transition == 1'b1) ? i_input_data[914 % IN_WIDTH] : ping_storage_data_963 ^ i_input_data[914 % IN_WIDTH];
                default: ping_storage_data_963 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_963;
                endcase
            end else begin
                case (input_count)
                284 / IN_WIDTH: pong_storage_data_963 <= (fillup_transition == 1'b1) ? i_input_data[284 % IN_WIDTH] : pong_storage_data_963 ^ i_input_data[284 % IN_WIDTH];
                322 / IN_WIDTH: pong_storage_data_963 <= (fillup_transition == 1'b1) ? i_input_data[322 % IN_WIDTH] : pong_storage_data_963 ^ i_input_data[322 % IN_WIDTH];
                828 / IN_WIDTH: pong_storage_data_963 <= (fillup_transition == 1'b1) ? i_input_data[828 % IN_WIDTH] : pong_storage_data_963 ^ i_input_data[828 % IN_WIDTH];
                914 / IN_WIDTH: pong_storage_data_963 <= (fillup_transition == 1'b1) ? i_input_data[914 % IN_WIDTH] : pong_storage_data_963 ^ i_input_data[914 % IN_WIDTH];
                default: pong_storage_data_963 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_963;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_963 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_963;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_963 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_963;
            end
        end
    end
end

logic ping_storage_data_964;
logic pong_storage_data_964;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_964 <= 1'b0;
        pong_storage_data_964 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                285 / IN_WIDTH: ping_storage_data_964 <= (fillup_transition == 1'b1) ? i_input_data[285 % IN_WIDTH] : ping_storage_data_964 ^ i_input_data[285 % IN_WIDTH];
                323 / IN_WIDTH: ping_storage_data_964 <= (fillup_transition == 1'b1) ? i_input_data[323 % IN_WIDTH] : ping_storage_data_964 ^ i_input_data[323 % IN_WIDTH];
                829 / IN_WIDTH: ping_storage_data_964 <= (fillup_transition == 1'b1) ? i_input_data[829 % IN_WIDTH] : ping_storage_data_964 ^ i_input_data[829 % IN_WIDTH];
                915 / IN_WIDTH: ping_storage_data_964 <= (fillup_transition == 1'b1) ? i_input_data[915 % IN_WIDTH] : ping_storage_data_964 ^ i_input_data[915 % IN_WIDTH];
                default: ping_storage_data_964 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_964;
                endcase
            end else begin
                case (input_count)
                285 / IN_WIDTH: pong_storage_data_964 <= (fillup_transition == 1'b1) ? i_input_data[285 % IN_WIDTH] : pong_storage_data_964 ^ i_input_data[285 % IN_WIDTH];
                323 / IN_WIDTH: pong_storage_data_964 <= (fillup_transition == 1'b1) ? i_input_data[323 % IN_WIDTH] : pong_storage_data_964 ^ i_input_data[323 % IN_WIDTH];
                829 / IN_WIDTH: pong_storage_data_964 <= (fillup_transition == 1'b1) ? i_input_data[829 % IN_WIDTH] : pong_storage_data_964 ^ i_input_data[829 % IN_WIDTH];
                915 / IN_WIDTH: pong_storage_data_964 <= (fillup_transition == 1'b1) ? i_input_data[915 % IN_WIDTH] : pong_storage_data_964 ^ i_input_data[915 % IN_WIDTH];
                default: pong_storage_data_964 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_964;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_964 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_964;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_964 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_964;
            end
        end
    end
end

logic ping_storage_data_965;
logic pong_storage_data_965;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_965 <= 1'b0;
        pong_storage_data_965 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                286 / IN_WIDTH: ping_storage_data_965 <= (fillup_transition == 1'b1) ? i_input_data[286 % IN_WIDTH] : ping_storage_data_965 ^ i_input_data[286 % IN_WIDTH];
                324 / IN_WIDTH: ping_storage_data_965 <= (fillup_transition == 1'b1) ? i_input_data[324 % IN_WIDTH] : ping_storage_data_965 ^ i_input_data[324 % IN_WIDTH];
                830 / IN_WIDTH: ping_storage_data_965 <= (fillup_transition == 1'b1) ? i_input_data[830 % IN_WIDTH] : ping_storage_data_965 ^ i_input_data[830 % IN_WIDTH];
                916 / IN_WIDTH: ping_storage_data_965 <= (fillup_transition == 1'b1) ? i_input_data[916 % IN_WIDTH] : ping_storage_data_965 ^ i_input_data[916 % IN_WIDTH];
                default: ping_storage_data_965 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_965;
                endcase
            end else begin
                case (input_count)
                286 / IN_WIDTH: pong_storage_data_965 <= (fillup_transition == 1'b1) ? i_input_data[286 % IN_WIDTH] : pong_storage_data_965 ^ i_input_data[286 % IN_WIDTH];
                324 / IN_WIDTH: pong_storage_data_965 <= (fillup_transition == 1'b1) ? i_input_data[324 % IN_WIDTH] : pong_storage_data_965 ^ i_input_data[324 % IN_WIDTH];
                830 / IN_WIDTH: pong_storage_data_965 <= (fillup_transition == 1'b1) ? i_input_data[830 % IN_WIDTH] : pong_storage_data_965 ^ i_input_data[830 % IN_WIDTH];
                916 / IN_WIDTH: pong_storage_data_965 <= (fillup_transition == 1'b1) ? i_input_data[916 % IN_WIDTH] : pong_storage_data_965 ^ i_input_data[916 % IN_WIDTH];
                default: pong_storage_data_965 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_965;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_965 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_965;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_965 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_965;
            end
        end
    end
end

logic ping_storage_data_966;
logic pong_storage_data_966;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_966 <= 1'b0;
        pong_storage_data_966 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                287 / IN_WIDTH: ping_storage_data_966 <= (fillup_transition == 1'b1) ? i_input_data[287 % IN_WIDTH] : ping_storage_data_966 ^ i_input_data[287 % IN_WIDTH];
                325 / IN_WIDTH: ping_storage_data_966 <= (fillup_transition == 1'b1) ? i_input_data[325 % IN_WIDTH] : ping_storage_data_966 ^ i_input_data[325 % IN_WIDTH];
                831 / IN_WIDTH: ping_storage_data_966 <= (fillup_transition == 1'b1) ? i_input_data[831 % IN_WIDTH] : ping_storage_data_966 ^ i_input_data[831 % IN_WIDTH];
                917 / IN_WIDTH: ping_storage_data_966 <= (fillup_transition == 1'b1) ? i_input_data[917 % IN_WIDTH] : ping_storage_data_966 ^ i_input_data[917 % IN_WIDTH];
                default: ping_storage_data_966 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_966;
                endcase
            end else begin
                case (input_count)
                287 / IN_WIDTH: pong_storage_data_966 <= (fillup_transition == 1'b1) ? i_input_data[287 % IN_WIDTH] : pong_storage_data_966 ^ i_input_data[287 % IN_WIDTH];
                325 / IN_WIDTH: pong_storage_data_966 <= (fillup_transition == 1'b1) ? i_input_data[325 % IN_WIDTH] : pong_storage_data_966 ^ i_input_data[325 % IN_WIDTH];
                831 / IN_WIDTH: pong_storage_data_966 <= (fillup_transition == 1'b1) ? i_input_data[831 % IN_WIDTH] : pong_storage_data_966 ^ i_input_data[831 % IN_WIDTH];
                917 / IN_WIDTH: pong_storage_data_966 <= (fillup_transition == 1'b1) ? i_input_data[917 % IN_WIDTH] : pong_storage_data_966 ^ i_input_data[917 % IN_WIDTH];
                default: pong_storage_data_966 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_966;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_966 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_966;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_966 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_966;
            end
        end
    end
end

logic ping_storage_data_967;
logic pong_storage_data_967;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_967 <= 1'b0;
        pong_storage_data_967 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                192 / IN_WIDTH: ping_storage_data_967 <= (fillup_transition == 1'b1) ? i_input_data[192 % IN_WIDTH] : ping_storage_data_967 ^ i_input_data[192 % IN_WIDTH];
                326 / IN_WIDTH: ping_storage_data_967 <= (fillup_transition == 1'b1) ? i_input_data[326 % IN_WIDTH] : ping_storage_data_967 ^ i_input_data[326 % IN_WIDTH];
                832 / IN_WIDTH: ping_storage_data_967 <= (fillup_transition == 1'b1) ? i_input_data[832 % IN_WIDTH] : ping_storage_data_967 ^ i_input_data[832 % IN_WIDTH];
                918 / IN_WIDTH: ping_storage_data_967 <= (fillup_transition == 1'b1) ? i_input_data[918 % IN_WIDTH] : ping_storage_data_967 ^ i_input_data[918 % IN_WIDTH];
                default: ping_storage_data_967 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_967;
                endcase
            end else begin
                case (input_count)
                192 / IN_WIDTH: pong_storage_data_967 <= (fillup_transition == 1'b1) ? i_input_data[192 % IN_WIDTH] : pong_storage_data_967 ^ i_input_data[192 % IN_WIDTH];
                326 / IN_WIDTH: pong_storage_data_967 <= (fillup_transition == 1'b1) ? i_input_data[326 % IN_WIDTH] : pong_storage_data_967 ^ i_input_data[326 % IN_WIDTH];
                832 / IN_WIDTH: pong_storage_data_967 <= (fillup_transition == 1'b1) ? i_input_data[832 % IN_WIDTH] : pong_storage_data_967 ^ i_input_data[832 % IN_WIDTH];
                918 / IN_WIDTH: pong_storage_data_967 <= (fillup_transition == 1'b1) ? i_input_data[918 % IN_WIDTH] : pong_storage_data_967 ^ i_input_data[918 % IN_WIDTH];
                default: pong_storage_data_967 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_967;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_967 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_967;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_967 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_967;
            end
        end
    end
end

logic ping_storage_data_968;
logic pong_storage_data_968;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_968 <= 1'b0;
        pong_storage_data_968 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                193 / IN_WIDTH: ping_storage_data_968 <= (fillup_transition == 1'b1) ? i_input_data[193 % IN_WIDTH] : ping_storage_data_968 ^ i_input_data[193 % IN_WIDTH];
                327 / IN_WIDTH: ping_storage_data_968 <= (fillup_transition == 1'b1) ? i_input_data[327 % IN_WIDTH] : ping_storage_data_968 ^ i_input_data[327 % IN_WIDTH];
                833 / IN_WIDTH: ping_storage_data_968 <= (fillup_transition == 1'b1) ? i_input_data[833 % IN_WIDTH] : ping_storage_data_968 ^ i_input_data[833 % IN_WIDTH];
                919 / IN_WIDTH: ping_storage_data_968 <= (fillup_transition == 1'b1) ? i_input_data[919 % IN_WIDTH] : ping_storage_data_968 ^ i_input_data[919 % IN_WIDTH];
                default: ping_storage_data_968 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_968;
                endcase
            end else begin
                case (input_count)
                193 / IN_WIDTH: pong_storage_data_968 <= (fillup_transition == 1'b1) ? i_input_data[193 % IN_WIDTH] : pong_storage_data_968 ^ i_input_data[193 % IN_WIDTH];
                327 / IN_WIDTH: pong_storage_data_968 <= (fillup_transition == 1'b1) ? i_input_data[327 % IN_WIDTH] : pong_storage_data_968 ^ i_input_data[327 % IN_WIDTH];
                833 / IN_WIDTH: pong_storage_data_968 <= (fillup_transition == 1'b1) ? i_input_data[833 % IN_WIDTH] : pong_storage_data_968 ^ i_input_data[833 % IN_WIDTH];
                919 / IN_WIDTH: pong_storage_data_968 <= (fillup_transition == 1'b1) ? i_input_data[919 % IN_WIDTH] : pong_storage_data_968 ^ i_input_data[919 % IN_WIDTH];
                default: pong_storage_data_968 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_968;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_968 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_968;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_968 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_968;
            end
        end
    end
end

logic ping_storage_data_969;
logic pong_storage_data_969;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_969 <= 1'b0;
        pong_storage_data_969 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                194 / IN_WIDTH: ping_storage_data_969 <= (fillup_transition == 1'b1) ? i_input_data[194 % IN_WIDTH] : ping_storage_data_969 ^ i_input_data[194 % IN_WIDTH];
                328 / IN_WIDTH: ping_storage_data_969 <= (fillup_transition == 1'b1) ? i_input_data[328 % IN_WIDTH] : ping_storage_data_969 ^ i_input_data[328 % IN_WIDTH];
                834 / IN_WIDTH: ping_storage_data_969 <= (fillup_transition == 1'b1) ? i_input_data[834 % IN_WIDTH] : ping_storage_data_969 ^ i_input_data[834 % IN_WIDTH];
                920 / IN_WIDTH: ping_storage_data_969 <= (fillup_transition == 1'b1) ? i_input_data[920 % IN_WIDTH] : ping_storage_data_969 ^ i_input_data[920 % IN_WIDTH];
                default: ping_storage_data_969 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_969;
                endcase
            end else begin
                case (input_count)
                194 / IN_WIDTH: pong_storage_data_969 <= (fillup_transition == 1'b1) ? i_input_data[194 % IN_WIDTH] : pong_storage_data_969 ^ i_input_data[194 % IN_WIDTH];
                328 / IN_WIDTH: pong_storage_data_969 <= (fillup_transition == 1'b1) ? i_input_data[328 % IN_WIDTH] : pong_storage_data_969 ^ i_input_data[328 % IN_WIDTH];
                834 / IN_WIDTH: pong_storage_data_969 <= (fillup_transition == 1'b1) ? i_input_data[834 % IN_WIDTH] : pong_storage_data_969 ^ i_input_data[834 % IN_WIDTH];
                920 / IN_WIDTH: pong_storage_data_969 <= (fillup_transition == 1'b1) ? i_input_data[920 % IN_WIDTH] : pong_storage_data_969 ^ i_input_data[920 % IN_WIDTH];
                default: pong_storage_data_969 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_969;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_969 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_969;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_969 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_969;
            end
        end
    end
end

logic ping_storage_data_970;
logic pong_storage_data_970;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_970 <= 1'b0;
        pong_storage_data_970 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                195 / IN_WIDTH: ping_storage_data_970 <= (fillup_transition == 1'b1) ? i_input_data[195 % IN_WIDTH] : ping_storage_data_970 ^ i_input_data[195 % IN_WIDTH];
                329 / IN_WIDTH: ping_storage_data_970 <= (fillup_transition == 1'b1) ? i_input_data[329 % IN_WIDTH] : ping_storage_data_970 ^ i_input_data[329 % IN_WIDTH];
                835 / IN_WIDTH: ping_storage_data_970 <= (fillup_transition == 1'b1) ? i_input_data[835 % IN_WIDTH] : ping_storage_data_970 ^ i_input_data[835 % IN_WIDTH];
                921 / IN_WIDTH: ping_storage_data_970 <= (fillup_transition == 1'b1) ? i_input_data[921 % IN_WIDTH] : ping_storage_data_970 ^ i_input_data[921 % IN_WIDTH];
                default: ping_storage_data_970 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_970;
                endcase
            end else begin
                case (input_count)
                195 / IN_WIDTH: pong_storage_data_970 <= (fillup_transition == 1'b1) ? i_input_data[195 % IN_WIDTH] : pong_storage_data_970 ^ i_input_data[195 % IN_WIDTH];
                329 / IN_WIDTH: pong_storage_data_970 <= (fillup_transition == 1'b1) ? i_input_data[329 % IN_WIDTH] : pong_storage_data_970 ^ i_input_data[329 % IN_WIDTH];
                835 / IN_WIDTH: pong_storage_data_970 <= (fillup_transition == 1'b1) ? i_input_data[835 % IN_WIDTH] : pong_storage_data_970 ^ i_input_data[835 % IN_WIDTH];
                921 / IN_WIDTH: pong_storage_data_970 <= (fillup_transition == 1'b1) ? i_input_data[921 % IN_WIDTH] : pong_storage_data_970 ^ i_input_data[921 % IN_WIDTH];
                default: pong_storage_data_970 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_970;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_970 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_970;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_970 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_970;
            end
        end
    end
end

logic ping_storage_data_971;
logic pong_storage_data_971;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_971 <= 1'b0;
        pong_storage_data_971 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                196 / IN_WIDTH: ping_storage_data_971 <= (fillup_transition == 1'b1) ? i_input_data[196 % IN_WIDTH] : ping_storage_data_971 ^ i_input_data[196 % IN_WIDTH];
                330 / IN_WIDTH: ping_storage_data_971 <= (fillup_transition == 1'b1) ? i_input_data[330 % IN_WIDTH] : ping_storage_data_971 ^ i_input_data[330 % IN_WIDTH];
                836 / IN_WIDTH: ping_storage_data_971 <= (fillup_transition == 1'b1) ? i_input_data[836 % IN_WIDTH] : ping_storage_data_971 ^ i_input_data[836 % IN_WIDTH];
                922 / IN_WIDTH: ping_storage_data_971 <= (fillup_transition == 1'b1) ? i_input_data[922 % IN_WIDTH] : ping_storage_data_971 ^ i_input_data[922 % IN_WIDTH];
                default: ping_storage_data_971 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_971;
                endcase
            end else begin
                case (input_count)
                196 / IN_WIDTH: pong_storage_data_971 <= (fillup_transition == 1'b1) ? i_input_data[196 % IN_WIDTH] : pong_storage_data_971 ^ i_input_data[196 % IN_WIDTH];
                330 / IN_WIDTH: pong_storage_data_971 <= (fillup_transition == 1'b1) ? i_input_data[330 % IN_WIDTH] : pong_storage_data_971 ^ i_input_data[330 % IN_WIDTH];
                836 / IN_WIDTH: pong_storage_data_971 <= (fillup_transition == 1'b1) ? i_input_data[836 % IN_WIDTH] : pong_storage_data_971 ^ i_input_data[836 % IN_WIDTH];
                922 / IN_WIDTH: pong_storage_data_971 <= (fillup_transition == 1'b1) ? i_input_data[922 % IN_WIDTH] : pong_storage_data_971 ^ i_input_data[922 % IN_WIDTH];
                default: pong_storage_data_971 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_971;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_971 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_971;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_971 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_971;
            end
        end
    end
end

logic ping_storage_data_972;
logic pong_storage_data_972;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_972 <= 1'b0;
        pong_storage_data_972 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                197 / IN_WIDTH: ping_storage_data_972 <= (fillup_transition == 1'b1) ? i_input_data[197 % IN_WIDTH] : ping_storage_data_972 ^ i_input_data[197 % IN_WIDTH];
                331 / IN_WIDTH: ping_storage_data_972 <= (fillup_transition == 1'b1) ? i_input_data[331 % IN_WIDTH] : ping_storage_data_972 ^ i_input_data[331 % IN_WIDTH];
                837 / IN_WIDTH: ping_storage_data_972 <= (fillup_transition == 1'b1) ? i_input_data[837 % IN_WIDTH] : ping_storage_data_972 ^ i_input_data[837 % IN_WIDTH];
                923 / IN_WIDTH: ping_storage_data_972 <= (fillup_transition == 1'b1) ? i_input_data[923 % IN_WIDTH] : ping_storage_data_972 ^ i_input_data[923 % IN_WIDTH];
                default: ping_storage_data_972 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_972;
                endcase
            end else begin
                case (input_count)
                197 / IN_WIDTH: pong_storage_data_972 <= (fillup_transition == 1'b1) ? i_input_data[197 % IN_WIDTH] : pong_storage_data_972 ^ i_input_data[197 % IN_WIDTH];
                331 / IN_WIDTH: pong_storage_data_972 <= (fillup_transition == 1'b1) ? i_input_data[331 % IN_WIDTH] : pong_storage_data_972 ^ i_input_data[331 % IN_WIDTH];
                837 / IN_WIDTH: pong_storage_data_972 <= (fillup_transition == 1'b1) ? i_input_data[837 % IN_WIDTH] : pong_storage_data_972 ^ i_input_data[837 % IN_WIDTH];
                923 / IN_WIDTH: pong_storage_data_972 <= (fillup_transition == 1'b1) ? i_input_data[923 % IN_WIDTH] : pong_storage_data_972 ^ i_input_data[923 % IN_WIDTH];
                default: pong_storage_data_972 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_972;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_972 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_972;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_972 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_972;
            end
        end
    end
end

logic ping_storage_data_973;
logic pong_storage_data_973;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_973 <= 1'b0;
        pong_storage_data_973 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                198 / IN_WIDTH: ping_storage_data_973 <= (fillup_transition == 1'b1) ? i_input_data[198 % IN_WIDTH] : ping_storage_data_973 ^ i_input_data[198 % IN_WIDTH];
                332 / IN_WIDTH: ping_storage_data_973 <= (fillup_transition == 1'b1) ? i_input_data[332 % IN_WIDTH] : ping_storage_data_973 ^ i_input_data[332 % IN_WIDTH];
                838 / IN_WIDTH: ping_storage_data_973 <= (fillup_transition == 1'b1) ? i_input_data[838 % IN_WIDTH] : ping_storage_data_973 ^ i_input_data[838 % IN_WIDTH];
                924 / IN_WIDTH: ping_storage_data_973 <= (fillup_transition == 1'b1) ? i_input_data[924 % IN_WIDTH] : ping_storage_data_973 ^ i_input_data[924 % IN_WIDTH];
                default: ping_storage_data_973 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_973;
                endcase
            end else begin
                case (input_count)
                198 / IN_WIDTH: pong_storage_data_973 <= (fillup_transition == 1'b1) ? i_input_data[198 % IN_WIDTH] : pong_storage_data_973 ^ i_input_data[198 % IN_WIDTH];
                332 / IN_WIDTH: pong_storage_data_973 <= (fillup_transition == 1'b1) ? i_input_data[332 % IN_WIDTH] : pong_storage_data_973 ^ i_input_data[332 % IN_WIDTH];
                838 / IN_WIDTH: pong_storage_data_973 <= (fillup_transition == 1'b1) ? i_input_data[838 % IN_WIDTH] : pong_storage_data_973 ^ i_input_data[838 % IN_WIDTH];
                924 / IN_WIDTH: pong_storage_data_973 <= (fillup_transition == 1'b1) ? i_input_data[924 % IN_WIDTH] : pong_storage_data_973 ^ i_input_data[924 % IN_WIDTH];
                default: pong_storage_data_973 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_973;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_973 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_973;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_973 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_973;
            end
        end
    end
end

logic ping_storage_data_974;
logic pong_storage_data_974;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_974 <= 1'b0;
        pong_storage_data_974 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                199 / IN_WIDTH: ping_storage_data_974 <= (fillup_transition == 1'b1) ? i_input_data[199 % IN_WIDTH] : ping_storage_data_974 ^ i_input_data[199 % IN_WIDTH];
                333 / IN_WIDTH: ping_storage_data_974 <= (fillup_transition == 1'b1) ? i_input_data[333 % IN_WIDTH] : ping_storage_data_974 ^ i_input_data[333 % IN_WIDTH];
                839 / IN_WIDTH: ping_storage_data_974 <= (fillup_transition == 1'b1) ? i_input_data[839 % IN_WIDTH] : ping_storage_data_974 ^ i_input_data[839 % IN_WIDTH];
                925 / IN_WIDTH: ping_storage_data_974 <= (fillup_transition == 1'b1) ? i_input_data[925 % IN_WIDTH] : ping_storage_data_974 ^ i_input_data[925 % IN_WIDTH];
                default: ping_storage_data_974 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_974;
                endcase
            end else begin
                case (input_count)
                199 / IN_WIDTH: pong_storage_data_974 <= (fillup_transition == 1'b1) ? i_input_data[199 % IN_WIDTH] : pong_storage_data_974 ^ i_input_data[199 % IN_WIDTH];
                333 / IN_WIDTH: pong_storage_data_974 <= (fillup_transition == 1'b1) ? i_input_data[333 % IN_WIDTH] : pong_storage_data_974 ^ i_input_data[333 % IN_WIDTH];
                839 / IN_WIDTH: pong_storage_data_974 <= (fillup_transition == 1'b1) ? i_input_data[839 % IN_WIDTH] : pong_storage_data_974 ^ i_input_data[839 % IN_WIDTH];
                925 / IN_WIDTH: pong_storage_data_974 <= (fillup_transition == 1'b1) ? i_input_data[925 % IN_WIDTH] : pong_storage_data_974 ^ i_input_data[925 % IN_WIDTH];
                default: pong_storage_data_974 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_974;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_974 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_974;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_974 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_974;
            end
        end
    end
end

logic ping_storage_data_975;
logic pong_storage_data_975;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_975 <= 1'b0;
        pong_storage_data_975 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                200 / IN_WIDTH: ping_storage_data_975 <= (fillup_transition == 1'b1) ? i_input_data[200 % IN_WIDTH] : ping_storage_data_975 ^ i_input_data[200 % IN_WIDTH];
                334 / IN_WIDTH: ping_storage_data_975 <= (fillup_transition == 1'b1) ? i_input_data[334 % IN_WIDTH] : ping_storage_data_975 ^ i_input_data[334 % IN_WIDTH];
                840 / IN_WIDTH: ping_storage_data_975 <= (fillup_transition == 1'b1) ? i_input_data[840 % IN_WIDTH] : ping_storage_data_975 ^ i_input_data[840 % IN_WIDTH];
                926 / IN_WIDTH: ping_storage_data_975 <= (fillup_transition == 1'b1) ? i_input_data[926 % IN_WIDTH] : ping_storage_data_975 ^ i_input_data[926 % IN_WIDTH];
                default: ping_storage_data_975 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_975;
                endcase
            end else begin
                case (input_count)
                200 / IN_WIDTH: pong_storage_data_975 <= (fillup_transition == 1'b1) ? i_input_data[200 % IN_WIDTH] : pong_storage_data_975 ^ i_input_data[200 % IN_WIDTH];
                334 / IN_WIDTH: pong_storage_data_975 <= (fillup_transition == 1'b1) ? i_input_data[334 % IN_WIDTH] : pong_storage_data_975 ^ i_input_data[334 % IN_WIDTH];
                840 / IN_WIDTH: pong_storage_data_975 <= (fillup_transition == 1'b1) ? i_input_data[840 % IN_WIDTH] : pong_storage_data_975 ^ i_input_data[840 % IN_WIDTH];
                926 / IN_WIDTH: pong_storage_data_975 <= (fillup_transition == 1'b1) ? i_input_data[926 % IN_WIDTH] : pong_storage_data_975 ^ i_input_data[926 % IN_WIDTH];
                default: pong_storage_data_975 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_975;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_975 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_975;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_975 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_975;
            end
        end
    end
end

logic ping_storage_data_976;
logic pong_storage_data_976;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_976 <= 1'b0;
        pong_storage_data_976 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                201 / IN_WIDTH: ping_storage_data_976 <= (fillup_transition == 1'b1) ? i_input_data[201 % IN_WIDTH] : ping_storage_data_976 ^ i_input_data[201 % IN_WIDTH];
                335 / IN_WIDTH: ping_storage_data_976 <= (fillup_transition == 1'b1) ? i_input_data[335 % IN_WIDTH] : ping_storage_data_976 ^ i_input_data[335 % IN_WIDTH];
                841 / IN_WIDTH: ping_storage_data_976 <= (fillup_transition == 1'b1) ? i_input_data[841 % IN_WIDTH] : ping_storage_data_976 ^ i_input_data[841 % IN_WIDTH];
                927 / IN_WIDTH: ping_storage_data_976 <= (fillup_transition == 1'b1) ? i_input_data[927 % IN_WIDTH] : ping_storage_data_976 ^ i_input_data[927 % IN_WIDTH];
                default: ping_storage_data_976 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_976;
                endcase
            end else begin
                case (input_count)
                201 / IN_WIDTH: pong_storage_data_976 <= (fillup_transition == 1'b1) ? i_input_data[201 % IN_WIDTH] : pong_storage_data_976 ^ i_input_data[201 % IN_WIDTH];
                335 / IN_WIDTH: pong_storage_data_976 <= (fillup_transition == 1'b1) ? i_input_data[335 % IN_WIDTH] : pong_storage_data_976 ^ i_input_data[335 % IN_WIDTH];
                841 / IN_WIDTH: pong_storage_data_976 <= (fillup_transition == 1'b1) ? i_input_data[841 % IN_WIDTH] : pong_storage_data_976 ^ i_input_data[841 % IN_WIDTH];
                927 / IN_WIDTH: pong_storage_data_976 <= (fillup_transition == 1'b1) ? i_input_data[927 % IN_WIDTH] : pong_storage_data_976 ^ i_input_data[927 % IN_WIDTH];
                default: pong_storage_data_976 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_976;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_976 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_976;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_976 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_976;
            end
        end
    end
end

logic ping_storage_data_977;
logic pong_storage_data_977;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_977 <= 1'b0;
        pong_storage_data_977 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                202 / IN_WIDTH: ping_storage_data_977 <= (fillup_transition == 1'b1) ? i_input_data[202 % IN_WIDTH] : ping_storage_data_977 ^ i_input_data[202 % IN_WIDTH];
                336 / IN_WIDTH: ping_storage_data_977 <= (fillup_transition == 1'b1) ? i_input_data[336 % IN_WIDTH] : ping_storage_data_977 ^ i_input_data[336 % IN_WIDTH];
                842 / IN_WIDTH: ping_storage_data_977 <= (fillup_transition == 1'b1) ? i_input_data[842 % IN_WIDTH] : ping_storage_data_977 ^ i_input_data[842 % IN_WIDTH];
                928 / IN_WIDTH: ping_storage_data_977 <= (fillup_transition == 1'b1) ? i_input_data[928 % IN_WIDTH] : ping_storage_data_977 ^ i_input_data[928 % IN_WIDTH];
                default: ping_storage_data_977 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_977;
                endcase
            end else begin
                case (input_count)
                202 / IN_WIDTH: pong_storage_data_977 <= (fillup_transition == 1'b1) ? i_input_data[202 % IN_WIDTH] : pong_storage_data_977 ^ i_input_data[202 % IN_WIDTH];
                336 / IN_WIDTH: pong_storage_data_977 <= (fillup_transition == 1'b1) ? i_input_data[336 % IN_WIDTH] : pong_storage_data_977 ^ i_input_data[336 % IN_WIDTH];
                842 / IN_WIDTH: pong_storage_data_977 <= (fillup_transition == 1'b1) ? i_input_data[842 % IN_WIDTH] : pong_storage_data_977 ^ i_input_data[842 % IN_WIDTH];
                928 / IN_WIDTH: pong_storage_data_977 <= (fillup_transition == 1'b1) ? i_input_data[928 % IN_WIDTH] : pong_storage_data_977 ^ i_input_data[928 % IN_WIDTH];
                default: pong_storage_data_977 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_977;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_977 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_977;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_977 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_977;
            end
        end
    end
end

logic ping_storage_data_978;
logic pong_storage_data_978;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_978 <= 1'b0;
        pong_storage_data_978 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                203 / IN_WIDTH: ping_storage_data_978 <= (fillup_transition == 1'b1) ? i_input_data[203 % IN_WIDTH] : ping_storage_data_978 ^ i_input_data[203 % IN_WIDTH];
                337 / IN_WIDTH: ping_storage_data_978 <= (fillup_transition == 1'b1) ? i_input_data[337 % IN_WIDTH] : ping_storage_data_978 ^ i_input_data[337 % IN_WIDTH];
                843 / IN_WIDTH: ping_storage_data_978 <= (fillup_transition == 1'b1) ? i_input_data[843 % IN_WIDTH] : ping_storage_data_978 ^ i_input_data[843 % IN_WIDTH];
                929 / IN_WIDTH: ping_storage_data_978 <= (fillup_transition == 1'b1) ? i_input_data[929 % IN_WIDTH] : ping_storage_data_978 ^ i_input_data[929 % IN_WIDTH];
                default: ping_storage_data_978 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_978;
                endcase
            end else begin
                case (input_count)
                203 / IN_WIDTH: pong_storage_data_978 <= (fillup_transition == 1'b1) ? i_input_data[203 % IN_WIDTH] : pong_storage_data_978 ^ i_input_data[203 % IN_WIDTH];
                337 / IN_WIDTH: pong_storage_data_978 <= (fillup_transition == 1'b1) ? i_input_data[337 % IN_WIDTH] : pong_storage_data_978 ^ i_input_data[337 % IN_WIDTH];
                843 / IN_WIDTH: pong_storage_data_978 <= (fillup_transition == 1'b1) ? i_input_data[843 % IN_WIDTH] : pong_storage_data_978 ^ i_input_data[843 % IN_WIDTH];
                929 / IN_WIDTH: pong_storage_data_978 <= (fillup_transition == 1'b1) ? i_input_data[929 % IN_WIDTH] : pong_storage_data_978 ^ i_input_data[929 % IN_WIDTH];
                default: pong_storage_data_978 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_978;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_978 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_978;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_978 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_978;
            end
        end
    end
end

logic ping_storage_data_979;
logic pong_storage_data_979;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_979 <= 1'b0;
        pong_storage_data_979 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                204 / IN_WIDTH: ping_storage_data_979 <= (fillup_transition == 1'b1) ? i_input_data[204 % IN_WIDTH] : ping_storage_data_979 ^ i_input_data[204 % IN_WIDTH];
                338 / IN_WIDTH: ping_storage_data_979 <= (fillup_transition == 1'b1) ? i_input_data[338 % IN_WIDTH] : ping_storage_data_979 ^ i_input_data[338 % IN_WIDTH];
                844 / IN_WIDTH: ping_storage_data_979 <= (fillup_transition == 1'b1) ? i_input_data[844 % IN_WIDTH] : ping_storage_data_979 ^ i_input_data[844 % IN_WIDTH];
                930 / IN_WIDTH: ping_storage_data_979 <= (fillup_transition == 1'b1) ? i_input_data[930 % IN_WIDTH] : ping_storage_data_979 ^ i_input_data[930 % IN_WIDTH];
                default: ping_storage_data_979 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_979;
                endcase
            end else begin
                case (input_count)
                204 / IN_WIDTH: pong_storage_data_979 <= (fillup_transition == 1'b1) ? i_input_data[204 % IN_WIDTH] : pong_storage_data_979 ^ i_input_data[204 % IN_WIDTH];
                338 / IN_WIDTH: pong_storage_data_979 <= (fillup_transition == 1'b1) ? i_input_data[338 % IN_WIDTH] : pong_storage_data_979 ^ i_input_data[338 % IN_WIDTH];
                844 / IN_WIDTH: pong_storage_data_979 <= (fillup_transition == 1'b1) ? i_input_data[844 % IN_WIDTH] : pong_storage_data_979 ^ i_input_data[844 % IN_WIDTH];
                930 / IN_WIDTH: pong_storage_data_979 <= (fillup_transition == 1'b1) ? i_input_data[930 % IN_WIDTH] : pong_storage_data_979 ^ i_input_data[930 % IN_WIDTH];
                default: pong_storage_data_979 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_979;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_979 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_979;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_979 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_979;
            end
        end
    end
end

logic ping_storage_data_980;
logic pong_storage_data_980;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_980 <= 1'b0;
        pong_storage_data_980 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                205 / IN_WIDTH: ping_storage_data_980 <= (fillup_transition == 1'b1) ? i_input_data[205 % IN_WIDTH] : ping_storage_data_980 ^ i_input_data[205 % IN_WIDTH];
                339 / IN_WIDTH: ping_storage_data_980 <= (fillup_transition == 1'b1) ? i_input_data[339 % IN_WIDTH] : ping_storage_data_980 ^ i_input_data[339 % IN_WIDTH];
                845 / IN_WIDTH: ping_storage_data_980 <= (fillup_transition == 1'b1) ? i_input_data[845 % IN_WIDTH] : ping_storage_data_980 ^ i_input_data[845 % IN_WIDTH];
                931 / IN_WIDTH: ping_storage_data_980 <= (fillup_transition == 1'b1) ? i_input_data[931 % IN_WIDTH] : ping_storage_data_980 ^ i_input_data[931 % IN_WIDTH];
                default: ping_storage_data_980 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_980;
                endcase
            end else begin
                case (input_count)
                205 / IN_WIDTH: pong_storage_data_980 <= (fillup_transition == 1'b1) ? i_input_data[205 % IN_WIDTH] : pong_storage_data_980 ^ i_input_data[205 % IN_WIDTH];
                339 / IN_WIDTH: pong_storage_data_980 <= (fillup_transition == 1'b1) ? i_input_data[339 % IN_WIDTH] : pong_storage_data_980 ^ i_input_data[339 % IN_WIDTH];
                845 / IN_WIDTH: pong_storage_data_980 <= (fillup_transition == 1'b1) ? i_input_data[845 % IN_WIDTH] : pong_storage_data_980 ^ i_input_data[845 % IN_WIDTH];
                931 / IN_WIDTH: pong_storage_data_980 <= (fillup_transition == 1'b1) ? i_input_data[931 % IN_WIDTH] : pong_storage_data_980 ^ i_input_data[931 % IN_WIDTH];
                default: pong_storage_data_980 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_980;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_980 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_980;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_980 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_980;
            end
        end
    end
end

logic ping_storage_data_981;
logic pong_storage_data_981;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_981 <= 1'b0;
        pong_storage_data_981 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                206 / IN_WIDTH: ping_storage_data_981 <= (fillup_transition == 1'b1) ? i_input_data[206 % IN_WIDTH] : ping_storage_data_981 ^ i_input_data[206 % IN_WIDTH];
                340 / IN_WIDTH: ping_storage_data_981 <= (fillup_transition == 1'b1) ? i_input_data[340 % IN_WIDTH] : ping_storage_data_981 ^ i_input_data[340 % IN_WIDTH];
                846 / IN_WIDTH: ping_storage_data_981 <= (fillup_transition == 1'b1) ? i_input_data[846 % IN_WIDTH] : ping_storage_data_981 ^ i_input_data[846 % IN_WIDTH];
                932 / IN_WIDTH: ping_storage_data_981 <= (fillup_transition == 1'b1) ? i_input_data[932 % IN_WIDTH] : ping_storage_data_981 ^ i_input_data[932 % IN_WIDTH];
                default: ping_storage_data_981 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_981;
                endcase
            end else begin
                case (input_count)
                206 / IN_WIDTH: pong_storage_data_981 <= (fillup_transition == 1'b1) ? i_input_data[206 % IN_WIDTH] : pong_storage_data_981 ^ i_input_data[206 % IN_WIDTH];
                340 / IN_WIDTH: pong_storage_data_981 <= (fillup_transition == 1'b1) ? i_input_data[340 % IN_WIDTH] : pong_storage_data_981 ^ i_input_data[340 % IN_WIDTH];
                846 / IN_WIDTH: pong_storage_data_981 <= (fillup_transition == 1'b1) ? i_input_data[846 % IN_WIDTH] : pong_storage_data_981 ^ i_input_data[846 % IN_WIDTH];
                932 / IN_WIDTH: pong_storage_data_981 <= (fillup_transition == 1'b1) ? i_input_data[932 % IN_WIDTH] : pong_storage_data_981 ^ i_input_data[932 % IN_WIDTH];
                default: pong_storage_data_981 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_981;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_981 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_981;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_981 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_981;
            end
        end
    end
end

logic ping_storage_data_982;
logic pong_storage_data_982;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_982 <= 1'b0;
        pong_storage_data_982 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                207 / IN_WIDTH: ping_storage_data_982 <= (fillup_transition == 1'b1) ? i_input_data[207 % IN_WIDTH] : ping_storage_data_982 ^ i_input_data[207 % IN_WIDTH];
                341 / IN_WIDTH: ping_storage_data_982 <= (fillup_transition == 1'b1) ? i_input_data[341 % IN_WIDTH] : ping_storage_data_982 ^ i_input_data[341 % IN_WIDTH];
                847 / IN_WIDTH: ping_storage_data_982 <= (fillup_transition == 1'b1) ? i_input_data[847 % IN_WIDTH] : ping_storage_data_982 ^ i_input_data[847 % IN_WIDTH];
                933 / IN_WIDTH: ping_storage_data_982 <= (fillup_transition == 1'b1) ? i_input_data[933 % IN_WIDTH] : ping_storage_data_982 ^ i_input_data[933 % IN_WIDTH];
                default: ping_storage_data_982 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_982;
                endcase
            end else begin
                case (input_count)
                207 / IN_WIDTH: pong_storage_data_982 <= (fillup_transition == 1'b1) ? i_input_data[207 % IN_WIDTH] : pong_storage_data_982 ^ i_input_data[207 % IN_WIDTH];
                341 / IN_WIDTH: pong_storage_data_982 <= (fillup_transition == 1'b1) ? i_input_data[341 % IN_WIDTH] : pong_storage_data_982 ^ i_input_data[341 % IN_WIDTH];
                847 / IN_WIDTH: pong_storage_data_982 <= (fillup_transition == 1'b1) ? i_input_data[847 % IN_WIDTH] : pong_storage_data_982 ^ i_input_data[847 % IN_WIDTH];
                933 / IN_WIDTH: pong_storage_data_982 <= (fillup_transition == 1'b1) ? i_input_data[933 % IN_WIDTH] : pong_storage_data_982 ^ i_input_data[933 % IN_WIDTH];
                default: pong_storage_data_982 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_982;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_982 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_982;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_982 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_982;
            end
        end
    end
end

logic ping_storage_data_983;
logic pong_storage_data_983;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_983 <= 1'b0;
        pong_storage_data_983 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                208 / IN_WIDTH: ping_storage_data_983 <= (fillup_transition == 1'b1) ? i_input_data[208 % IN_WIDTH] : ping_storage_data_983 ^ i_input_data[208 % IN_WIDTH];
                342 / IN_WIDTH: ping_storage_data_983 <= (fillup_transition == 1'b1) ? i_input_data[342 % IN_WIDTH] : ping_storage_data_983 ^ i_input_data[342 % IN_WIDTH];
                848 / IN_WIDTH: ping_storage_data_983 <= (fillup_transition == 1'b1) ? i_input_data[848 % IN_WIDTH] : ping_storage_data_983 ^ i_input_data[848 % IN_WIDTH];
                934 / IN_WIDTH: ping_storage_data_983 <= (fillup_transition == 1'b1) ? i_input_data[934 % IN_WIDTH] : ping_storage_data_983 ^ i_input_data[934 % IN_WIDTH];
                default: ping_storage_data_983 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_983;
                endcase
            end else begin
                case (input_count)
                208 / IN_WIDTH: pong_storage_data_983 <= (fillup_transition == 1'b1) ? i_input_data[208 % IN_WIDTH] : pong_storage_data_983 ^ i_input_data[208 % IN_WIDTH];
                342 / IN_WIDTH: pong_storage_data_983 <= (fillup_transition == 1'b1) ? i_input_data[342 % IN_WIDTH] : pong_storage_data_983 ^ i_input_data[342 % IN_WIDTH];
                848 / IN_WIDTH: pong_storage_data_983 <= (fillup_transition == 1'b1) ? i_input_data[848 % IN_WIDTH] : pong_storage_data_983 ^ i_input_data[848 % IN_WIDTH];
                934 / IN_WIDTH: pong_storage_data_983 <= (fillup_transition == 1'b1) ? i_input_data[934 % IN_WIDTH] : pong_storage_data_983 ^ i_input_data[934 % IN_WIDTH];
                default: pong_storage_data_983 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_983;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_983 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_983;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_983 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_983;
            end
        end
    end
end

logic ping_storage_data_984;
logic pong_storage_data_984;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_984 <= 1'b0;
        pong_storage_data_984 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                209 / IN_WIDTH: ping_storage_data_984 <= (fillup_transition == 1'b1) ? i_input_data[209 % IN_WIDTH] : ping_storage_data_984 ^ i_input_data[209 % IN_WIDTH];
                343 / IN_WIDTH: ping_storage_data_984 <= (fillup_transition == 1'b1) ? i_input_data[343 % IN_WIDTH] : ping_storage_data_984 ^ i_input_data[343 % IN_WIDTH];
                849 / IN_WIDTH: ping_storage_data_984 <= (fillup_transition == 1'b1) ? i_input_data[849 % IN_WIDTH] : ping_storage_data_984 ^ i_input_data[849 % IN_WIDTH];
                935 / IN_WIDTH: ping_storage_data_984 <= (fillup_transition == 1'b1) ? i_input_data[935 % IN_WIDTH] : ping_storage_data_984 ^ i_input_data[935 % IN_WIDTH];
                default: ping_storage_data_984 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_984;
                endcase
            end else begin
                case (input_count)
                209 / IN_WIDTH: pong_storage_data_984 <= (fillup_transition == 1'b1) ? i_input_data[209 % IN_WIDTH] : pong_storage_data_984 ^ i_input_data[209 % IN_WIDTH];
                343 / IN_WIDTH: pong_storage_data_984 <= (fillup_transition == 1'b1) ? i_input_data[343 % IN_WIDTH] : pong_storage_data_984 ^ i_input_data[343 % IN_WIDTH];
                849 / IN_WIDTH: pong_storage_data_984 <= (fillup_transition == 1'b1) ? i_input_data[849 % IN_WIDTH] : pong_storage_data_984 ^ i_input_data[849 % IN_WIDTH];
                935 / IN_WIDTH: pong_storage_data_984 <= (fillup_transition == 1'b1) ? i_input_data[935 % IN_WIDTH] : pong_storage_data_984 ^ i_input_data[935 % IN_WIDTH];
                default: pong_storage_data_984 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_984;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_984 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_984;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_984 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_984;
            end
        end
    end
end

logic ping_storage_data_985;
logic pong_storage_data_985;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_985 <= 1'b0;
        pong_storage_data_985 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                210 / IN_WIDTH: ping_storage_data_985 <= (fillup_transition == 1'b1) ? i_input_data[210 % IN_WIDTH] : ping_storage_data_985 ^ i_input_data[210 % IN_WIDTH];
                344 / IN_WIDTH: ping_storage_data_985 <= (fillup_transition == 1'b1) ? i_input_data[344 % IN_WIDTH] : ping_storage_data_985 ^ i_input_data[344 % IN_WIDTH];
                850 / IN_WIDTH: ping_storage_data_985 <= (fillup_transition == 1'b1) ? i_input_data[850 % IN_WIDTH] : ping_storage_data_985 ^ i_input_data[850 % IN_WIDTH];
                936 / IN_WIDTH: ping_storage_data_985 <= (fillup_transition == 1'b1) ? i_input_data[936 % IN_WIDTH] : ping_storage_data_985 ^ i_input_data[936 % IN_WIDTH];
                default: ping_storage_data_985 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_985;
                endcase
            end else begin
                case (input_count)
                210 / IN_WIDTH: pong_storage_data_985 <= (fillup_transition == 1'b1) ? i_input_data[210 % IN_WIDTH] : pong_storage_data_985 ^ i_input_data[210 % IN_WIDTH];
                344 / IN_WIDTH: pong_storage_data_985 <= (fillup_transition == 1'b1) ? i_input_data[344 % IN_WIDTH] : pong_storage_data_985 ^ i_input_data[344 % IN_WIDTH];
                850 / IN_WIDTH: pong_storage_data_985 <= (fillup_transition == 1'b1) ? i_input_data[850 % IN_WIDTH] : pong_storage_data_985 ^ i_input_data[850 % IN_WIDTH];
                936 / IN_WIDTH: pong_storage_data_985 <= (fillup_transition == 1'b1) ? i_input_data[936 % IN_WIDTH] : pong_storage_data_985 ^ i_input_data[936 % IN_WIDTH];
                default: pong_storage_data_985 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_985;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_985 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_985;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_985 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_985;
            end
        end
    end
end

logic ping_storage_data_986;
logic pong_storage_data_986;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_986 <= 1'b0;
        pong_storage_data_986 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                211 / IN_WIDTH: ping_storage_data_986 <= (fillup_transition == 1'b1) ? i_input_data[211 % IN_WIDTH] : ping_storage_data_986 ^ i_input_data[211 % IN_WIDTH];
                345 / IN_WIDTH: ping_storage_data_986 <= (fillup_transition == 1'b1) ? i_input_data[345 % IN_WIDTH] : ping_storage_data_986 ^ i_input_data[345 % IN_WIDTH];
                851 / IN_WIDTH: ping_storage_data_986 <= (fillup_transition == 1'b1) ? i_input_data[851 % IN_WIDTH] : ping_storage_data_986 ^ i_input_data[851 % IN_WIDTH];
                937 / IN_WIDTH: ping_storage_data_986 <= (fillup_transition == 1'b1) ? i_input_data[937 % IN_WIDTH] : ping_storage_data_986 ^ i_input_data[937 % IN_WIDTH];
                default: ping_storage_data_986 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_986;
                endcase
            end else begin
                case (input_count)
                211 / IN_WIDTH: pong_storage_data_986 <= (fillup_transition == 1'b1) ? i_input_data[211 % IN_WIDTH] : pong_storage_data_986 ^ i_input_data[211 % IN_WIDTH];
                345 / IN_WIDTH: pong_storage_data_986 <= (fillup_transition == 1'b1) ? i_input_data[345 % IN_WIDTH] : pong_storage_data_986 ^ i_input_data[345 % IN_WIDTH];
                851 / IN_WIDTH: pong_storage_data_986 <= (fillup_transition == 1'b1) ? i_input_data[851 % IN_WIDTH] : pong_storage_data_986 ^ i_input_data[851 % IN_WIDTH];
                937 / IN_WIDTH: pong_storage_data_986 <= (fillup_transition == 1'b1) ? i_input_data[937 % IN_WIDTH] : pong_storage_data_986 ^ i_input_data[937 % IN_WIDTH];
                default: pong_storage_data_986 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_986;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_986 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_986;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_986 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_986;
            end
        end
    end
end

logic ping_storage_data_987;
logic pong_storage_data_987;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_987 <= 1'b0;
        pong_storage_data_987 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                212 / IN_WIDTH: ping_storage_data_987 <= (fillup_transition == 1'b1) ? i_input_data[212 % IN_WIDTH] : ping_storage_data_987 ^ i_input_data[212 % IN_WIDTH];
                346 / IN_WIDTH: ping_storage_data_987 <= (fillup_transition == 1'b1) ? i_input_data[346 % IN_WIDTH] : ping_storage_data_987 ^ i_input_data[346 % IN_WIDTH];
                852 / IN_WIDTH: ping_storage_data_987 <= (fillup_transition == 1'b1) ? i_input_data[852 % IN_WIDTH] : ping_storage_data_987 ^ i_input_data[852 % IN_WIDTH];
                938 / IN_WIDTH: ping_storage_data_987 <= (fillup_transition == 1'b1) ? i_input_data[938 % IN_WIDTH] : ping_storage_data_987 ^ i_input_data[938 % IN_WIDTH];
                default: ping_storage_data_987 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_987;
                endcase
            end else begin
                case (input_count)
                212 / IN_WIDTH: pong_storage_data_987 <= (fillup_transition == 1'b1) ? i_input_data[212 % IN_WIDTH] : pong_storage_data_987 ^ i_input_data[212 % IN_WIDTH];
                346 / IN_WIDTH: pong_storage_data_987 <= (fillup_transition == 1'b1) ? i_input_data[346 % IN_WIDTH] : pong_storage_data_987 ^ i_input_data[346 % IN_WIDTH];
                852 / IN_WIDTH: pong_storage_data_987 <= (fillup_transition == 1'b1) ? i_input_data[852 % IN_WIDTH] : pong_storage_data_987 ^ i_input_data[852 % IN_WIDTH];
                938 / IN_WIDTH: pong_storage_data_987 <= (fillup_transition == 1'b1) ? i_input_data[938 % IN_WIDTH] : pong_storage_data_987 ^ i_input_data[938 % IN_WIDTH];
                default: pong_storage_data_987 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_987;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_987 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_987;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_987 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_987;
            end
        end
    end
end

logic ping_storage_data_988;
logic pong_storage_data_988;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_988 <= 1'b0;
        pong_storage_data_988 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                213 / IN_WIDTH: ping_storage_data_988 <= (fillup_transition == 1'b1) ? i_input_data[213 % IN_WIDTH] : ping_storage_data_988 ^ i_input_data[213 % IN_WIDTH];
                347 / IN_WIDTH: ping_storage_data_988 <= (fillup_transition == 1'b1) ? i_input_data[347 % IN_WIDTH] : ping_storage_data_988 ^ i_input_data[347 % IN_WIDTH];
                853 / IN_WIDTH: ping_storage_data_988 <= (fillup_transition == 1'b1) ? i_input_data[853 % IN_WIDTH] : ping_storage_data_988 ^ i_input_data[853 % IN_WIDTH];
                939 / IN_WIDTH: ping_storage_data_988 <= (fillup_transition == 1'b1) ? i_input_data[939 % IN_WIDTH] : ping_storage_data_988 ^ i_input_data[939 % IN_WIDTH];
                default: ping_storage_data_988 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_988;
                endcase
            end else begin
                case (input_count)
                213 / IN_WIDTH: pong_storage_data_988 <= (fillup_transition == 1'b1) ? i_input_data[213 % IN_WIDTH] : pong_storage_data_988 ^ i_input_data[213 % IN_WIDTH];
                347 / IN_WIDTH: pong_storage_data_988 <= (fillup_transition == 1'b1) ? i_input_data[347 % IN_WIDTH] : pong_storage_data_988 ^ i_input_data[347 % IN_WIDTH];
                853 / IN_WIDTH: pong_storage_data_988 <= (fillup_transition == 1'b1) ? i_input_data[853 % IN_WIDTH] : pong_storage_data_988 ^ i_input_data[853 % IN_WIDTH];
                939 / IN_WIDTH: pong_storage_data_988 <= (fillup_transition == 1'b1) ? i_input_data[939 % IN_WIDTH] : pong_storage_data_988 ^ i_input_data[939 % IN_WIDTH];
                default: pong_storage_data_988 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_988;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_988 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_988;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_988 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_988;
            end
        end
    end
end

logic ping_storage_data_989;
logic pong_storage_data_989;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_989 <= 1'b0;
        pong_storage_data_989 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                214 / IN_WIDTH: ping_storage_data_989 <= (fillup_transition == 1'b1) ? i_input_data[214 % IN_WIDTH] : ping_storage_data_989 ^ i_input_data[214 % IN_WIDTH];
                348 / IN_WIDTH: ping_storage_data_989 <= (fillup_transition == 1'b1) ? i_input_data[348 % IN_WIDTH] : ping_storage_data_989 ^ i_input_data[348 % IN_WIDTH];
                854 / IN_WIDTH: ping_storage_data_989 <= (fillup_transition == 1'b1) ? i_input_data[854 % IN_WIDTH] : ping_storage_data_989 ^ i_input_data[854 % IN_WIDTH];
                940 / IN_WIDTH: ping_storage_data_989 <= (fillup_transition == 1'b1) ? i_input_data[940 % IN_WIDTH] : ping_storage_data_989 ^ i_input_data[940 % IN_WIDTH];
                default: ping_storage_data_989 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_989;
                endcase
            end else begin
                case (input_count)
                214 / IN_WIDTH: pong_storage_data_989 <= (fillup_transition == 1'b1) ? i_input_data[214 % IN_WIDTH] : pong_storage_data_989 ^ i_input_data[214 % IN_WIDTH];
                348 / IN_WIDTH: pong_storage_data_989 <= (fillup_transition == 1'b1) ? i_input_data[348 % IN_WIDTH] : pong_storage_data_989 ^ i_input_data[348 % IN_WIDTH];
                854 / IN_WIDTH: pong_storage_data_989 <= (fillup_transition == 1'b1) ? i_input_data[854 % IN_WIDTH] : pong_storage_data_989 ^ i_input_data[854 % IN_WIDTH];
                940 / IN_WIDTH: pong_storage_data_989 <= (fillup_transition == 1'b1) ? i_input_data[940 % IN_WIDTH] : pong_storage_data_989 ^ i_input_data[940 % IN_WIDTH];
                default: pong_storage_data_989 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_989;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_989 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_989;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_989 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_989;
            end
        end
    end
end

logic ping_storage_data_990;
logic pong_storage_data_990;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_990 <= 1'b0;
        pong_storage_data_990 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                215 / IN_WIDTH: ping_storage_data_990 <= (fillup_transition == 1'b1) ? i_input_data[215 % IN_WIDTH] : ping_storage_data_990 ^ i_input_data[215 % IN_WIDTH];
                349 / IN_WIDTH: ping_storage_data_990 <= (fillup_transition == 1'b1) ? i_input_data[349 % IN_WIDTH] : ping_storage_data_990 ^ i_input_data[349 % IN_WIDTH];
                855 / IN_WIDTH: ping_storage_data_990 <= (fillup_transition == 1'b1) ? i_input_data[855 % IN_WIDTH] : ping_storage_data_990 ^ i_input_data[855 % IN_WIDTH];
                941 / IN_WIDTH: ping_storage_data_990 <= (fillup_transition == 1'b1) ? i_input_data[941 % IN_WIDTH] : ping_storage_data_990 ^ i_input_data[941 % IN_WIDTH];
                default: ping_storage_data_990 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_990;
                endcase
            end else begin
                case (input_count)
                215 / IN_WIDTH: pong_storage_data_990 <= (fillup_transition == 1'b1) ? i_input_data[215 % IN_WIDTH] : pong_storage_data_990 ^ i_input_data[215 % IN_WIDTH];
                349 / IN_WIDTH: pong_storage_data_990 <= (fillup_transition == 1'b1) ? i_input_data[349 % IN_WIDTH] : pong_storage_data_990 ^ i_input_data[349 % IN_WIDTH];
                855 / IN_WIDTH: pong_storage_data_990 <= (fillup_transition == 1'b1) ? i_input_data[855 % IN_WIDTH] : pong_storage_data_990 ^ i_input_data[855 % IN_WIDTH];
                941 / IN_WIDTH: pong_storage_data_990 <= (fillup_transition == 1'b1) ? i_input_data[941 % IN_WIDTH] : pong_storage_data_990 ^ i_input_data[941 % IN_WIDTH];
                default: pong_storage_data_990 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_990;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_990 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_990;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_990 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_990;
            end
        end
    end
end

logic ping_storage_data_991;
logic pong_storage_data_991;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_991 <= 1'b0;
        pong_storage_data_991 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                216 / IN_WIDTH: ping_storage_data_991 <= (fillup_transition == 1'b1) ? i_input_data[216 % IN_WIDTH] : ping_storage_data_991 ^ i_input_data[216 % IN_WIDTH];
                350 / IN_WIDTH: ping_storage_data_991 <= (fillup_transition == 1'b1) ? i_input_data[350 % IN_WIDTH] : ping_storage_data_991 ^ i_input_data[350 % IN_WIDTH];
                856 / IN_WIDTH: ping_storage_data_991 <= (fillup_transition == 1'b1) ? i_input_data[856 % IN_WIDTH] : ping_storage_data_991 ^ i_input_data[856 % IN_WIDTH];
                942 / IN_WIDTH: ping_storage_data_991 <= (fillup_transition == 1'b1) ? i_input_data[942 % IN_WIDTH] : ping_storage_data_991 ^ i_input_data[942 % IN_WIDTH];
                default: ping_storage_data_991 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_991;
                endcase
            end else begin
                case (input_count)
                216 / IN_WIDTH: pong_storage_data_991 <= (fillup_transition == 1'b1) ? i_input_data[216 % IN_WIDTH] : pong_storage_data_991 ^ i_input_data[216 % IN_WIDTH];
                350 / IN_WIDTH: pong_storage_data_991 <= (fillup_transition == 1'b1) ? i_input_data[350 % IN_WIDTH] : pong_storage_data_991 ^ i_input_data[350 % IN_WIDTH];
                856 / IN_WIDTH: pong_storage_data_991 <= (fillup_transition == 1'b1) ? i_input_data[856 % IN_WIDTH] : pong_storage_data_991 ^ i_input_data[856 % IN_WIDTH];
                942 / IN_WIDTH: pong_storage_data_991 <= (fillup_transition == 1'b1) ? i_input_data[942 % IN_WIDTH] : pong_storage_data_991 ^ i_input_data[942 % IN_WIDTH];
                default: pong_storage_data_991 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_991;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_991 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_991;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_991 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_991;
            end
        end
    end
end

logic ping_storage_data_992;
logic pong_storage_data_992;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_992 <= 1'b0;
        pong_storage_data_992 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                217 / IN_WIDTH: ping_storage_data_992 <= (fillup_transition == 1'b1) ? i_input_data[217 % IN_WIDTH] : ping_storage_data_992 ^ i_input_data[217 % IN_WIDTH];
                351 / IN_WIDTH: ping_storage_data_992 <= (fillup_transition == 1'b1) ? i_input_data[351 % IN_WIDTH] : ping_storage_data_992 ^ i_input_data[351 % IN_WIDTH];
                857 / IN_WIDTH: ping_storage_data_992 <= (fillup_transition == 1'b1) ? i_input_data[857 % IN_WIDTH] : ping_storage_data_992 ^ i_input_data[857 % IN_WIDTH];
                943 / IN_WIDTH: ping_storage_data_992 <= (fillup_transition == 1'b1) ? i_input_data[943 % IN_WIDTH] : ping_storage_data_992 ^ i_input_data[943 % IN_WIDTH];
                default: ping_storage_data_992 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_992;
                endcase
            end else begin
                case (input_count)
                217 / IN_WIDTH: pong_storage_data_992 <= (fillup_transition == 1'b1) ? i_input_data[217 % IN_WIDTH] : pong_storage_data_992 ^ i_input_data[217 % IN_WIDTH];
                351 / IN_WIDTH: pong_storage_data_992 <= (fillup_transition == 1'b1) ? i_input_data[351 % IN_WIDTH] : pong_storage_data_992 ^ i_input_data[351 % IN_WIDTH];
                857 / IN_WIDTH: pong_storage_data_992 <= (fillup_transition == 1'b1) ? i_input_data[857 % IN_WIDTH] : pong_storage_data_992 ^ i_input_data[857 % IN_WIDTH];
                943 / IN_WIDTH: pong_storage_data_992 <= (fillup_transition == 1'b1) ? i_input_data[943 % IN_WIDTH] : pong_storage_data_992 ^ i_input_data[943 % IN_WIDTH];
                default: pong_storage_data_992 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_992;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_992 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_992;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_992 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_992;
            end
        end
    end
end

logic ping_storage_data_993;
logic pong_storage_data_993;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_993 <= 1'b0;
        pong_storage_data_993 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                218 / IN_WIDTH: ping_storage_data_993 <= (fillup_transition == 1'b1) ? i_input_data[218 % IN_WIDTH] : ping_storage_data_993 ^ i_input_data[218 % IN_WIDTH];
                352 / IN_WIDTH: ping_storage_data_993 <= (fillup_transition == 1'b1) ? i_input_data[352 % IN_WIDTH] : ping_storage_data_993 ^ i_input_data[352 % IN_WIDTH];
                858 / IN_WIDTH: ping_storage_data_993 <= (fillup_transition == 1'b1) ? i_input_data[858 % IN_WIDTH] : ping_storage_data_993 ^ i_input_data[858 % IN_WIDTH];
                944 / IN_WIDTH: ping_storage_data_993 <= (fillup_transition == 1'b1) ? i_input_data[944 % IN_WIDTH] : ping_storage_data_993 ^ i_input_data[944 % IN_WIDTH];
                default: ping_storage_data_993 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_993;
                endcase
            end else begin
                case (input_count)
                218 / IN_WIDTH: pong_storage_data_993 <= (fillup_transition == 1'b1) ? i_input_data[218 % IN_WIDTH] : pong_storage_data_993 ^ i_input_data[218 % IN_WIDTH];
                352 / IN_WIDTH: pong_storage_data_993 <= (fillup_transition == 1'b1) ? i_input_data[352 % IN_WIDTH] : pong_storage_data_993 ^ i_input_data[352 % IN_WIDTH];
                858 / IN_WIDTH: pong_storage_data_993 <= (fillup_transition == 1'b1) ? i_input_data[858 % IN_WIDTH] : pong_storage_data_993 ^ i_input_data[858 % IN_WIDTH];
                944 / IN_WIDTH: pong_storage_data_993 <= (fillup_transition == 1'b1) ? i_input_data[944 % IN_WIDTH] : pong_storage_data_993 ^ i_input_data[944 % IN_WIDTH];
                default: pong_storage_data_993 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_993;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_993 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_993;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_993 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_993;
            end
        end
    end
end

logic ping_storage_data_994;
logic pong_storage_data_994;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_994 <= 1'b0;
        pong_storage_data_994 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                219 / IN_WIDTH: ping_storage_data_994 <= (fillup_transition == 1'b1) ? i_input_data[219 % IN_WIDTH] : ping_storage_data_994 ^ i_input_data[219 % IN_WIDTH];
                353 / IN_WIDTH: ping_storage_data_994 <= (fillup_transition == 1'b1) ? i_input_data[353 % IN_WIDTH] : ping_storage_data_994 ^ i_input_data[353 % IN_WIDTH];
                859 / IN_WIDTH: ping_storage_data_994 <= (fillup_transition == 1'b1) ? i_input_data[859 % IN_WIDTH] : ping_storage_data_994 ^ i_input_data[859 % IN_WIDTH];
                945 / IN_WIDTH: ping_storage_data_994 <= (fillup_transition == 1'b1) ? i_input_data[945 % IN_WIDTH] : ping_storage_data_994 ^ i_input_data[945 % IN_WIDTH];
                default: ping_storage_data_994 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_994;
                endcase
            end else begin
                case (input_count)
                219 / IN_WIDTH: pong_storage_data_994 <= (fillup_transition == 1'b1) ? i_input_data[219 % IN_WIDTH] : pong_storage_data_994 ^ i_input_data[219 % IN_WIDTH];
                353 / IN_WIDTH: pong_storage_data_994 <= (fillup_transition == 1'b1) ? i_input_data[353 % IN_WIDTH] : pong_storage_data_994 ^ i_input_data[353 % IN_WIDTH];
                859 / IN_WIDTH: pong_storage_data_994 <= (fillup_transition == 1'b1) ? i_input_data[859 % IN_WIDTH] : pong_storage_data_994 ^ i_input_data[859 % IN_WIDTH];
                945 / IN_WIDTH: pong_storage_data_994 <= (fillup_transition == 1'b1) ? i_input_data[945 % IN_WIDTH] : pong_storage_data_994 ^ i_input_data[945 % IN_WIDTH];
                default: pong_storage_data_994 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_994;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_994 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_994;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_994 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_994;
            end
        end
    end
end

logic ping_storage_data_995;
logic pong_storage_data_995;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_995 <= 1'b0;
        pong_storage_data_995 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                220 / IN_WIDTH: ping_storage_data_995 <= (fillup_transition == 1'b1) ? i_input_data[220 % IN_WIDTH] : ping_storage_data_995 ^ i_input_data[220 % IN_WIDTH];
                354 / IN_WIDTH: ping_storage_data_995 <= (fillup_transition == 1'b1) ? i_input_data[354 % IN_WIDTH] : ping_storage_data_995 ^ i_input_data[354 % IN_WIDTH];
                860 / IN_WIDTH: ping_storage_data_995 <= (fillup_transition == 1'b1) ? i_input_data[860 % IN_WIDTH] : ping_storage_data_995 ^ i_input_data[860 % IN_WIDTH];
                946 / IN_WIDTH: ping_storage_data_995 <= (fillup_transition == 1'b1) ? i_input_data[946 % IN_WIDTH] : ping_storage_data_995 ^ i_input_data[946 % IN_WIDTH];
                default: ping_storage_data_995 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_995;
                endcase
            end else begin
                case (input_count)
                220 / IN_WIDTH: pong_storage_data_995 <= (fillup_transition == 1'b1) ? i_input_data[220 % IN_WIDTH] : pong_storage_data_995 ^ i_input_data[220 % IN_WIDTH];
                354 / IN_WIDTH: pong_storage_data_995 <= (fillup_transition == 1'b1) ? i_input_data[354 % IN_WIDTH] : pong_storage_data_995 ^ i_input_data[354 % IN_WIDTH];
                860 / IN_WIDTH: pong_storage_data_995 <= (fillup_transition == 1'b1) ? i_input_data[860 % IN_WIDTH] : pong_storage_data_995 ^ i_input_data[860 % IN_WIDTH];
                946 / IN_WIDTH: pong_storage_data_995 <= (fillup_transition == 1'b1) ? i_input_data[946 % IN_WIDTH] : pong_storage_data_995 ^ i_input_data[946 % IN_WIDTH];
                default: pong_storage_data_995 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_995;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_995 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_995;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_995 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_995;
            end
        end
    end
end

logic ping_storage_data_996;
logic pong_storage_data_996;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_996 <= 1'b0;
        pong_storage_data_996 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                221 / IN_WIDTH: ping_storage_data_996 <= (fillup_transition == 1'b1) ? i_input_data[221 % IN_WIDTH] : ping_storage_data_996 ^ i_input_data[221 % IN_WIDTH];
                355 / IN_WIDTH: ping_storage_data_996 <= (fillup_transition == 1'b1) ? i_input_data[355 % IN_WIDTH] : ping_storage_data_996 ^ i_input_data[355 % IN_WIDTH];
                861 / IN_WIDTH: ping_storage_data_996 <= (fillup_transition == 1'b1) ? i_input_data[861 % IN_WIDTH] : ping_storage_data_996 ^ i_input_data[861 % IN_WIDTH];
                947 / IN_WIDTH: ping_storage_data_996 <= (fillup_transition == 1'b1) ? i_input_data[947 % IN_WIDTH] : ping_storage_data_996 ^ i_input_data[947 % IN_WIDTH];
                default: ping_storage_data_996 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_996;
                endcase
            end else begin
                case (input_count)
                221 / IN_WIDTH: pong_storage_data_996 <= (fillup_transition == 1'b1) ? i_input_data[221 % IN_WIDTH] : pong_storage_data_996 ^ i_input_data[221 % IN_WIDTH];
                355 / IN_WIDTH: pong_storage_data_996 <= (fillup_transition == 1'b1) ? i_input_data[355 % IN_WIDTH] : pong_storage_data_996 ^ i_input_data[355 % IN_WIDTH];
                861 / IN_WIDTH: pong_storage_data_996 <= (fillup_transition == 1'b1) ? i_input_data[861 % IN_WIDTH] : pong_storage_data_996 ^ i_input_data[861 % IN_WIDTH];
                947 / IN_WIDTH: pong_storage_data_996 <= (fillup_transition == 1'b1) ? i_input_data[947 % IN_WIDTH] : pong_storage_data_996 ^ i_input_data[947 % IN_WIDTH];
                default: pong_storage_data_996 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_996;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_996 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_996;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_996 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_996;
            end
        end
    end
end

logic ping_storage_data_997;
logic pong_storage_data_997;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_997 <= 1'b0;
        pong_storage_data_997 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                222 / IN_WIDTH: ping_storage_data_997 <= (fillup_transition == 1'b1) ? i_input_data[222 % IN_WIDTH] : ping_storage_data_997 ^ i_input_data[222 % IN_WIDTH];
                356 / IN_WIDTH: ping_storage_data_997 <= (fillup_transition == 1'b1) ? i_input_data[356 % IN_WIDTH] : ping_storage_data_997 ^ i_input_data[356 % IN_WIDTH];
                862 / IN_WIDTH: ping_storage_data_997 <= (fillup_transition == 1'b1) ? i_input_data[862 % IN_WIDTH] : ping_storage_data_997 ^ i_input_data[862 % IN_WIDTH];
                948 / IN_WIDTH: ping_storage_data_997 <= (fillup_transition == 1'b1) ? i_input_data[948 % IN_WIDTH] : ping_storage_data_997 ^ i_input_data[948 % IN_WIDTH];
                default: ping_storage_data_997 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_997;
                endcase
            end else begin
                case (input_count)
                222 / IN_WIDTH: pong_storage_data_997 <= (fillup_transition == 1'b1) ? i_input_data[222 % IN_WIDTH] : pong_storage_data_997 ^ i_input_data[222 % IN_WIDTH];
                356 / IN_WIDTH: pong_storage_data_997 <= (fillup_transition == 1'b1) ? i_input_data[356 % IN_WIDTH] : pong_storage_data_997 ^ i_input_data[356 % IN_WIDTH];
                862 / IN_WIDTH: pong_storage_data_997 <= (fillup_transition == 1'b1) ? i_input_data[862 % IN_WIDTH] : pong_storage_data_997 ^ i_input_data[862 % IN_WIDTH];
                948 / IN_WIDTH: pong_storage_data_997 <= (fillup_transition == 1'b1) ? i_input_data[948 % IN_WIDTH] : pong_storage_data_997 ^ i_input_data[948 % IN_WIDTH];
                default: pong_storage_data_997 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_997;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_997 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_997;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_997 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_997;
            end
        end
    end
end

logic ping_storage_data_998;
logic pong_storage_data_998;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_998 <= 1'b0;
        pong_storage_data_998 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                223 / IN_WIDTH: ping_storage_data_998 <= (fillup_transition == 1'b1) ? i_input_data[223 % IN_WIDTH] : ping_storage_data_998 ^ i_input_data[223 % IN_WIDTH];
                357 / IN_WIDTH: ping_storage_data_998 <= (fillup_transition == 1'b1) ? i_input_data[357 % IN_WIDTH] : ping_storage_data_998 ^ i_input_data[357 % IN_WIDTH];
                863 / IN_WIDTH: ping_storage_data_998 <= (fillup_transition == 1'b1) ? i_input_data[863 % IN_WIDTH] : ping_storage_data_998 ^ i_input_data[863 % IN_WIDTH];
                949 / IN_WIDTH: ping_storage_data_998 <= (fillup_transition == 1'b1) ? i_input_data[949 % IN_WIDTH] : ping_storage_data_998 ^ i_input_data[949 % IN_WIDTH];
                default: ping_storage_data_998 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_998;
                endcase
            end else begin
                case (input_count)
                223 / IN_WIDTH: pong_storage_data_998 <= (fillup_transition == 1'b1) ? i_input_data[223 % IN_WIDTH] : pong_storage_data_998 ^ i_input_data[223 % IN_WIDTH];
                357 / IN_WIDTH: pong_storage_data_998 <= (fillup_transition == 1'b1) ? i_input_data[357 % IN_WIDTH] : pong_storage_data_998 ^ i_input_data[357 % IN_WIDTH];
                863 / IN_WIDTH: pong_storage_data_998 <= (fillup_transition == 1'b1) ? i_input_data[863 % IN_WIDTH] : pong_storage_data_998 ^ i_input_data[863 % IN_WIDTH];
                949 / IN_WIDTH: pong_storage_data_998 <= (fillup_transition == 1'b1) ? i_input_data[949 % IN_WIDTH] : pong_storage_data_998 ^ i_input_data[949 % IN_WIDTH];
                default: pong_storage_data_998 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_998;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_998 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_998;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_998 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_998;
            end
        end
    end
end

logic ping_storage_data_999;
logic pong_storage_data_999;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_999 <= 1'b0;
        pong_storage_data_999 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                224 / IN_WIDTH: ping_storage_data_999 <= (fillup_transition == 1'b1) ? i_input_data[224 % IN_WIDTH] : ping_storage_data_999 ^ i_input_data[224 % IN_WIDTH];
                358 / IN_WIDTH: ping_storage_data_999 <= (fillup_transition == 1'b1) ? i_input_data[358 % IN_WIDTH] : ping_storage_data_999 ^ i_input_data[358 % IN_WIDTH];
                768 / IN_WIDTH: ping_storage_data_999 <= (fillup_transition == 1'b1) ? i_input_data[768 % IN_WIDTH] : ping_storage_data_999 ^ i_input_data[768 % IN_WIDTH];
                950 / IN_WIDTH: ping_storage_data_999 <= (fillup_transition == 1'b1) ? i_input_data[950 % IN_WIDTH] : ping_storage_data_999 ^ i_input_data[950 % IN_WIDTH];
                default: ping_storage_data_999 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_999;
                endcase
            end else begin
                case (input_count)
                224 / IN_WIDTH: pong_storage_data_999 <= (fillup_transition == 1'b1) ? i_input_data[224 % IN_WIDTH] : pong_storage_data_999 ^ i_input_data[224 % IN_WIDTH];
                358 / IN_WIDTH: pong_storage_data_999 <= (fillup_transition == 1'b1) ? i_input_data[358 % IN_WIDTH] : pong_storage_data_999 ^ i_input_data[358 % IN_WIDTH];
                768 / IN_WIDTH: pong_storage_data_999 <= (fillup_transition == 1'b1) ? i_input_data[768 % IN_WIDTH] : pong_storage_data_999 ^ i_input_data[768 % IN_WIDTH];
                950 / IN_WIDTH: pong_storage_data_999 <= (fillup_transition == 1'b1) ? i_input_data[950 % IN_WIDTH] : pong_storage_data_999 ^ i_input_data[950 % IN_WIDTH];
                default: pong_storage_data_999 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_999;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_999 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_999;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_999 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_999;
            end
        end
    end
end

logic ping_storage_data_1000;
logic pong_storage_data_1000;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1000 <= 1'b0;
        pong_storage_data_1000 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                225 / IN_WIDTH: ping_storage_data_1000 <= (fillup_transition == 1'b1) ? i_input_data[225 % IN_WIDTH] : ping_storage_data_1000 ^ i_input_data[225 % IN_WIDTH];
                359 / IN_WIDTH: ping_storage_data_1000 <= (fillup_transition == 1'b1) ? i_input_data[359 % IN_WIDTH] : ping_storage_data_1000 ^ i_input_data[359 % IN_WIDTH];
                769 / IN_WIDTH: ping_storage_data_1000 <= (fillup_transition == 1'b1) ? i_input_data[769 % IN_WIDTH] : ping_storage_data_1000 ^ i_input_data[769 % IN_WIDTH];
                951 / IN_WIDTH: ping_storage_data_1000 <= (fillup_transition == 1'b1) ? i_input_data[951 % IN_WIDTH] : ping_storage_data_1000 ^ i_input_data[951 % IN_WIDTH];
                default: ping_storage_data_1000 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1000;
                endcase
            end else begin
                case (input_count)
                225 / IN_WIDTH: pong_storage_data_1000 <= (fillup_transition == 1'b1) ? i_input_data[225 % IN_WIDTH] : pong_storage_data_1000 ^ i_input_data[225 % IN_WIDTH];
                359 / IN_WIDTH: pong_storage_data_1000 <= (fillup_transition == 1'b1) ? i_input_data[359 % IN_WIDTH] : pong_storage_data_1000 ^ i_input_data[359 % IN_WIDTH];
                769 / IN_WIDTH: pong_storage_data_1000 <= (fillup_transition == 1'b1) ? i_input_data[769 % IN_WIDTH] : pong_storage_data_1000 ^ i_input_data[769 % IN_WIDTH];
                951 / IN_WIDTH: pong_storage_data_1000 <= (fillup_transition == 1'b1) ? i_input_data[951 % IN_WIDTH] : pong_storage_data_1000 ^ i_input_data[951 % IN_WIDTH];
                default: pong_storage_data_1000 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1000;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1000 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1000;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1000 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1000;
            end
        end
    end
end

logic ping_storage_data_1001;
logic pong_storage_data_1001;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1001 <= 1'b0;
        pong_storage_data_1001 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                226 / IN_WIDTH: ping_storage_data_1001 <= (fillup_transition == 1'b1) ? i_input_data[226 % IN_WIDTH] : ping_storage_data_1001 ^ i_input_data[226 % IN_WIDTH];
                360 / IN_WIDTH: ping_storage_data_1001 <= (fillup_transition == 1'b1) ? i_input_data[360 % IN_WIDTH] : ping_storage_data_1001 ^ i_input_data[360 % IN_WIDTH];
                770 / IN_WIDTH: ping_storage_data_1001 <= (fillup_transition == 1'b1) ? i_input_data[770 % IN_WIDTH] : ping_storage_data_1001 ^ i_input_data[770 % IN_WIDTH];
                952 / IN_WIDTH: ping_storage_data_1001 <= (fillup_transition == 1'b1) ? i_input_data[952 % IN_WIDTH] : ping_storage_data_1001 ^ i_input_data[952 % IN_WIDTH];
                default: ping_storage_data_1001 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1001;
                endcase
            end else begin
                case (input_count)
                226 / IN_WIDTH: pong_storage_data_1001 <= (fillup_transition == 1'b1) ? i_input_data[226 % IN_WIDTH] : pong_storage_data_1001 ^ i_input_data[226 % IN_WIDTH];
                360 / IN_WIDTH: pong_storage_data_1001 <= (fillup_transition == 1'b1) ? i_input_data[360 % IN_WIDTH] : pong_storage_data_1001 ^ i_input_data[360 % IN_WIDTH];
                770 / IN_WIDTH: pong_storage_data_1001 <= (fillup_transition == 1'b1) ? i_input_data[770 % IN_WIDTH] : pong_storage_data_1001 ^ i_input_data[770 % IN_WIDTH];
                952 / IN_WIDTH: pong_storage_data_1001 <= (fillup_transition == 1'b1) ? i_input_data[952 % IN_WIDTH] : pong_storage_data_1001 ^ i_input_data[952 % IN_WIDTH];
                default: pong_storage_data_1001 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1001;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1001 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1001;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1001 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1001;
            end
        end
    end
end

logic ping_storage_data_1002;
logic pong_storage_data_1002;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1002 <= 1'b0;
        pong_storage_data_1002 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                227 / IN_WIDTH: ping_storage_data_1002 <= (fillup_transition == 1'b1) ? i_input_data[227 % IN_WIDTH] : ping_storage_data_1002 ^ i_input_data[227 % IN_WIDTH];
                361 / IN_WIDTH: ping_storage_data_1002 <= (fillup_transition == 1'b1) ? i_input_data[361 % IN_WIDTH] : ping_storage_data_1002 ^ i_input_data[361 % IN_WIDTH];
                771 / IN_WIDTH: ping_storage_data_1002 <= (fillup_transition == 1'b1) ? i_input_data[771 % IN_WIDTH] : ping_storage_data_1002 ^ i_input_data[771 % IN_WIDTH];
                953 / IN_WIDTH: ping_storage_data_1002 <= (fillup_transition == 1'b1) ? i_input_data[953 % IN_WIDTH] : ping_storage_data_1002 ^ i_input_data[953 % IN_WIDTH];
                default: ping_storage_data_1002 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1002;
                endcase
            end else begin
                case (input_count)
                227 / IN_WIDTH: pong_storage_data_1002 <= (fillup_transition == 1'b1) ? i_input_data[227 % IN_WIDTH] : pong_storage_data_1002 ^ i_input_data[227 % IN_WIDTH];
                361 / IN_WIDTH: pong_storage_data_1002 <= (fillup_transition == 1'b1) ? i_input_data[361 % IN_WIDTH] : pong_storage_data_1002 ^ i_input_data[361 % IN_WIDTH];
                771 / IN_WIDTH: pong_storage_data_1002 <= (fillup_transition == 1'b1) ? i_input_data[771 % IN_WIDTH] : pong_storage_data_1002 ^ i_input_data[771 % IN_WIDTH];
                953 / IN_WIDTH: pong_storage_data_1002 <= (fillup_transition == 1'b1) ? i_input_data[953 % IN_WIDTH] : pong_storage_data_1002 ^ i_input_data[953 % IN_WIDTH];
                default: pong_storage_data_1002 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1002;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1002 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1002;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1002 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1002;
            end
        end
    end
end

logic ping_storage_data_1003;
logic pong_storage_data_1003;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1003 <= 1'b0;
        pong_storage_data_1003 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                228 / IN_WIDTH: ping_storage_data_1003 <= (fillup_transition == 1'b1) ? i_input_data[228 % IN_WIDTH] : ping_storage_data_1003 ^ i_input_data[228 % IN_WIDTH];
                362 / IN_WIDTH: ping_storage_data_1003 <= (fillup_transition == 1'b1) ? i_input_data[362 % IN_WIDTH] : ping_storage_data_1003 ^ i_input_data[362 % IN_WIDTH];
                772 / IN_WIDTH: ping_storage_data_1003 <= (fillup_transition == 1'b1) ? i_input_data[772 % IN_WIDTH] : ping_storage_data_1003 ^ i_input_data[772 % IN_WIDTH];
                954 / IN_WIDTH: ping_storage_data_1003 <= (fillup_transition == 1'b1) ? i_input_data[954 % IN_WIDTH] : ping_storage_data_1003 ^ i_input_data[954 % IN_WIDTH];
                default: ping_storage_data_1003 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1003;
                endcase
            end else begin
                case (input_count)
                228 / IN_WIDTH: pong_storage_data_1003 <= (fillup_transition == 1'b1) ? i_input_data[228 % IN_WIDTH] : pong_storage_data_1003 ^ i_input_data[228 % IN_WIDTH];
                362 / IN_WIDTH: pong_storage_data_1003 <= (fillup_transition == 1'b1) ? i_input_data[362 % IN_WIDTH] : pong_storage_data_1003 ^ i_input_data[362 % IN_WIDTH];
                772 / IN_WIDTH: pong_storage_data_1003 <= (fillup_transition == 1'b1) ? i_input_data[772 % IN_WIDTH] : pong_storage_data_1003 ^ i_input_data[772 % IN_WIDTH];
                954 / IN_WIDTH: pong_storage_data_1003 <= (fillup_transition == 1'b1) ? i_input_data[954 % IN_WIDTH] : pong_storage_data_1003 ^ i_input_data[954 % IN_WIDTH];
                default: pong_storage_data_1003 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1003;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1003 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1003;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1003 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1003;
            end
        end
    end
end

logic ping_storage_data_1004;
logic pong_storage_data_1004;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1004 <= 1'b0;
        pong_storage_data_1004 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                229 / IN_WIDTH: ping_storage_data_1004 <= (fillup_transition == 1'b1) ? i_input_data[229 % IN_WIDTH] : ping_storage_data_1004 ^ i_input_data[229 % IN_WIDTH];
                363 / IN_WIDTH: ping_storage_data_1004 <= (fillup_transition == 1'b1) ? i_input_data[363 % IN_WIDTH] : ping_storage_data_1004 ^ i_input_data[363 % IN_WIDTH];
                773 / IN_WIDTH: ping_storage_data_1004 <= (fillup_transition == 1'b1) ? i_input_data[773 % IN_WIDTH] : ping_storage_data_1004 ^ i_input_data[773 % IN_WIDTH];
                955 / IN_WIDTH: ping_storage_data_1004 <= (fillup_transition == 1'b1) ? i_input_data[955 % IN_WIDTH] : ping_storage_data_1004 ^ i_input_data[955 % IN_WIDTH];
                default: ping_storage_data_1004 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1004;
                endcase
            end else begin
                case (input_count)
                229 / IN_WIDTH: pong_storage_data_1004 <= (fillup_transition == 1'b1) ? i_input_data[229 % IN_WIDTH] : pong_storage_data_1004 ^ i_input_data[229 % IN_WIDTH];
                363 / IN_WIDTH: pong_storage_data_1004 <= (fillup_transition == 1'b1) ? i_input_data[363 % IN_WIDTH] : pong_storage_data_1004 ^ i_input_data[363 % IN_WIDTH];
                773 / IN_WIDTH: pong_storage_data_1004 <= (fillup_transition == 1'b1) ? i_input_data[773 % IN_WIDTH] : pong_storage_data_1004 ^ i_input_data[773 % IN_WIDTH];
                955 / IN_WIDTH: pong_storage_data_1004 <= (fillup_transition == 1'b1) ? i_input_data[955 % IN_WIDTH] : pong_storage_data_1004 ^ i_input_data[955 % IN_WIDTH];
                default: pong_storage_data_1004 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1004;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1004 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1004;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1004 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1004;
            end
        end
    end
end

logic ping_storage_data_1005;
logic pong_storage_data_1005;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1005 <= 1'b0;
        pong_storage_data_1005 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                230 / IN_WIDTH: ping_storage_data_1005 <= (fillup_transition == 1'b1) ? i_input_data[230 % IN_WIDTH] : ping_storage_data_1005 ^ i_input_data[230 % IN_WIDTH];
                364 / IN_WIDTH: ping_storage_data_1005 <= (fillup_transition == 1'b1) ? i_input_data[364 % IN_WIDTH] : ping_storage_data_1005 ^ i_input_data[364 % IN_WIDTH];
                774 / IN_WIDTH: ping_storage_data_1005 <= (fillup_transition == 1'b1) ? i_input_data[774 % IN_WIDTH] : ping_storage_data_1005 ^ i_input_data[774 % IN_WIDTH];
                956 / IN_WIDTH: ping_storage_data_1005 <= (fillup_transition == 1'b1) ? i_input_data[956 % IN_WIDTH] : ping_storage_data_1005 ^ i_input_data[956 % IN_WIDTH];
                default: ping_storage_data_1005 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1005;
                endcase
            end else begin
                case (input_count)
                230 / IN_WIDTH: pong_storage_data_1005 <= (fillup_transition == 1'b1) ? i_input_data[230 % IN_WIDTH] : pong_storage_data_1005 ^ i_input_data[230 % IN_WIDTH];
                364 / IN_WIDTH: pong_storage_data_1005 <= (fillup_transition == 1'b1) ? i_input_data[364 % IN_WIDTH] : pong_storage_data_1005 ^ i_input_data[364 % IN_WIDTH];
                774 / IN_WIDTH: pong_storage_data_1005 <= (fillup_transition == 1'b1) ? i_input_data[774 % IN_WIDTH] : pong_storage_data_1005 ^ i_input_data[774 % IN_WIDTH];
                956 / IN_WIDTH: pong_storage_data_1005 <= (fillup_transition == 1'b1) ? i_input_data[956 % IN_WIDTH] : pong_storage_data_1005 ^ i_input_data[956 % IN_WIDTH];
                default: pong_storage_data_1005 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1005;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1005 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1005;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1005 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1005;
            end
        end
    end
end

logic ping_storage_data_1006;
logic pong_storage_data_1006;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1006 <= 1'b0;
        pong_storage_data_1006 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                231 / IN_WIDTH: ping_storage_data_1006 <= (fillup_transition == 1'b1) ? i_input_data[231 % IN_WIDTH] : ping_storage_data_1006 ^ i_input_data[231 % IN_WIDTH];
                365 / IN_WIDTH: ping_storage_data_1006 <= (fillup_transition == 1'b1) ? i_input_data[365 % IN_WIDTH] : ping_storage_data_1006 ^ i_input_data[365 % IN_WIDTH];
                775 / IN_WIDTH: ping_storage_data_1006 <= (fillup_transition == 1'b1) ? i_input_data[775 % IN_WIDTH] : ping_storage_data_1006 ^ i_input_data[775 % IN_WIDTH];
                957 / IN_WIDTH: ping_storage_data_1006 <= (fillup_transition == 1'b1) ? i_input_data[957 % IN_WIDTH] : ping_storage_data_1006 ^ i_input_data[957 % IN_WIDTH];
                default: ping_storage_data_1006 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1006;
                endcase
            end else begin
                case (input_count)
                231 / IN_WIDTH: pong_storage_data_1006 <= (fillup_transition == 1'b1) ? i_input_data[231 % IN_WIDTH] : pong_storage_data_1006 ^ i_input_data[231 % IN_WIDTH];
                365 / IN_WIDTH: pong_storage_data_1006 <= (fillup_transition == 1'b1) ? i_input_data[365 % IN_WIDTH] : pong_storage_data_1006 ^ i_input_data[365 % IN_WIDTH];
                775 / IN_WIDTH: pong_storage_data_1006 <= (fillup_transition == 1'b1) ? i_input_data[775 % IN_WIDTH] : pong_storage_data_1006 ^ i_input_data[775 % IN_WIDTH];
                957 / IN_WIDTH: pong_storage_data_1006 <= (fillup_transition == 1'b1) ? i_input_data[957 % IN_WIDTH] : pong_storage_data_1006 ^ i_input_data[957 % IN_WIDTH];
                default: pong_storage_data_1006 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1006;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1006 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1006;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1006 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1006;
            end
        end
    end
end

logic ping_storage_data_1007;
logic pong_storage_data_1007;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1007 <= 1'b0;
        pong_storage_data_1007 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                232 / IN_WIDTH: ping_storage_data_1007 <= (fillup_transition == 1'b1) ? i_input_data[232 % IN_WIDTH] : ping_storage_data_1007 ^ i_input_data[232 % IN_WIDTH];
                366 / IN_WIDTH: ping_storage_data_1007 <= (fillup_transition == 1'b1) ? i_input_data[366 % IN_WIDTH] : ping_storage_data_1007 ^ i_input_data[366 % IN_WIDTH];
                776 / IN_WIDTH: ping_storage_data_1007 <= (fillup_transition == 1'b1) ? i_input_data[776 % IN_WIDTH] : ping_storage_data_1007 ^ i_input_data[776 % IN_WIDTH];
                958 / IN_WIDTH: ping_storage_data_1007 <= (fillup_transition == 1'b1) ? i_input_data[958 % IN_WIDTH] : ping_storage_data_1007 ^ i_input_data[958 % IN_WIDTH];
                default: ping_storage_data_1007 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1007;
                endcase
            end else begin
                case (input_count)
                232 / IN_WIDTH: pong_storage_data_1007 <= (fillup_transition == 1'b1) ? i_input_data[232 % IN_WIDTH] : pong_storage_data_1007 ^ i_input_data[232 % IN_WIDTH];
                366 / IN_WIDTH: pong_storage_data_1007 <= (fillup_transition == 1'b1) ? i_input_data[366 % IN_WIDTH] : pong_storage_data_1007 ^ i_input_data[366 % IN_WIDTH];
                776 / IN_WIDTH: pong_storage_data_1007 <= (fillup_transition == 1'b1) ? i_input_data[776 % IN_WIDTH] : pong_storage_data_1007 ^ i_input_data[776 % IN_WIDTH];
                958 / IN_WIDTH: pong_storage_data_1007 <= (fillup_transition == 1'b1) ? i_input_data[958 % IN_WIDTH] : pong_storage_data_1007 ^ i_input_data[958 % IN_WIDTH];
                default: pong_storage_data_1007 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1007;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1007 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1007;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1007 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1007;
            end
        end
    end
end

logic ping_storage_data_1008;
logic pong_storage_data_1008;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1008 <= 1'b0;
        pong_storage_data_1008 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                233 / IN_WIDTH: ping_storage_data_1008 <= (fillup_transition == 1'b1) ? i_input_data[233 % IN_WIDTH] : ping_storage_data_1008 ^ i_input_data[233 % IN_WIDTH];
                367 / IN_WIDTH: ping_storage_data_1008 <= (fillup_transition == 1'b1) ? i_input_data[367 % IN_WIDTH] : ping_storage_data_1008 ^ i_input_data[367 % IN_WIDTH];
                777 / IN_WIDTH: ping_storage_data_1008 <= (fillup_transition == 1'b1) ? i_input_data[777 % IN_WIDTH] : ping_storage_data_1008 ^ i_input_data[777 % IN_WIDTH];
                959 / IN_WIDTH: ping_storage_data_1008 <= (fillup_transition == 1'b1) ? i_input_data[959 % IN_WIDTH] : ping_storage_data_1008 ^ i_input_data[959 % IN_WIDTH];
                default: ping_storage_data_1008 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1008;
                endcase
            end else begin
                case (input_count)
                233 / IN_WIDTH: pong_storage_data_1008 <= (fillup_transition == 1'b1) ? i_input_data[233 % IN_WIDTH] : pong_storage_data_1008 ^ i_input_data[233 % IN_WIDTH];
                367 / IN_WIDTH: pong_storage_data_1008 <= (fillup_transition == 1'b1) ? i_input_data[367 % IN_WIDTH] : pong_storage_data_1008 ^ i_input_data[367 % IN_WIDTH];
                777 / IN_WIDTH: pong_storage_data_1008 <= (fillup_transition == 1'b1) ? i_input_data[777 % IN_WIDTH] : pong_storage_data_1008 ^ i_input_data[777 % IN_WIDTH];
                959 / IN_WIDTH: pong_storage_data_1008 <= (fillup_transition == 1'b1) ? i_input_data[959 % IN_WIDTH] : pong_storage_data_1008 ^ i_input_data[959 % IN_WIDTH];
                default: pong_storage_data_1008 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1008;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1008 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1008;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1008 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1008;
            end
        end
    end
end

logic ping_storage_data_1009;
logic pong_storage_data_1009;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1009 <= 1'b0;
        pong_storage_data_1009 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                234 / IN_WIDTH: ping_storage_data_1009 <= (fillup_transition == 1'b1) ? i_input_data[234 % IN_WIDTH] : ping_storage_data_1009 ^ i_input_data[234 % IN_WIDTH];
                368 / IN_WIDTH: ping_storage_data_1009 <= (fillup_transition == 1'b1) ? i_input_data[368 % IN_WIDTH] : ping_storage_data_1009 ^ i_input_data[368 % IN_WIDTH];
                778 / IN_WIDTH: ping_storage_data_1009 <= (fillup_transition == 1'b1) ? i_input_data[778 % IN_WIDTH] : ping_storage_data_1009 ^ i_input_data[778 % IN_WIDTH];
                864 / IN_WIDTH: ping_storage_data_1009 <= (fillup_transition == 1'b1) ? i_input_data[864 % IN_WIDTH] : ping_storage_data_1009 ^ i_input_data[864 % IN_WIDTH];
                default: ping_storage_data_1009 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1009;
                endcase
            end else begin
                case (input_count)
                234 / IN_WIDTH: pong_storage_data_1009 <= (fillup_transition == 1'b1) ? i_input_data[234 % IN_WIDTH] : pong_storage_data_1009 ^ i_input_data[234 % IN_WIDTH];
                368 / IN_WIDTH: pong_storage_data_1009 <= (fillup_transition == 1'b1) ? i_input_data[368 % IN_WIDTH] : pong_storage_data_1009 ^ i_input_data[368 % IN_WIDTH];
                778 / IN_WIDTH: pong_storage_data_1009 <= (fillup_transition == 1'b1) ? i_input_data[778 % IN_WIDTH] : pong_storage_data_1009 ^ i_input_data[778 % IN_WIDTH];
                864 / IN_WIDTH: pong_storage_data_1009 <= (fillup_transition == 1'b1) ? i_input_data[864 % IN_WIDTH] : pong_storage_data_1009 ^ i_input_data[864 % IN_WIDTH];
                default: pong_storage_data_1009 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1009;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1009 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1009;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1009 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1009;
            end
        end
    end
end

logic ping_storage_data_1010;
logic pong_storage_data_1010;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1010 <= 1'b0;
        pong_storage_data_1010 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                235 / IN_WIDTH: ping_storage_data_1010 <= (fillup_transition == 1'b1) ? i_input_data[235 % IN_WIDTH] : ping_storage_data_1010 ^ i_input_data[235 % IN_WIDTH];
                369 / IN_WIDTH: ping_storage_data_1010 <= (fillup_transition == 1'b1) ? i_input_data[369 % IN_WIDTH] : ping_storage_data_1010 ^ i_input_data[369 % IN_WIDTH];
                779 / IN_WIDTH: ping_storage_data_1010 <= (fillup_transition == 1'b1) ? i_input_data[779 % IN_WIDTH] : ping_storage_data_1010 ^ i_input_data[779 % IN_WIDTH];
                865 / IN_WIDTH: ping_storage_data_1010 <= (fillup_transition == 1'b1) ? i_input_data[865 % IN_WIDTH] : ping_storage_data_1010 ^ i_input_data[865 % IN_WIDTH];
                default: ping_storage_data_1010 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1010;
                endcase
            end else begin
                case (input_count)
                235 / IN_WIDTH: pong_storage_data_1010 <= (fillup_transition == 1'b1) ? i_input_data[235 % IN_WIDTH] : pong_storage_data_1010 ^ i_input_data[235 % IN_WIDTH];
                369 / IN_WIDTH: pong_storage_data_1010 <= (fillup_transition == 1'b1) ? i_input_data[369 % IN_WIDTH] : pong_storage_data_1010 ^ i_input_data[369 % IN_WIDTH];
                779 / IN_WIDTH: pong_storage_data_1010 <= (fillup_transition == 1'b1) ? i_input_data[779 % IN_WIDTH] : pong_storage_data_1010 ^ i_input_data[779 % IN_WIDTH];
                865 / IN_WIDTH: pong_storage_data_1010 <= (fillup_transition == 1'b1) ? i_input_data[865 % IN_WIDTH] : pong_storage_data_1010 ^ i_input_data[865 % IN_WIDTH];
                default: pong_storage_data_1010 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1010;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1010 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1010;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1010 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1010;
            end
        end
    end
end

logic ping_storage_data_1011;
logic pong_storage_data_1011;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1011 <= 1'b0;
        pong_storage_data_1011 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                236 / IN_WIDTH: ping_storage_data_1011 <= (fillup_transition == 1'b1) ? i_input_data[236 % IN_WIDTH] : ping_storage_data_1011 ^ i_input_data[236 % IN_WIDTH];
                370 / IN_WIDTH: ping_storage_data_1011 <= (fillup_transition == 1'b1) ? i_input_data[370 % IN_WIDTH] : ping_storage_data_1011 ^ i_input_data[370 % IN_WIDTH];
                780 / IN_WIDTH: ping_storage_data_1011 <= (fillup_transition == 1'b1) ? i_input_data[780 % IN_WIDTH] : ping_storage_data_1011 ^ i_input_data[780 % IN_WIDTH];
                866 / IN_WIDTH: ping_storage_data_1011 <= (fillup_transition == 1'b1) ? i_input_data[866 % IN_WIDTH] : ping_storage_data_1011 ^ i_input_data[866 % IN_WIDTH];
                default: ping_storage_data_1011 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1011;
                endcase
            end else begin
                case (input_count)
                236 / IN_WIDTH: pong_storage_data_1011 <= (fillup_transition == 1'b1) ? i_input_data[236 % IN_WIDTH] : pong_storage_data_1011 ^ i_input_data[236 % IN_WIDTH];
                370 / IN_WIDTH: pong_storage_data_1011 <= (fillup_transition == 1'b1) ? i_input_data[370 % IN_WIDTH] : pong_storage_data_1011 ^ i_input_data[370 % IN_WIDTH];
                780 / IN_WIDTH: pong_storage_data_1011 <= (fillup_transition == 1'b1) ? i_input_data[780 % IN_WIDTH] : pong_storage_data_1011 ^ i_input_data[780 % IN_WIDTH];
                866 / IN_WIDTH: pong_storage_data_1011 <= (fillup_transition == 1'b1) ? i_input_data[866 % IN_WIDTH] : pong_storage_data_1011 ^ i_input_data[866 % IN_WIDTH];
                default: pong_storage_data_1011 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1011;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1011 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1011;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1011 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1011;
            end
        end
    end
end

logic ping_storage_data_1012;
logic pong_storage_data_1012;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1012 <= 1'b0;
        pong_storage_data_1012 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                237 / IN_WIDTH: ping_storage_data_1012 <= (fillup_transition == 1'b1) ? i_input_data[237 % IN_WIDTH] : ping_storage_data_1012 ^ i_input_data[237 % IN_WIDTH];
                371 / IN_WIDTH: ping_storage_data_1012 <= (fillup_transition == 1'b1) ? i_input_data[371 % IN_WIDTH] : ping_storage_data_1012 ^ i_input_data[371 % IN_WIDTH];
                781 / IN_WIDTH: ping_storage_data_1012 <= (fillup_transition == 1'b1) ? i_input_data[781 % IN_WIDTH] : ping_storage_data_1012 ^ i_input_data[781 % IN_WIDTH];
                867 / IN_WIDTH: ping_storage_data_1012 <= (fillup_transition == 1'b1) ? i_input_data[867 % IN_WIDTH] : ping_storage_data_1012 ^ i_input_data[867 % IN_WIDTH];
                default: ping_storage_data_1012 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1012;
                endcase
            end else begin
                case (input_count)
                237 / IN_WIDTH: pong_storage_data_1012 <= (fillup_transition == 1'b1) ? i_input_data[237 % IN_WIDTH] : pong_storage_data_1012 ^ i_input_data[237 % IN_WIDTH];
                371 / IN_WIDTH: pong_storage_data_1012 <= (fillup_transition == 1'b1) ? i_input_data[371 % IN_WIDTH] : pong_storage_data_1012 ^ i_input_data[371 % IN_WIDTH];
                781 / IN_WIDTH: pong_storage_data_1012 <= (fillup_transition == 1'b1) ? i_input_data[781 % IN_WIDTH] : pong_storage_data_1012 ^ i_input_data[781 % IN_WIDTH];
                867 / IN_WIDTH: pong_storage_data_1012 <= (fillup_transition == 1'b1) ? i_input_data[867 % IN_WIDTH] : pong_storage_data_1012 ^ i_input_data[867 % IN_WIDTH];
                default: pong_storage_data_1012 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1012;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1012 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1012;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1012 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1012;
            end
        end
    end
end

logic ping_storage_data_1013;
logic pong_storage_data_1013;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1013 <= 1'b0;
        pong_storage_data_1013 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                238 / IN_WIDTH: ping_storage_data_1013 <= (fillup_transition == 1'b1) ? i_input_data[238 % IN_WIDTH] : ping_storage_data_1013 ^ i_input_data[238 % IN_WIDTH];
                372 / IN_WIDTH: ping_storage_data_1013 <= (fillup_transition == 1'b1) ? i_input_data[372 % IN_WIDTH] : ping_storage_data_1013 ^ i_input_data[372 % IN_WIDTH];
                782 / IN_WIDTH: ping_storage_data_1013 <= (fillup_transition == 1'b1) ? i_input_data[782 % IN_WIDTH] : ping_storage_data_1013 ^ i_input_data[782 % IN_WIDTH];
                868 / IN_WIDTH: ping_storage_data_1013 <= (fillup_transition == 1'b1) ? i_input_data[868 % IN_WIDTH] : ping_storage_data_1013 ^ i_input_data[868 % IN_WIDTH];
                default: ping_storage_data_1013 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1013;
                endcase
            end else begin
                case (input_count)
                238 / IN_WIDTH: pong_storage_data_1013 <= (fillup_transition == 1'b1) ? i_input_data[238 % IN_WIDTH] : pong_storage_data_1013 ^ i_input_data[238 % IN_WIDTH];
                372 / IN_WIDTH: pong_storage_data_1013 <= (fillup_transition == 1'b1) ? i_input_data[372 % IN_WIDTH] : pong_storage_data_1013 ^ i_input_data[372 % IN_WIDTH];
                782 / IN_WIDTH: pong_storage_data_1013 <= (fillup_transition == 1'b1) ? i_input_data[782 % IN_WIDTH] : pong_storage_data_1013 ^ i_input_data[782 % IN_WIDTH];
                868 / IN_WIDTH: pong_storage_data_1013 <= (fillup_transition == 1'b1) ? i_input_data[868 % IN_WIDTH] : pong_storage_data_1013 ^ i_input_data[868 % IN_WIDTH];
                default: pong_storage_data_1013 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1013;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1013 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1013;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1013 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1013;
            end
        end
    end
end

logic ping_storage_data_1014;
logic pong_storage_data_1014;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1014 <= 1'b0;
        pong_storage_data_1014 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                239 / IN_WIDTH: ping_storage_data_1014 <= (fillup_transition == 1'b1) ? i_input_data[239 % IN_WIDTH] : ping_storage_data_1014 ^ i_input_data[239 % IN_WIDTH];
                373 / IN_WIDTH: ping_storage_data_1014 <= (fillup_transition == 1'b1) ? i_input_data[373 % IN_WIDTH] : ping_storage_data_1014 ^ i_input_data[373 % IN_WIDTH];
                783 / IN_WIDTH: ping_storage_data_1014 <= (fillup_transition == 1'b1) ? i_input_data[783 % IN_WIDTH] : ping_storage_data_1014 ^ i_input_data[783 % IN_WIDTH];
                869 / IN_WIDTH: ping_storage_data_1014 <= (fillup_transition == 1'b1) ? i_input_data[869 % IN_WIDTH] : ping_storage_data_1014 ^ i_input_data[869 % IN_WIDTH];
                default: ping_storage_data_1014 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1014;
                endcase
            end else begin
                case (input_count)
                239 / IN_WIDTH: pong_storage_data_1014 <= (fillup_transition == 1'b1) ? i_input_data[239 % IN_WIDTH] : pong_storage_data_1014 ^ i_input_data[239 % IN_WIDTH];
                373 / IN_WIDTH: pong_storage_data_1014 <= (fillup_transition == 1'b1) ? i_input_data[373 % IN_WIDTH] : pong_storage_data_1014 ^ i_input_data[373 % IN_WIDTH];
                783 / IN_WIDTH: pong_storage_data_1014 <= (fillup_transition == 1'b1) ? i_input_data[783 % IN_WIDTH] : pong_storage_data_1014 ^ i_input_data[783 % IN_WIDTH];
                869 / IN_WIDTH: pong_storage_data_1014 <= (fillup_transition == 1'b1) ? i_input_data[869 % IN_WIDTH] : pong_storage_data_1014 ^ i_input_data[869 % IN_WIDTH];
                default: pong_storage_data_1014 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1014;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1014 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1014;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1014 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1014;
            end
        end
    end
end

logic ping_storage_data_1015;
logic pong_storage_data_1015;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1015 <= 1'b0;
        pong_storage_data_1015 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                240 / IN_WIDTH: ping_storage_data_1015 <= (fillup_transition == 1'b1) ? i_input_data[240 % IN_WIDTH] : ping_storage_data_1015 ^ i_input_data[240 % IN_WIDTH];
                374 / IN_WIDTH: ping_storage_data_1015 <= (fillup_transition == 1'b1) ? i_input_data[374 % IN_WIDTH] : ping_storage_data_1015 ^ i_input_data[374 % IN_WIDTH];
                784 / IN_WIDTH: ping_storage_data_1015 <= (fillup_transition == 1'b1) ? i_input_data[784 % IN_WIDTH] : ping_storage_data_1015 ^ i_input_data[784 % IN_WIDTH];
                870 / IN_WIDTH: ping_storage_data_1015 <= (fillup_transition == 1'b1) ? i_input_data[870 % IN_WIDTH] : ping_storage_data_1015 ^ i_input_data[870 % IN_WIDTH];
                default: ping_storage_data_1015 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1015;
                endcase
            end else begin
                case (input_count)
                240 / IN_WIDTH: pong_storage_data_1015 <= (fillup_transition == 1'b1) ? i_input_data[240 % IN_WIDTH] : pong_storage_data_1015 ^ i_input_data[240 % IN_WIDTH];
                374 / IN_WIDTH: pong_storage_data_1015 <= (fillup_transition == 1'b1) ? i_input_data[374 % IN_WIDTH] : pong_storage_data_1015 ^ i_input_data[374 % IN_WIDTH];
                784 / IN_WIDTH: pong_storage_data_1015 <= (fillup_transition == 1'b1) ? i_input_data[784 % IN_WIDTH] : pong_storage_data_1015 ^ i_input_data[784 % IN_WIDTH];
                870 / IN_WIDTH: pong_storage_data_1015 <= (fillup_transition == 1'b1) ? i_input_data[870 % IN_WIDTH] : pong_storage_data_1015 ^ i_input_data[870 % IN_WIDTH];
                default: pong_storage_data_1015 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1015;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1015 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1015;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1015 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1015;
            end
        end
    end
end

logic ping_storage_data_1016;
logic pong_storage_data_1016;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1016 <= 1'b0;
        pong_storage_data_1016 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                241 / IN_WIDTH: ping_storage_data_1016 <= (fillup_transition == 1'b1) ? i_input_data[241 % IN_WIDTH] : ping_storage_data_1016 ^ i_input_data[241 % IN_WIDTH];
                375 / IN_WIDTH: ping_storage_data_1016 <= (fillup_transition == 1'b1) ? i_input_data[375 % IN_WIDTH] : ping_storage_data_1016 ^ i_input_data[375 % IN_WIDTH];
                785 / IN_WIDTH: ping_storage_data_1016 <= (fillup_transition == 1'b1) ? i_input_data[785 % IN_WIDTH] : ping_storage_data_1016 ^ i_input_data[785 % IN_WIDTH];
                871 / IN_WIDTH: ping_storage_data_1016 <= (fillup_transition == 1'b1) ? i_input_data[871 % IN_WIDTH] : ping_storage_data_1016 ^ i_input_data[871 % IN_WIDTH];
                default: ping_storage_data_1016 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1016;
                endcase
            end else begin
                case (input_count)
                241 / IN_WIDTH: pong_storage_data_1016 <= (fillup_transition == 1'b1) ? i_input_data[241 % IN_WIDTH] : pong_storage_data_1016 ^ i_input_data[241 % IN_WIDTH];
                375 / IN_WIDTH: pong_storage_data_1016 <= (fillup_transition == 1'b1) ? i_input_data[375 % IN_WIDTH] : pong_storage_data_1016 ^ i_input_data[375 % IN_WIDTH];
                785 / IN_WIDTH: pong_storage_data_1016 <= (fillup_transition == 1'b1) ? i_input_data[785 % IN_WIDTH] : pong_storage_data_1016 ^ i_input_data[785 % IN_WIDTH];
                871 / IN_WIDTH: pong_storage_data_1016 <= (fillup_transition == 1'b1) ? i_input_data[871 % IN_WIDTH] : pong_storage_data_1016 ^ i_input_data[871 % IN_WIDTH];
                default: pong_storage_data_1016 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1016;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1016 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1016;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1016 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1016;
            end
        end
    end
end

logic ping_storage_data_1017;
logic pong_storage_data_1017;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1017 <= 1'b0;
        pong_storage_data_1017 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                242 / IN_WIDTH: ping_storage_data_1017 <= (fillup_transition == 1'b1) ? i_input_data[242 % IN_WIDTH] : ping_storage_data_1017 ^ i_input_data[242 % IN_WIDTH];
                376 / IN_WIDTH: ping_storage_data_1017 <= (fillup_transition == 1'b1) ? i_input_data[376 % IN_WIDTH] : ping_storage_data_1017 ^ i_input_data[376 % IN_WIDTH];
                786 / IN_WIDTH: ping_storage_data_1017 <= (fillup_transition == 1'b1) ? i_input_data[786 % IN_WIDTH] : ping_storage_data_1017 ^ i_input_data[786 % IN_WIDTH];
                872 / IN_WIDTH: ping_storage_data_1017 <= (fillup_transition == 1'b1) ? i_input_data[872 % IN_WIDTH] : ping_storage_data_1017 ^ i_input_data[872 % IN_WIDTH];
                default: ping_storage_data_1017 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1017;
                endcase
            end else begin
                case (input_count)
                242 / IN_WIDTH: pong_storage_data_1017 <= (fillup_transition == 1'b1) ? i_input_data[242 % IN_WIDTH] : pong_storage_data_1017 ^ i_input_data[242 % IN_WIDTH];
                376 / IN_WIDTH: pong_storage_data_1017 <= (fillup_transition == 1'b1) ? i_input_data[376 % IN_WIDTH] : pong_storage_data_1017 ^ i_input_data[376 % IN_WIDTH];
                786 / IN_WIDTH: pong_storage_data_1017 <= (fillup_transition == 1'b1) ? i_input_data[786 % IN_WIDTH] : pong_storage_data_1017 ^ i_input_data[786 % IN_WIDTH];
                872 / IN_WIDTH: pong_storage_data_1017 <= (fillup_transition == 1'b1) ? i_input_data[872 % IN_WIDTH] : pong_storage_data_1017 ^ i_input_data[872 % IN_WIDTH];
                default: pong_storage_data_1017 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1017;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1017 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1017;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1017 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1017;
            end
        end
    end
end

logic ping_storage_data_1018;
logic pong_storage_data_1018;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1018 <= 1'b0;
        pong_storage_data_1018 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                243 / IN_WIDTH: ping_storage_data_1018 <= (fillup_transition == 1'b1) ? i_input_data[243 % IN_WIDTH] : ping_storage_data_1018 ^ i_input_data[243 % IN_WIDTH];
                377 / IN_WIDTH: ping_storage_data_1018 <= (fillup_transition == 1'b1) ? i_input_data[377 % IN_WIDTH] : ping_storage_data_1018 ^ i_input_data[377 % IN_WIDTH];
                787 / IN_WIDTH: ping_storage_data_1018 <= (fillup_transition == 1'b1) ? i_input_data[787 % IN_WIDTH] : ping_storage_data_1018 ^ i_input_data[787 % IN_WIDTH];
                873 / IN_WIDTH: ping_storage_data_1018 <= (fillup_transition == 1'b1) ? i_input_data[873 % IN_WIDTH] : ping_storage_data_1018 ^ i_input_data[873 % IN_WIDTH];
                default: ping_storage_data_1018 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1018;
                endcase
            end else begin
                case (input_count)
                243 / IN_WIDTH: pong_storage_data_1018 <= (fillup_transition == 1'b1) ? i_input_data[243 % IN_WIDTH] : pong_storage_data_1018 ^ i_input_data[243 % IN_WIDTH];
                377 / IN_WIDTH: pong_storage_data_1018 <= (fillup_transition == 1'b1) ? i_input_data[377 % IN_WIDTH] : pong_storage_data_1018 ^ i_input_data[377 % IN_WIDTH];
                787 / IN_WIDTH: pong_storage_data_1018 <= (fillup_transition == 1'b1) ? i_input_data[787 % IN_WIDTH] : pong_storage_data_1018 ^ i_input_data[787 % IN_WIDTH];
                873 / IN_WIDTH: pong_storage_data_1018 <= (fillup_transition == 1'b1) ? i_input_data[873 % IN_WIDTH] : pong_storage_data_1018 ^ i_input_data[873 % IN_WIDTH];
                default: pong_storage_data_1018 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1018;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1018 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1018;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1018 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1018;
            end
        end
    end
end

logic ping_storage_data_1019;
logic pong_storage_data_1019;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1019 <= 1'b0;
        pong_storage_data_1019 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                244 / IN_WIDTH: ping_storage_data_1019 <= (fillup_transition == 1'b1) ? i_input_data[244 % IN_WIDTH] : ping_storage_data_1019 ^ i_input_data[244 % IN_WIDTH];
                378 / IN_WIDTH: ping_storage_data_1019 <= (fillup_transition == 1'b1) ? i_input_data[378 % IN_WIDTH] : ping_storage_data_1019 ^ i_input_data[378 % IN_WIDTH];
                788 / IN_WIDTH: ping_storage_data_1019 <= (fillup_transition == 1'b1) ? i_input_data[788 % IN_WIDTH] : ping_storage_data_1019 ^ i_input_data[788 % IN_WIDTH];
                874 / IN_WIDTH: ping_storage_data_1019 <= (fillup_transition == 1'b1) ? i_input_data[874 % IN_WIDTH] : ping_storage_data_1019 ^ i_input_data[874 % IN_WIDTH];
                default: ping_storage_data_1019 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1019;
                endcase
            end else begin
                case (input_count)
                244 / IN_WIDTH: pong_storage_data_1019 <= (fillup_transition == 1'b1) ? i_input_data[244 % IN_WIDTH] : pong_storage_data_1019 ^ i_input_data[244 % IN_WIDTH];
                378 / IN_WIDTH: pong_storage_data_1019 <= (fillup_transition == 1'b1) ? i_input_data[378 % IN_WIDTH] : pong_storage_data_1019 ^ i_input_data[378 % IN_WIDTH];
                788 / IN_WIDTH: pong_storage_data_1019 <= (fillup_transition == 1'b1) ? i_input_data[788 % IN_WIDTH] : pong_storage_data_1019 ^ i_input_data[788 % IN_WIDTH];
                874 / IN_WIDTH: pong_storage_data_1019 <= (fillup_transition == 1'b1) ? i_input_data[874 % IN_WIDTH] : pong_storage_data_1019 ^ i_input_data[874 % IN_WIDTH];
                default: pong_storage_data_1019 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1019;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1019 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1019;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1019 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1019;
            end
        end
    end
end

logic ping_storage_data_1020;
logic pong_storage_data_1020;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1020 <= 1'b0;
        pong_storage_data_1020 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                245 / IN_WIDTH: ping_storage_data_1020 <= (fillup_transition == 1'b1) ? i_input_data[245 % IN_WIDTH] : ping_storage_data_1020 ^ i_input_data[245 % IN_WIDTH];
                379 / IN_WIDTH: ping_storage_data_1020 <= (fillup_transition == 1'b1) ? i_input_data[379 % IN_WIDTH] : ping_storage_data_1020 ^ i_input_data[379 % IN_WIDTH];
                789 / IN_WIDTH: ping_storage_data_1020 <= (fillup_transition == 1'b1) ? i_input_data[789 % IN_WIDTH] : ping_storage_data_1020 ^ i_input_data[789 % IN_WIDTH];
                875 / IN_WIDTH: ping_storage_data_1020 <= (fillup_transition == 1'b1) ? i_input_data[875 % IN_WIDTH] : ping_storage_data_1020 ^ i_input_data[875 % IN_WIDTH];
                default: ping_storage_data_1020 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1020;
                endcase
            end else begin
                case (input_count)
                245 / IN_WIDTH: pong_storage_data_1020 <= (fillup_transition == 1'b1) ? i_input_data[245 % IN_WIDTH] : pong_storage_data_1020 ^ i_input_data[245 % IN_WIDTH];
                379 / IN_WIDTH: pong_storage_data_1020 <= (fillup_transition == 1'b1) ? i_input_data[379 % IN_WIDTH] : pong_storage_data_1020 ^ i_input_data[379 % IN_WIDTH];
                789 / IN_WIDTH: pong_storage_data_1020 <= (fillup_transition == 1'b1) ? i_input_data[789 % IN_WIDTH] : pong_storage_data_1020 ^ i_input_data[789 % IN_WIDTH];
                875 / IN_WIDTH: pong_storage_data_1020 <= (fillup_transition == 1'b1) ? i_input_data[875 % IN_WIDTH] : pong_storage_data_1020 ^ i_input_data[875 % IN_WIDTH];
                default: pong_storage_data_1020 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1020;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1020 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1020;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1020 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1020;
            end
        end
    end
end

logic ping_storage_data_1021;
logic pong_storage_data_1021;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1021 <= 1'b0;
        pong_storage_data_1021 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                246 / IN_WIDTH: ping_storage_data_1021 <= (fillup_transition == 1'b1) ? i_input_data[246 % IN_WIDTH] : ping_storage_data_1021 ^ i_input_data[246 % IN_WIDTH];
                380 / IN_WIDTH: ping_storage_data_1021 <= (fillup_transition == 1'b1) ? i_input_data[380 % IN_WIDTH] : ping_storage_data_1021 ^ i_input_data[380 % IN_WIDTH];
                790 / IN_WIDTH: ping_storage_data_1021 <= (fillup_transition == 1'b1) ? i_input_data[790 % IN_WIDTH] : ping_storage_data_1021 ^ i_input_data[790 % IN_WIDTH];
                876 / IN_WIDTH: ping_storage_data_1021 <= (fillup_transition == 1'b1) ? i_input_data[876 % IN_WIDTH] : ping_storage_data_1021 ^ i_input_data[876 % IN_WIDTH];
                default: ping_storage_data_1021 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1021;
                endcase
            end else begin
                case (input_count)
                246 / IN_WIDTH: pong_storage_data_1021 <= (fillup_transition == 1'b1) ? i_input_data[246 % IN_WIDTH] : pong_storage_data_1021 ^ i_input_data[246 % IN_WIDTH];
                380 / IN_WIDTH: pong_storage_data_1021 <= (fillup_transition == 1'b1) ? i_input_data[380 % IN_WIDTH] : pong_storage_data_1021 ^ i_input_data[380 % IN_WIDTH];
                790 / IN_WIDTH: pong_storage_data_1021 <= (fillup_transition == 1'b1) ? i_input_data[790 % IN_WIDTH] : pong_storage_data_1021 ^ i_input_data[790 % IN_WIDTH];
                876 / IN_WIDTH: pong_storage_data_1021 <= (fillup_transition == 1'b1) ? i_input_data[876 % IN_WIDTH] : pong_storage_data_1021 ^ i_input_data[876 % IN_WIDTH];
                default: pong_storage_data_1021 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1021;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1021 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1021;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1021 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1021;
            end
        end
    end
end

logic ping_storage_data_1022;
logic pong_storage_data_1022;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1022 <= 1'b0;
        pong_storage_data_1022 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                247 / IN_WIDTH: ping_storage_data_1022 <= (fillup_transition == 1'b1) ? i_input_data[247 % IN_WIDTH] : ping_storage_data_1022 ^ i_input_data[247 % IN_WIDTH];
                381 / IN_WIDTH: ping_storage_data_1022 <= (fillup_transition == 1'b1) ? i_input_data[381 % IN_WIDTH] : ping_storage_data_1022 ^ i_input_data[381 % IN_WIDTH];
                791 / IN_WIDTH: ping_storage_data_1022 <= (fillup_transition == 1'b1) ? i_input_data[791 % IN_WIDTH] : ping_storage_data_1022 ^ i_input_data[791 % IN_WIDTH];
                877 / IN_WIDTH: ping_storage_data_1022 <= (fillup_transition == 1'b1) ? i_input_data[877 % IN_WIDTH] : ping_storage_data_1022 ^ i_input_data[877 % IN_WIDTH];
                default: ping_storage_data_1022 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1022;
                endcase
            end else begin
                case (input_count)
                247 / IN_WIDTH: pong_storage_data_1022 <= (fillup_transition == 1'b1) ? i_input_data[247 % IN_WIDTH] : pong_storage_data_1022 ^ i_input_data[247 % IN_WIDTH];
                381 / IN_WIDTH: pong_storage_data_1022 <= (fillup_transition == 1'b1) ? i_input_data[381 % IN_WIDTH] : pong_storage_data_1022 ^ i_input_data[381 % IN_WIDTH];
                791 / IN_WIDTH: pong_storage_data_1022 <= (fillup_transition == 1'b1) ? i_input_data[791 % IN_WIDTH] : pong_storage_data_1022 ^ i_input_data[791 % IN_WIDTH];
                877 / IN_WIDTH: pong_storage_data_1022 <= (fillup_transition == 1'b1) ? i_input_data[877 % IN_WIDTH] : pong_storage_data_1022 ^ i_input_data[877 % IN_WIDTH];
                default: pong_storage_data_1022 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1022;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1022 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1022;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1022 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1022;
            end
        end
    end
end

logic ping_storage_data_1023;
logic pong_storage_data_1023;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1023 <= 1'b0;
        pong_storage_data_1023 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                248 / IN_WIDTH: ping_storage_data_1023 <= (fillup_transition == 1'b1) ? i_input_data[248 % IN_WIDTH] : ping_storage_data_1023 ^ i_input_data[248 % IN_WIDTH];
                382 / IN_WIDTH: ping_storage_data_1023 <= (fillup_transition == 1'b1) ? i_input_data[382 % IN_WIDTH] : ping_storage_data_1023 ^ i_input_data[382 % IN_WIDTH];
                792 / IN_WIDTH: ping_storage_data_1023 <= (fillup_transition == 1'b1) ? i_input_data[792 % IN_WIDTH] : ping_storage_data_1023 ^ i_input_data[792 % IN_WIDTH];
                878 / IN_WIDTH: ping_storage_data_1023 <= (fillup_transition == 1'b1) ? i_input_data[878 % IN_WIDTH] : ping_storage_data_1023 ^ i_input_data[878 % IN_WIDTH];
                default: ping_storage_data_1023 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1023;
                endcase
            end else begin
                case (input_count)
                248 / IN_WIDTH: pong_storage_data_1023 <= (fillup_transition == 1'b1) ? i_input_data[248 % IN_WIDTH] : pong_storage_data_1023 ^ i_input_data[248 % IN_WIDTH];
                382 / IN_WIDTH: pong_storage_data_1023 <= (fillup_transition == 1'b1) ? i_input_data[382 % IN_WIDTH] : pong_storage_data_1023 ^ i_input_data[382 % IN_WIDTH];
                792 / IN_WIDTH: pong_storage_data_1023 <= (fillup_transition == 1'b1) ? i_input_data[792 % IN_WIDTH] : pong_storage_data_1023 ^ i_input_data[792 % IN_WIDTH];
                878 / IN_WIDTH: pong_storage_data_1023 <= (fillup_transition == 1'b1) ? i_input_data[878 % IN_WIDTH] : pong_storage_data_1023 ^ i_input_data[878 % IN_WIDTH];
                default: pong_storage_data_1023 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1023;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1023 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1023;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1023 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1023;
            end
        end
    end
end

logic ping_storage_data_1024;
logic pong_storage_data_1024;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1024 <= 1'b0;
        pong_storage_data_1024 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                249 / IN_WIDTH: ping_storage_data_1024 <= (fillup_transition == 1'b1) ? i_input_data[249 % IN_WIDTH] : ping_storage_data_1024 ^ i_input_data[249 % IN_WIDTH];
                383 / IN_WIDTH: ping_storage_data_1024 <= (fillup_transition == 1'b1) ? i_input_data[383 % IN_WIDTH] : ping_storage_data_1024 ^ i_input_data[383 % IN_WIDTH];
                793 / IN_WIDTH: ping_storage_data_1024 <= (fillup_transition == 1'b1) ? i_input_data[793 % IN_WIDTH] : ping_storage_data_1024 ^ i_input_data[793 % IN_WIDTH];
                879 / IN_WIDTH: ping_storage_data_1024 <= (fillup_transition == 1'b1) ? i_input_data[879 % IN_WIDTH] : ping_storage_data_1024 ^ i_input_data[879 % IN_WIDTH];
                default: ping_storage_data_1024 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1024;
                endcase
            end else begin
                case (input_count)
                249 / IN_WIDTH: pong_storage_data_1024 <= (fillup_transition == 1'b1) ? i_input_data[249 % IN_WIDTH] : pong_storage_data_1024 ^ i_input_data[249 % IN_WIDTH];
                383 / IN_WIDTH: pong_storage_data_1024 <= (fillup_transition == 1'b1) ? i_input_data[383 % IN_WIDTH] : pong_storage_data_1024 ^ i_input_data[383 % IN_WIDTH];
                793 / IN_WIDTH: pong_storage_data_1024 <= (fillup_transition == 1'b1) ? i_input_data[793 % IN_WIDTH] : pong_storage_data_1024 ^ i_input_data[793 % IN_WIDTH];
                879 / IN_WIDTH: pong_storage_data_1024 <= (fillup_transition == 1'b1) ? i_input_data[879 % IN_WIDTH] : pong_storage_data_1024 ^ i_input_data[879 % IN_WIDTH];
                default: pong_storage_data_1024 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1024;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1024 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1024;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1024 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1024;
            end
        end
    end
end

logic ping_storage_data_1025;
logic pong_storage_data_1025;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1025 <= 1'b0;
        pong_storage_data_1025 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                250 / IN_WIDTH: ping_storage_data_1025 <= (fillup_transition == 1'b1) ? i_input_data[250 % IN_WIDTH] : ping_storage_data_1025 ^ i_input_data[250 % IN_WIDTH];
                288 / IN_WIDTH: ping_storage_data_1025 <= (fillup_transition == 1'b1) ? i_input_data[288 % IN_WIDTH] : ping_storage_data_1025 ^ i_input_data[288 % IN_WIDTH];
                794 / IN_WIDTH: ping_storage_data_1025 <= (fillup_transition == 1'b1) ? i_input_data[794 % IN_WIDTH] : ping_storage_data_1025 ^ i_input_data[794 % IN_WIDTH];
                880 / IN_WIDTH: ping_storage_data_1025 <= (fillup_transition == 1'b1) ? i_input_data[880 % IN_WIDTH] : ping_storage_data_1025 ^ i_input_data[880 % IN_WIDTH];
                default: ping_storage_data_1025 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1025;
                endcase
            end else begin
                case (input_count)
                250 / IN_WIDTH: pong_storage_data_1025 <= (fillup_transition == 1'b1) ? i_input_data[250 % IN_WIDTH] : pong_storage_data_1025 ^ i_input_data[250 % IN_WIDTH];
                288 / IN_WIDTH: pong_storage_data_1025 <= (fillup_transition == 1'b1) ? i_input_data[288 % IN_WIDTH] : pong_storage_data_1025 ^ i_input_data[288 % IN_WIDTH];
                794 / IN_WIDTH: pong_storage_data_1025 <= (fillup_transition == 1'b1) ? i_input_data[794 % IN_WIDTH] : pong_storage_data_1025 ^ i_input_data[794 % IN_WIDTH];
                880 / IN_WIDTH: pong_storage_data_1025 <= (fillup_transition == 1'b1) ? i_input_data[880 % IN_WIDTH] : pong_storage_data_1025 ^ i_input_data[880 % IN_WIDTH];
                default: pong_storage_data_1025 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1025;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1025 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1025;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1025 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1025;
            end
        end
    end
end

logic ping_storage_data_1026;
logic pong_storage_data_1026;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1026 <= 1'b0;
        pong_storage_data_1026 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                251 / IN_WIDTH: ping_storage_data_1026 <= (fillup_transition == 1'b1) ? i_input_data[251 % IN_WIDTH] : ping_storage_data_1026 ^ i_input_data[251 % IN_WIDTH];
                289 / IN_WIDTH: ping_storage_data_1026 <= (fillup_transition == 1'b1) ? i_input_data[289 % IN_WIDTH] : ping_storage_data_1026 ^ i_input_data[289 % IN_WIDTH];
                795 / IN_WIDTH: ping_storage_data_1026 <= (fillup_transition == 1'b1) ? i_input_data[795 % IN_WIDTH] : ping_storage_data_1026 ^ i_input_data[795 % IN_WIDTH];
                881 / IN_WIDTH: ping_storage_data_1026 <= (fillup_transition == 1'b1) ? i_input_data[881 % IN_WIDTH] : ping_storage_data_1026 ^ i_input_data[881 % IN_WIDTH];
                default: ping_storage_data_1026 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1026;
                endcase
            end else begin
                case (input_count)
                251 / IN_WIDTH: pong_storage_data_1026 <= (fillup_transition == 1'b1) ? i_input_data[251 % IN_WIDTH] : pong_storage_data_1026 ^ i_input_data[251 % IN_WIDTH];
                289 / IN_WIDTH: pong_storage_data_1026 <= (fillup_transition == 1'b1) ? i_input_data[289 % IN_WIDTH] : pong_storage_data_1026 ^ i_input_data[289 % IN_WIDTH];
                795 / IN_WIDTH: pong_storage_data_1026 <= (fillup_transition == 1'b1) ? i_input_data[795 % IN_WIDTH] : pong_storage_data_1026 ^ i_input_data[795 % IN_WIDTH];
                881 / IN_WIDTH: pong_storage_data_1026 <= (fillup_transition == 1'b1) ? i_input_data[881 % IN_WIDTH] : pong_storage_data_1026 ^ i_input_data[881 % IN_WIDTH];
                default: pong_storage_data_1026 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1026;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1026 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1026;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1026 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1026;
            end
        end
    end
end

logic ping_storage_data_1027;
logic pong_storage_data_1027;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1027 <= 1'b0;
        pong_storage_data_1027 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                252 / IN_WIDTH: ping_storage_data_1027 <= (fillup_transition == 1'b1) ? i_input_data[252 % IN_WIDTH] : ping_storage_data_1027 ^ i_input_data[252 % IN_WIDTH];
                290 / IN_WIDTH: ping_storage_data_1027 <= (fillup_transition == 1'b1) ? i_input_data[290 % IN_WIDTH] : ping_storage_data_1027 ^ i_input_data[290 % IN_WIDTH];
                796 / IN_WIDTH: ping_storage_data_1027 <= (fillup_transition == 1'b1) ? i_input_data[796 % IN_WIDTH] : ping_storage_data_1027 ^ i_input_data[796 % IN_WIDTH];
                882 / IN_WIDTH: ping_storage_data_1027 <= (fillup_transition == 1'b1) ? i_input_data[882 % IN_WIDTH] : ping_storage_data_1027 ^ i_input_data[882 % IN_WIDTH];
                default: ping_storage_data_1027 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1027;
                endcase
            end else begin
                case (input_count)
                252 / IN_WIDTH: pong_storage_data_1027 <= (fillup_transition == 1'b1) ? i_input_data[252 % IN_WIDTH] : pong_storage_data_1027 ^ i_input_data[252 % IN_WIDTH];
                290 / IN_WIDTH: pong_storage_data_1027 <= (fillup_transition == 1'b1) ? i_input_data[290 % IN_WIDTH] : pong_storage_data_1027 ^ i_input_data[290 % IN_WIDTH];
                796 / IN_WIDTH: pong_storage_data_1027 <= (fillup_transition == 1'b1) ? i_input_data[796 % IN_WIDTH] : pong_storage_data_1027 ^ i_input_data[796 % IN_WIDTH];
                882 / IN_WIDTH: pong_storage_data_1027 <= (fillup_transition == 1'b1) ? i_input_data[882 % IN_WIDTH] : pong_storage_data_1027 ^ i_input_data[882 % IN_WIDTH];
                default: pong_storage_data_1027 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1027;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1027 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1027;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1027 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1027;
            end
        end
    end
end

logic ping_storage_data_1028;
logic pong_storage_data_1028;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1028 <= 1'b0;
        pong_storage_data_1028 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                253 / IN_WIDTH: ping_storage_data_1028 <= (fillup_transition == 1'b1) ? i_input_data[253 % IN_WIDTH] : ping_storage_data_1028 ^ i_input_data[253 % IN_WIDTH];
                291 / IN_WIDTH: ping_storage_data_1028 <= (fillup_transition == 1'b1) ? i_input_data[291 % IN_WIDTH] : ping_storage_data_1028 ^ i_input_data[291 % IN_WIDTH];
                797 / IN_WIDTH: ping_storage_data_1028 <= (fillup_transition == 1'b1) ? i_input_data[797 % IN_WIDTH] : ping_storage_data_1028 ^ i_input_data[797 % IN_WIDTH];
                883 / IN_WIDTH: ping_storage_data_1028 <= (fillup_transition == 1'b1) ? i_input_data[883 % IN_WIDTH] : ping_storage_data_1028 ^ i_input_data[883 % IN_WIDTH];
                default: ping_storage_data_1028 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1028;
                endcase
            end else begin
                case (input_count)
                253 / IN_WIDTH: pong_storage_data_1028 <= (fillup_transition == 1'b1) ? i_input_data[253 % IN_WIDTH] : pong_storage_data_1028 ^ i_input_data[253 % IN_WIDTH];
                291 / IN_WIDTH: pong_storage_data_1028 <= (fillup_transition == 1'b1) ? i_input_data[291 % IN_WIDTH] : pong_storage_data_1028 ^ i_input_data[291 % IN_WIDTH];
                797 / IN_WIDTH: pong_storage_data_1028 <= (fillup_transition == 1'b1) ? i_input_data[797 % IN_WIDTH] : pong_storage_data_1028 ^ i_input_data[797 % IN_WIDTH];
                883 / IN_WIDTH: pong_storage_data_1028 <= (fillup_transition == 1'b1) ? i_input_data[883 % IN_WIDTH] : pong_storage_data_1028 ^ i_input_data[883 % IN_WIDTH];
                default: pong_storage_data_1028 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1028;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1028 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1028;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1028 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1028;
            end
        end
    end
end

logic ping_storage_data_1029;
logic pong_storage_data_1029;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1029 <= 1'b0;
        pong_storage_data_1029 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                254 / IN_WIDTH: ping_storage_data_1029 <= (fillup_transition == 1'b1) ? i_input_data[254 % IN_WIDTH] : ping_storage_data_1029 ^ i_input_data[254 % IN_WIDTH];
                292 / IN_WIDTH: ping_storage_data_1029 <= (fillup_transition == 1'b1) ? i_input_data[292 % IN_WIDTH] : ping_storage_data_1029 ^ i_input_data[292 % IN_WIDTH];
                798 / IN_WIDTH: ping_storage_data_1029 <= (fillup_transition == 1'b1) ? i_input_data[798 % IN_WIDTH] : ping_storage_data_1029 ^ i_input_data[798 % IN_WIDTH];
                884 / IN_WIDTH: ping_storage_data_1029 <= (fillup_transition == 1'b1) ? i_input_data[884 % IN_WIDTH] : ping_storage_data_1029 ^ i_input_data[884 % IN_WIDTH];
                default: ping_storage_data_1029 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1029;
                endcase
            end else begin
                case (input_count)
                254 / IN_WIDTH: pong_storage_data_1029 <= (fillup_transition == 1'b1) ? i_input_data[254 % IN_WIDTH] : pong_storage_data_1029 ^ i_input_data[254 % IN_WIDTH];
                292 / IN_WIDTH: pong_storage_data_1029 <= (fillup_transition == 1'b1) ? i_input_data[292 % IN_WIDTH] : pong_storage_data_1029 ^ i_input_data[292 % IN_WIDTH];
                798 / IN_WIDTH: pong_storage_data_1029 <= (fillup_transition == 1'b1) ? i_input_data[798 % IN_WIDTH] : pong_storage_data_1029 ^ i_input_data[798 % IN_WIDTH];
                884 / IN_WIDTH: pong_storage_data_1029 <= (fillup_transition == 1'b1) ? i_input_data[884 % IN_WIDTH] : pong_storage_data_1029 ^ i_input_data[884 % IN_WIDTH];
                default: pong_storage_data_1029 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1029;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1029 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1029;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1029 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1029;
            end
        end
    end
end

logic ping_storage_data_1030;
logic pong_storage_data_1030;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1030 <= 1'b0;
        pong_storage_data_1030 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                255 / IN_WIDTH: ping_storage_data_1030 <= (fillup_transition == 1'b1) ? i_input_data[255 % IN_WIDTH] : ping_storage_data_1030 ^ i_input_data[255 % IN_WIDTH];
                293 / IN_WIDTH: ping_storage_data_1030 <= (fillup_transition == 1'b1) ? i_input_data[293 % IN_WIDTH] : ping_storage_data_1030 ^ i_input_data[293 % IN_WIDTH];
                799 / IN_WIDTH: ping_storage_data_1030 <= (fillup_transition == 1'b1) ? i_input_data[799 % IN_WIDTH] : ping_storage_data_1030 ^ i_input_data[799 % IN_WIDTH];
                885 / IN_WIDTH: ping_storage_data_1030 <= (fillup_transition == 1'b1) ? i_input_data[885 % IN_WIDTH] : ping_storage_data_1030 ^ i_input_data[885 % IN_WIDTH];
                default: ping_storage_data_1030 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1030;
                endcase
            end else begin
                case (input_count)
                255 / IN_WIDTH: pong_storage_data_1030 <= (fillup_transition == 1'b1) ? i_input_data[255 % IN_WIDTH] : pong_storage_data_1030 ^ i_input_data[255 % IN_WIDTH];
                293 / IN_WIDTH: pong_storage_data_1030 <= (fillup_transition == 1'b1) ? i_input_data[293 % IN_WIDTH] : pong_storage_data_1030 ^ i_input_data[293 % IN_WIDTH];
                799 / IN_WIDTH: pong_storage_data_1030 <= (fillup_transition == 1'b1) ? i_input_data[799 % IN_WIDTH] : pong_storage_data_1030 ^ i_input_data[799 % IN_WIDTH];
                885 / IN_WIDTH: pong_storage_data_1030 <= (fillup_transition == 1'b1) ? i_input_data[885 % IN_WIDTH] : pong_storage_data_1030 ^ i_input_data[885 % IN_WIDTH];
                default: pong_storage_data_1030 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1030;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1030 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1030;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1030 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1030;
            end
        end
    end
end

logic ping_storage_data_1031;
logic pong_storage_data_1031;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1031 <= 1'b0;
        pong_storage_data_1031 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                256 / IN_WIDTH: ping_storage_data_1031 <= (fillup_transition == 1'b1) ? i_input_data[256 % IN_WIDTH] : ping_storage_data_1031 ^ i_input_data[256 % IN_WIDTH];
                294 / IN_WIDTH: ping_storage_data_1031 <= (fillup_transition == 1'b1) ? i_input_data[294 % IN_WIDTH] : ping_storage_data_1031 ^ i_input_data[294 % IN_WIDTH];
                800 / IN_WIDTH: ping_storage_data_1031 <= (fillup_transition == 1'b1) ? i_input_data[800 % IN_WIDTH] : ping_storage_data_1031 ^ i_input_data[800 % IN_WIDTH];
                886 / IN_WIDTH: ping_storage_data_1031 <= (fillup_transition == 1'b1) ? i_input_data[886 % IN_WIDTH] : ping_storage_data_1031 ^ i_input_data[886 % IN_WIDTH];
                default: ping_storage_data_1031 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1031;
                endcase
            end else begin
                case (input_count)
                256 / IN_WIDTH: pong_storage_data_1031 <= (fillup_transition == 1'b1) ? i_input_data[256 % IN_WIDTH] : pong_storage_data_1031 ^ i_input_data[256 % IN_WIDTH];
                294 / IN_WIDTH: pong_storage_data_1031 <= (fillup_transition == 1'b1) ? i_input_data[294 % IN_WIDTH] : pong_storage_data_1031 ^ i_input_data[294 % IN_WIDTH];
                800 / IN_WIDTH: pong_storage_data_1031 <= (fillup_transition == 1'b1) ? i_input_data[800 % IN_WIDTH] : pong_storage_data_1031 ^ i_input_data[800 % IN_WIDTH];
                886 / IN_WIDTH: pong_storage_data_1031 <= (fillup_transition == 1'b1) ? i_input_data[886 % IN_WIDTH] : pong_storage_data_1031 ^ i_input_data[886 % IN_WIDTH];
                default: pong_storage_data_1031 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1031;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1031 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1031;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1031 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1031;
            end
        end
    end
end

logic ping_storage_data_1032;
logic pong_storage_data_1032;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1032 <= 1'b0;
        pong_storage_data_1032 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                257 / IN_WIDTH: ping_storage_data_1032 <= (fillup_transition == 1'b1) ? i_input_data[257 % IN_WIDTH] : ping_storage_data_1032 ^ i_input_data[257 % IN_WIDTH];
                295 / IN_WIDTH: ping_storage_data_1032 <= (fillup_transition == 1'b1) ? i_input_data[295 % IN_WIDTH] : ping_storage_data_1032 ^ i_input_data[295 % IN_WIDTH];
                801 / IN_WIDTH: ping_storage_data_1032 <= (fillup_transition == 1'b1) ? i_input_data[801 % IN_WIDTH] : ping_storage_data_1032 ^ i_input_data[801 % IN_WIDTH];
                887 / IN_WIDTH: ping_storage_data_1032 <= (fillup_transition == 1'b1) ? i_input_data[887 % IN_WIDTH] : ping_storage_data_1032 ^ i_input_data[887 % IN_WIDTH];
                default: ping_storage_data_1032 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1032;
                endcase
            end else begin
                case (input_count)
                257 / IN_WIDTH: pong_storage_data_1032 <= (fillup_transition == 1'b1) ? i_input_data[257 % IN_WIDTH] : pong_storage_data_1032 ^ i_input_data[257 % IN_WIDTH];
                295 / IN_WIDTH: pong_storage_data_1032 <= (fillup_transition == 1'b1) ? i_input_data[295 % IN_WIDTH] : pong_storage_data_1032 ^ i_input_data[295 % IN_WIDTH];
                801 / IN_WIDTH: pong_storage_data_1032 <= (fillup_transition == 1'b1) ? i_input_data[801 % IN_WIDTH] : pong_storage_data_1032 ^ i_input_data[801 % IN_WIDTH];
                887 / IN_WIDTH: pong_storage_data_1032 <= (fillup_transition == 1'b1) ? i_input_data[887 % IN_WIDTH] : pong_storage_data_1032 ^ i_input_data[887 % IN_WIDTH];
                default: pong_storage_data_1032 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1032;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1032 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1032;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1032 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1032;
            end
        end
    end
end

logic ping_storage_data_1033;
logic pong_storage_data_1033;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1033 <= 1'b0;
        pong_storage_data_1033 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                258 / IN_WIDTH: ping_storage_data_1033 <= (fillup_transition == 1'b1) ? i_input_data[258 % IN_WIDTH] : ping_storage_data_1033 ^ i_input_data[258 % IN_WIDTH];
                296 / IN_WIDTH: ping_storage_data_1033 <= (fillup_transition == 1'b1) ? i_input_data[296 % IN_WIDTH] : ping_storage_data_1033 ^ i_input_data[296 % IN_WIDTH];
                802 / IN_WIDTH: ping_storage_data_1033 <= (fillup_transition == 1'b1) ? i_input_data[802 % IN_WIDTH] : ping_storage_data_1033 ^ i_input_data[802 % IN_WIDTH];
                888 / IN_WIDTH: ping_storage_data_1033 <= (fillup_transition == 1'b1) ? i_input_data[888 % IN_WIDTH] : ping_storage_data_1033 ^ i_input_data[888 % IN_WIDTH];
                default: ping_storage_data_1033 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1033;
                endcase
            end else begin
                case (input_count)
                258 / IN_WIDTH: pong_storage_data_1033 <= (fillup_transition == 1'b1) ? i_input_data[258 % IN_WIDTH] : pong_storage_data_1033 ^ i_input_data[258 % IN_WIDTH];
                296 / IN_WIDTH: pong_storage_data_1033 <= (fillup_transition == 1'b1) ? i_input_data[296 % IN_WIDTH] : pong_storage_data_1033 ^ i_input_data[296 % IN_WIDTH];
                802 / IN_WIDTH: pong_storage_data_1033 <= (fillup_transition == 1'b1) ? i_input_data[802 % IN_WIDTH] : pong_storage_data_1033 ^ i_input_data[802 % IN_WIDTH];
                888 / IN_WIDTH: pong_storage_data_1033 <= (fillup_transition == 1'b1) ? i_input_data[888 % IN_WIDTH] : pong_storage_data_1033 ^ i_input_data[888 % IN_WIDTH];
                default: pong_storage_data_1033 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1033;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1033 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1033;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1033 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1033;
            end
        end
    end
end

logic ping_storage_data_1034;
logic pong_storage_data_1034;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1034 <= 1'b0;
        pong_storage_data_1034 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                259 / IN_WIDTH: ping_storage_data_1034 <= (fillup_transition == 1'b1) ? i_input_data[259 % IN_WIDTH] : ping_storage_data_1034 ^ i_input_data[259 % IN_WIDTH];
                297 / IN_WIDTH: ping_storage_data_1034 <= (fillup_transition == 1'b1) ? i_input_data[297 % IN_WIDTH] : ping_storage_data_1034 ^ i_input_data[297 % IN_WIDTH];
                803 / IN_WIDTH: ping_storage_data_1034 <= (fillup_transition == 1'b1) ? i_input_data[803 % IN_WIDTH] : ping_storage_data_1034 ^ i_input_data[803 % IN_WIDTH];
                889 / IN_WIDTH: ping_storage_data_1034 <= (fillup_transition == 1'b1) ? i_input_data[889 % IN_WIDTH] : ping_storage_data_1034 ^ i_input_data[889 % IN_WIDTH];
                default: ping_storage_data_1034 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1034;
                endcase
            end else begin
                case (input_count)
                259 / IN_WIDTH: pong_storage_data_1034 <= (fillup_transition == 1'b1) ? i_input_data[259 % IN_WIDTH] : pong_storage_data_1034 ^ i_input_data[259 % IN_WIDTH];
                297 / IN_WIDTH: pong_storage_data_1034 <= (fillup_transition == 1'b1) ? i_input_data[297 % IN_WIDTH] : pong_storage_data_1034 ^ i_input_data[297 % IN_WIDTH];
                803 / IN_WIDTH: pong_storage_data_1034 <= (fillup_transition == 1'b1) ? i_input_data[803 % IN_WIDTH] : pong_storage_data_1034 ^ i_input_data[803 % IN_WIDTH];
                889 / IN_WIDTH: pong_storage_data_1034 <= (fillup_transition == 1'b1) ? i_input_data[889 % IN_WIDTH] : pong_storage_data_1034 ^ i_input_data[889 % IN_WIDTH];
                default: pong_storage_data_1034 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1034;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1034 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1034;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1034 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1034;
            end
        end
    end
end

logic ping_storage_data_1035;
logic pong_storage_data_1035;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1035 <= 1'b0;
        pong_storage_data_1035 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                260 / IN_WIDTH: ping_storage_data_1035 <= (fillup_transition == 1'b1) ? i_input_data[260 % IN_WIDTH] : ping_storage_data_1035 ^ i_input_data[260 % IN_WIDTH];
                298 / IN_WIDTH: ping_storage_data_1035 <= (fillup_transition == 1'b1) ? i_input_data[298 % IN_WIDTH] : ping_storage_data_1035 ^ i_input_data[298 % IN_WIDTH];
                804 / IN_WIDTH: ping_storage_data_1035 <= (fillup_transition == 1'b1) ? i_input_data[804 % IN_WIDTH] : ping_storage_data_1035 ^ i_input_data[804 % IN_WIDTH];
                890 / IN_WIDTH: ping_storage_data_1035 <= (fillup_transition == 1'b1) ? i_input_data[890 % IN_WIDTH] : ping_storage_data_1035 ^ i_input_data[890 % IN_WIDTH];
                default: ping_storage_data_1035 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1035;
                endcase
            end else begin
                case (input_count)
                260 / IN_WIDTH: pong_storage_data_1035 <= (fillup_transition == 1'b1) ? i_input_data[260 % IN_WIDTH] : pong_storage_data_1035 ^ i_input_data[260 % IN_WIDTH];
                298 / IN_WIDTH: pong_storage_data_1035 <= (fillup_transition == 1'b1) ? i_input_data[298 % IN_WIDTH] : pong_storage_data_1035 ^ i_input_data[298 % IN_WIDTH];
                804 / IN_WIDTH: pong_storage_data_1035 <= (fillup_transition == 1'b1) ? i_input_data[804 % IN_WIDTH] : pong_storage_data_1035 ^ i_input_data[804 % IN_WIDTH];
                890 / IN_WIDTH: pong_storage_data_1035 <= (fillup_transition == 1'b1) ? i_input_data[890 % IN_WIDTH] : pong_storage_data_1035 ^ i_input_data[890 % IN_WIDTH];
                default: pong_storage_data_1035 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1035;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1035 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1035;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1035 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1035;
            end
        end
    end
end

logic ping_storage_data_1036;
logic pong_storage_data_1036;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1036 <= 1'b0;
        pong_storage_data_1036 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                261 / IN_WIDTH: ping_storage_data_1036 <= (fillup_transition == 1'b1) ? i_input_data[261 % IN_WIDTH] : ping_storage_data_1036 ^ i_input_data[261 % IN_WIDTH];
                299 / IN_WIDTH: ping_storage_data_1036 <= (fillup_transition == 1'b1) ? i_input_data[299 % IN_WIDTH] : ping_storage_data_1036 ^ i_input_data[299 % IN_WIDTH];
                805 / IN_WIDTH: ping_storage_data_1036 <= (fillup_transition == 1'b1) ? i_input_data[805 % IN_WIDTH] : ping_storage_data_1036 ^ i_input_data[805 % IN_WIDTH];
                891 / IN_WIDTH: ping_storage_data_1036 <= (fillup_transition == 1'b1) ? i_input_data[891 % IN_WIDTH] : ping_storage_data_1036 ^ i_input_data[891 % IN_WIDTH];
                default: ping_storage_data_1036 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1036;
                endcase
            end else begin
                case (input_count)
                261 / IN_WIDTH: pong_storage_data_1036 <= (fillup_transition == 1'b1) ? i_input_data[261 % IN_WIDTH] : pong_storage_data_1036 ^ i_input_data[261 % IN_WIDTH];
                299 / IN_WIDTH: pong_storage_data_1036 <= (fillup_transition == 1'b1) ? i_input_data[299 % IN_WIDTH] : pong_storage_data_1036 ^ i_input_data[299 % IN_WIDTH];
                805 / IN_WIDTH: pong_storage_data_1036 <= (fillup_transition == 1'b1) ? i_input_data[805 % IN_WIDTH] : pong_storage_data_1036 ^ i_input_data[805 % IN_WIDTH];
                891 / IN_WIDTH: pong_storage_data_1036 <= (fillup_transition == 1'b1) ? i_input_data[891 % IN_WIDTH] : pong_storage_data_1036 ^ i_input_data[891 % IN_WIDTH];
                default: pong_storage_data_1036 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1036;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1036 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1036;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1036 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1036;
            end
        end
    end
end

logic ping_storage_data_1037;
logic pong_storage_data_1037;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1037 <= 1'b0;
        pong_storage_data_1037 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                262 / IN_WIDTH: ping_storage_data_1037 <= (fillup_transition == 1'b1) ? i_input_data[262 % IN_WIDTH] : ping_storage_data_1037 ^ i_input_data[262 % IN_WIDTH];
                300 / IN_WIDTH: ping_storage_data_1037 <= (fillup_transition == 1'b1) ? i_input_data[300 % IN_WIDTH] : ping_storage_data_1037 ^ i_input_data[300 % IN_WIDTH];
                806 / IN_WIDTH: ping_storage_data_1037 <= (fillup_transition == 1'b1) ? i_input_data[806 % IN_WIDTH] : ping_storage_data_1037 ^ i_input_data[806 % IN_WIDTH];
                892 / IN_WIDTH: ping_storage_data_1037 <= (fillup_transition == 1'b1) ? i_input_data[892 % IN_WIDTH] : ping_storage_data_1037 ^ i_input_data[892 % IN_WIDTH];
                default: ping_storage_data_1037 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1037;
                endcase
            end else begin
                case (input_count)
                262 / IN_WIDTH: pong_storage_data_1037 <= (fillup_transition == 1'b1) ? i_input_data[262 % IN_WIDTH] : pong_storage_data_1037 ^ i_input_data[262 % IN_WIDTH];
                300 / IN_WIDTH: pong_storage_data_1037 <= (fillup_transition == 1'b1) ? i_input_data[300 % IN_WIDTH] : pong_storage_data_1037 ^ i_input_data[300 % IN_WIDTH];
                806 / IN_WIDTH: pong_storage_data_1037 <= (fillup_transition == 1'b1) ? i_input_data[806 % IN_WIDTH] : pong_storage_data_1037 ^ i_input_data[806 % IN_WIDTH];
                892 / IN_WIDTH: pong_storage_data_1037 <= (fillup_transition == 1'b1) ? i_input_data[892 % IN_WIDTH] : pong_storage_data_1037 ^ i_input_data[892 % IN_WIDTH];
                default: pong_storage_data_1037 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1037;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1037 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1037;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1037 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1037;
            end
        end
    end
end

logic ping_storage_data_1038;
logic pong_storage_data_1038;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1038 <= 1'b0;
        pong_storage_data_1038 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                263 / IN_WIDTH: ping_storage_data_1038 <= (fillup_transition == 1'b1) ? i_input_data[263 % IN_WIDTH] : ping_storage_data_1038 ^ i_input_data[263 % IN_WIDTH];
                301 / IN_WIDTH: ping_storage_data_1038 <= (fillup_transition == 1'b1) ? i_input_data[301 % IN_WIDTH] : ping_storage_data_1038 ^ i_input_data[301 % IN_WIDTH];
                807 / IN_WIDTH: ping_storage_data_1038 <= (fillup_transition == 1'b1) ? i_input_data[807 % IN_WIDTH] : ping_storage_data_1038 ^ i_input_data[807 % IN_WIDTH];
                893 / IN_WIDTH: ping_storage_data_1038 <= (fillup_transition == 1'b1) ? i_input_data[893 % IN_WIDTH] : ping_storage_data_1038 ^ i_input_data[893 % IN_WIDTH];
                default: ping_storage_data_1038 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1038;
                endcase
            end else begin
                case (input_count)
                263 / IN_WIDTH: pong_storage_data_1038 <= (fillup_transition == 1'b1) ? i_input_data[263 % IN_WIDTH] : pong_storage_data_1038 ^ i_input_data[263 % IN_WIDTH];
                301 / IN_WIDTH: pong_storage_data_1038 <= (fillup_transition == 1'b1) ? i_input_data[301 % IN_WIDTH] : pong_storage_data_1038 ^ i_input_data[301 % IN_WIDTH];
                807 / IN_WIDTH: pong_storage_data_1038 <= (fillup_transition == 1'b1) ? i_input_data[807 % IN_WIDTH] : pong_storage_data_1038 ^ i_input_data[807 % IN_WIDTH];
                893 / IN_WIDTH: pong_storage_data_1038 <= (fillup_transition == 1'b1) ? i_input_data[893 % IN_WIDTH] : pong_storage_data_1038 ^ i_input_data[893 % IN_WIDTH];
                default: pong_storage_data_1038 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1038;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1038 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1038;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1038 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1038;
            end
        end
    end
end

logic ping_storage_data_1039;
logic pong_storage_data_1039;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1039 <= 1'b0;
        pong_storage_data_1039 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                264 / IN_WIDTH: ping_storage_data_1039 <= (fillup_transition == 1'b1) ? i_input_data[264 % IN_WIDTH] : ping_storage_data_1039 ^ i_input_data[264 % IN_WIDTH];
                302 / IN_WIDTH: ping_storage_data_1039 <= (fillup_transition == 1'b1) ? i_input_data[302 % IN_WIDTH] : ping_storage_data_1039 ^ i_input_data[302 % IN_WIDTH];
                808 / IN_WIDTH: ping_storage_data_1039 <= (fillup_transition == 1'b1) ? i_input_data[808 % IN_WIDTH] : ping_storage_data_1039 ^ i_input_data[808 % IN_WIDTH];
                894 / IN_WIDTH: ping_storage_data_1039 <= (fillup_transition == 1'b1) ? i_input_data[894 % IN_WIDTH] : ping_storage_data_1039 ^ i_input_data[894 % IN_WIDTH];
                default: ping_storage_data_1039 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1039;
                endcase
            end else begin
                case (input_count)
                264 / IN_WIDTH: pong_storage_data_1039 <= (fillup_transition == 1'b1) ? i_input_data[264 % IN_WIDTH] : pong_storage_data_1039 ^ i_input_data[264 % IN_WIDTH];
                302 / IN_WIDTH: pong_storage_data_1039 <= (fillup_transition == 1'b1) ? i_input_data[302 % IN_WIDTH] : pong_storage_data_1039 ^ i_input_data[302 % IN_WIDTH];
                808 / IN_WIDTH: pong_storage_data_1039 <= (fillup_transition == 1'b1) ? i_input_data[808 % IN_WIDTH] : pong_storage_data_1039 ^ i_input_data[808 % IN_WIDTH];
                894 / IN_WIDTH: pong_storage_data_1039 <= (fillup_transition == 1'b1) ? i_input_data[894 % IN_WIDTH] : pong_storage_data_1039 ^ i_input_data[894 % IN_WIDTH];
                default: pong_storage_data_1039 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1039;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1039 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1039;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1039 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1039;
            end
        end
    end
end

logic ping_storage_data_1040;
logic pong_storage_data_1040;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1040 <= 1'b0;
        pong_storage_data_1040 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                265 / IN_WIDTH: ping_storage_data_1040 <= (fillup_transition == 1'b1) ? i_input_data[265 % IN_WIDTH] : ping_storage_data_1040 ^ i_input_data[265 % IN_WIDTH];
                303 / IN_WIDTH: ping_storage_data_1040 <= (fillup_transition == 1'b1) ? i_input_data[303 % IN_WIDTH] : ping_storage_data_1040 ^ i_input_data[303 % IN_WIDTH];
                809 / IN_WIDTH: ping_storage_data_1040 <= (fillup_transition == 1'b1) ? i_input_data[809 % IN_WIDTH] : ping_storage_data_1040 ^ i_input_data[809 % IN_WIDTH];
                895 / IN_WIDTH: ping_storage_data_1040 <= (fillup_transition == 1'b1) ? i_input_data[895 % IN_WIDTH] : ping_storage_data_1040 ^ i_input_data[895 % IN_WIDTH];
                default: ping_storage_data_1040 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1040;
                endcase
            end else begin
                case (input_count)
                265 / IN_WIDTH: pong_storage_data_1040 <= (fillup_transition == 1'b1) ? i_input_data[265 % IN_WIDTH] : pong_storage_data_1040 ^ i_input_data[265 % IN_WIDTH];
                303 / IN_WIDTH: pong_storage_data_1040 <= (fillup_transition == 1'b1) ? i_input_data[303 % IN_WIDTH] : pong_storage_data_1040 ^ i_input_data[303 % IN_WIDTH];
                809 / IN_WIDTH: pong_storage_data_1040 <= (fillup_transition == 1'b1) ? i_input_data[809 % IN_WIDTH] : pong_storage_data_1040 ^ i_input_data[809 % IN_WIDTH];
                895 / IN_WIDTH: pong_storage_data_1040 <= (fillup_transition == 1'b1) ? i_input_data[895 % IN_WIDTH] : pong_storage_data_1040 ^ i_input_data[895 % IN_WIDTH];
                default: pong_storage_data_1040 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1040;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1040 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1040;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1040 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1040;
            end
        end
    end
end

logic ping_storage_data_1041;
logic pong_storage_data_1041;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1041 <= 1'b0;
        pong_storage_data_1041 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                266 / IN_WIDTH: ping_storage_data_1041 <= (fillup_transition == 1'b1) ? i_input_data[266 % IN_WIDTH] : ping_storage_data_1041 ^ i_input_data[266 % IN_WIDTH];
                304 / IN_WIDTH: ping_storage_data_1041 <= (fillup_transition == 1'b1) ? i_input_data[304 % IN_WIDTH] : ping_storage_data_1041 ^ i_input_data[304 % IN_WIDTH];
                810 / IN_WIDTH: ping_storage_data_1041 <= (fillup_transition == 1'b1) ? i_input_data[810 % IN_WIDTH] : ping_storage_data_1041 ^ i_input_data[810 % IN_WIDTH];
                896 / IN_WIDTH: ping_storage_data_1041 <= (fillup_transition == 1'b1) ? i_input_data[896 % IN_WIDTH] : ping_storage_data_1041 ^ i_input_data[896 % IN_WIDTH];
                default: ping_storage_data_1041 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1041;
                endcase
            end else begin
                case (input_count)
                266 / IN_WIDTH: pong_storage_data_1041 <= (fillup_transition == 1'b1) ? i_input_data[266 % IN_WIDTH] : pong_storage_data_1041 ^ i_input_data[266 % IN_WIDTH];
                304 / IN_WIDTH: pong_storage_data_1041 <= (fillup_transition == 1'b1) ? i_input_data[304 % IN_WIDTH] : pong_storage_data_1041 ^ i_input_data[304 % IN_WIDTH];
                810 / IN_WIDTH: pong_storage_data_1041 <= (fillup_transition == 1'b1) ? i_input_data[810 % IN_WIDTH] : pong_storage_data_1041 ^ i_input_data[810 % IN_WIDTH];
                896 / IN_WIDTH: pong_storage_data_1041 <= (fillup_transition == 1'b1) ? i_input_data[896 % IN_WIDTH] : pong_storage_data_1041 ^ i_input_data[896 % IN_WIDTH];
                default: pong_storage_data_1041 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1041;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1041 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1041;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1041 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1041;
            end
        end
    end
end

logic ping_storage_data_1042;
logic pong_storage_data_1042;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1042 <= 1'b0;
        pong_storage_data_1042 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                267 / IN_WIDTH: ping_storage_data_1042 <= (fillup_transition == 1'b1) ? i_input_data[267 % IN_WIDTH] : ping_storage_data_1042 ^ i_input_data[267 % IN_WIDTH];
                305 / IN_WIDTH: ping_storage_data_1042 <= (fillup_transition == 1'b1) ? i_input_data[305 % IN_WIDTH] : ping_storage_data_1042 ^ i_input_data[305 % IN_WIDTH];
                811 / IN_WIDTH: ping_storage_data_1042 <= (fillup_transition == 1'b1) ? i_input_data[811 % IN_WIDTH] : ping_storage_data_1042 ^ i_input_data[811 % IN_WIDTH];
                897 / IN_WIDTH: ping_storage_data_1042 <= (fillup_transition == 1'b1) ? i_input_data[897 % IN_WIDTH] : ping_storage_data_1042 ^ i_input_data[897 % IN_WIDTH];
                default: ping_storage_data_1042 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1042;
                endcase
            end else begin
                case (input_count)
                267 / IN_WIDTH: pong_storage_data_1042 <= (fillup_transition == 1'b1) ? i_input_data[267 % IN_WIDTH] : pong_storage_data_1042 ^ i_input_data[267 % IN_WIDTH];
                305 / IN_WIDTH: pong_storage_data_1042 <= (fillup_transition == 1'b1) ? i_input_data[305 % IN_WIDTH] : pong_storage_data_1042 ^ i_input_data[305 % IN_WIDTH];
                811 / IN_WIDTH: pong_storage_data_1042 <= (fillup_transition == 1'b1) ? i_input_data[811 % IN_WIDTH] : pong_storage_data_1042 ^ i_input_data[811 % IN_WIDTH];
                897 / IN_WIDTH: pong_storage_data_1042 <= (fillup_transition == 1'b1) ? i_input_data[897 % IN_WIDTH] : pong_storage_data_1042 ^ i_input_data[897 % IN_WIDTH];
                default: pong_storage_data_1042 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1042;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1042 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1042;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1042 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1042;
            end
        end
    end
end

logic ping_storage_data_1043;
logic pong_storage_data_1043;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1043 <= 1'b0;
        pong_storage_data_1043 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                268 / IN_WIDTH: ping_storage_data_1043 <= (fillup_transition == 1'b1) ? i_input_data[268 % IN_WIDTH] : ping_storage_data_1043 ^ i_input_data[268 % IN_WIDTH];
                306 / IN_WIDTH: ping_storage_data_1043 <= (fillup_transition == 1'b1) ? i_input_data[306 % IN_WIDTH] : ping_storage_data_1043 ^ i_input_data[306 % IN_WIDTH];
                812 / IN_WIDTH: ping_storage_data_1043 <= (fillup_transition == 1'b1) ? i_input_data[812 % IN_WIDTH] : ping_storage_data_1043 ^ i_input_data[812 % IN_WIDTH];
                898 / IN_WIDTH: ping_storage_data_1043 <= (fillup_transition == 1'b1) ? i_input_data[898 % IN_WIDTH] : ping_storage_data_1043 ^ i_input_data[898 % IN_WIDTH];
                default: ping_storage_data_1043 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1043;
                endcase
            end else begin
                case (input_count)
                268 / IN_WIDTH: pong_storage_data_1043 <= (fillup_transition == 1'b1) ? i_input_data[268 % IN_WIDTH] : pong_storage_data_1043 ^ i_input_data[268 % IN_WIDTH];
                306 / IN_WIDTH: pong_storage_data_1043 <= (fillup_transition == 1'b1) ? i_input_data[306 % IN_WIDTH] : pong_storage_data_1043 ^ i_input_data[306 % IN_WIDTH];
                812 / IN_WIDTH: pong_storage_data_1043 <= (fillup_transition == 1'b1) ? i_input_data[812 % IN_WIDTH] : pong_storage_data_1043 ^ i_input_data[812 % IN_WIDTH];
                898 / IN_WIDTH: pong_storage_data_1043 <= (fillup_transition == 1'b1) ? i_input_data[898 % IN_WIDTH] : pong_storage_data_1043 ^ i_input_data[898 % IN_WIDTH];
                default: pong_storage_data_1043 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1043;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1043 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1043;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1043 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1043;
            end
        end
    end
end

logic ping_storage_data_1044;
logic pong_storage_data_1044;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1044 <= 1'b0;
        pong_storage_data_1044 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                269 / IN_WIDTH: ping_storage_data_1044 <= (fillup_transition == 1'b1) ? i_input_data[269 % IN_WIDTH] : ping_storage_data_1044 ^ i_input_data[269 % IN_WIDTH];
                307 / IN_WIDTH: ping_storage_data_1044 <= (fillup_transition == 1'b1) ? i_input_data[307 % IN_WIDTH] : ping_storage_data_1044 ^ i_input_data[307 % IN_WIDTH];
                813 / IN_WIDTH: ping_storage_data_1044 <= (fillup_transition == 1'b1) ? i_input_data[813 % IN_WIDTH] : ping_storage_data_1044 ^ i_input_data[813 % IN_WIDTH];
                899 / IN_WIDTH: ping_storage_data_1044 <= (fillup_transition == 1'b1) ? i_input_data[899 % IN_WIDTH] : ping_storage_data_1044 ^ i_input_data[899 % IN_WIDTH];
                default: ping_storage_data_1044 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1044;
                endcase
            end else begin
                case (input_count)
                269 / IN_WIDTH: pong_storage_data_1044 <= (fillup_transition == 1'b1) ? i_input_data[269 % IN_WIDTH] : pong_storage_data_1044 ^ i_input_data[269 % IN_WIDTH];
                307 / IN_WIDTH: pong_storage_data_1044 <= (fillup_transition == 1'b1) ? i_input_data[307 % IN_WIDTH] : pong_storage_data_1044 ^ i_input_data[307 % IN_WIDTH];
                813 / IN_WIDTH: pong_storage_data_1044 <= (fillup_transition == 1'b1) ? i_input_data[813 % IN_WIDTH] : pong_storage_data_1044 ^ i_input_data[813 % IN_WIDTH];
                899 / IN_WIDTH: pong_storage_data_1044 <= (fillup_transition == 1'b1) ? i_input_data[899 % IN_WIDTH] : pong_storage_data_1044 ^ i_input_data[899 % IN_WIDTH];
                default: pong_storage_data_1044 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1044;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1044 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1044;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1044 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1044;
            end
        end
    end
end

logic ping_storage_data_1045;
logic pong_storage_data_1045;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1045 <= 1'b0;
        pong_storage_data_1045 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                270 / IN_WIDTH: ping_storage_data_1045 <= (fillup_transition == 1'b1) ? i_input_data[270 % IN_WIDTH] : ping_storage_data_1045 ^ i_input_data[270 % IN_WIDTH];
                308 / IN_WIDTH: ping_storage_data_1045 <= (fillup_transition == 1'b1) ? i_input_data[308 % IN_WIDTH] : ping_storage_data_1045 ^ i_input_data[308 % IN_WIDTH];
                814 / IN_WIDTH: ping_storage_data_1045 <= (fillup_transition == 1'b1) ? i_input_data[814 % IN_WIDTH] : ping_storage_data_1045 ^ i_input_data[814 % IN_WIDTH];
                900 / IN_WIDTH: ping_storage_data_1045 <= (fillup_transition == 1'b1) ? i_input_data[900 % IN_WIDTH] : ping_storage_data_1045 ^ i_input_data[900 % IN_WIDTH];
                default: ping_storage_data_1045 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1045;
                endcase
            end else begin
                case (input_count)
                270 / IN_WIDTH: pong_storage_data_1045 <= (fillup_transition == 1'b1) ? i_input_data[270 % IN_WIDTH] : pong_storage_data_1045 ^ i_input_data[270 % IN_WIDTH];
                308 / IN_WIDTH: pong_storage_data_1045 <= (fillup_transition == 1'b1) ? i_input_data[308 % IN_WIDTH] : pong_storage_data_1045 ^ i_input_data[308 % IN_WIDTH];
                814 / IN_WIDTH: pong_storage_data_1045 <= (fillup_transition == 1'b1) ? i_input_data[814 % IN_WIDTH] : pong_storage_data_1045 ^ i_input_data[814 % IN_WIDTH];
                900 / IN_WIDTH: pong_storage_data_1045 <= (fillup_transition == 1'b1) ? i_input_data[900 % IN_WIDTH] : pong_storage_data_1045 ^ i_input_data[900 % IN_WIDTH];
                default: pong_storage_data_1045 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1045;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1045 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1045;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1045 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1045;
            end
        end
    end
end

logic ping_storage_data_1046;
logic pong_storage_data_1046;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1046 <= 1'b0;
        pong_storage_data_1046 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                271 / IN_WIDTH: ping_storage_data_1046 <= (fillup_transition == 1'b1) ? i_input_data[271 % IN_WIDTH] : ping_storage_data_1046 ^ i_input_data[271 % IN_WIDTH];
                309 / IN_WIDTH: ping_storage_data_1046 <= (fillup_transition == 1'b1) ? i_input_data[309 % IN_WIDTH] : ping_storage_data_1046 ^ i_input_data[309 % IN_WIDTH];
                815 / IN_WIDTH: ping_storage_data_1046 <= (fillup_transition == 1'b1) ? i_input_data[815 % IN_WIDTH] : ping_storage_data_1046 ^ i_input_data[815 % IN_WIDTH];
                901 / IN_WIDTH: ping_storage_data_1046 <= (fillup_transition == 1'b1) ? i_input_data[901 % IN_WIDTH] : ping_storage_data_1046 ^ i_input_data[901 % IN_WIDTH];
                default: ping_storage_data_1046 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1046;
                endcase
            end else begin
                case (input_count)
                271 / IN_WIDTH: pong_storage_data_1046 <= (fillup_transition == 1'b1) ? i_input_data[271 % IN_WIDTH] : pong_storage_data_1046 ^ i_input_data[271 % IN_WIDTH];
                309 / IN_WIDTH: pong_storage_data_1046 <= (fillup_transition == 1'b1) ? i_input_data[309 % IN_WIDTH] : pong_storage_data_1046 ^ i_input_data[309 % IN_WIDTH];
                815 / IN_WIDTH: pong_storage_data_1046 <= (fillup_transition == 1'b1) ? i_input_data[815 % IN_WIDTH] : pong_storage_data_1046 ^ i_input_data[815 % IN_WIDTH];
                901 / IN_WIDTH: pong_storage_data_1046 <= (fillup_transition == 1'b1) ? i_input_data[901 % IN_WIDTH] : pong_storage_data_1046 ^ i_input_data[901 % IN_WIDTH];
                default: pong_storage_data_1046 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1046;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1046 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1046;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1046 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1046;
            end
        end
    end
end

logic ping_storage_data_1047;
logic pong_storage_data_1047;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1047 <= 1'b0;
        pong_storage_data_1047 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                272 / IN_WIDTH: ping_storage_data_1047 <= (fillup_transition == 1'b1) ? i_input_data[272 % IN_WIDTH] : ping_storage_data_1047 ^ i_input_data[272 % IN_WIDTH];
                310 / IN_WIDTH: ping_storage_data_1047 <= (fillup_transition == 1'b1) ? i_input_data[310 % IN_WIDTH] : ping_storage_data_1047 ^ i_input_data[310 % IN_WIDTH];
                816 / IN_WIDTH: ping_storage_data_1047 <= (fillup_transition == 1'b1) ? i_input_data[816 % IN_WIDTH] : ping_storage_data_1047 ^ i_input_data[816 % IN_WIDTH];
                902 / IN_WIDTH: ping_storage_data_1047 <= (fillup_transition == 1'b1) ? i_input_data[902 % IN_WIDTH] : ping_storage_data_1047 ^ i_input_data[902 % IN_WIDTH];
                default: ping_storage_data_1047 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1047;
                endcase
            end else begin
                case (input_count)
                272 / IN_WIDTH: pong_storage_data_1047 <= (fillup_transition == 1'b1) ? i_input_data[272 % IN_WIDTH] : pong_storage_data_1047 ^ i_input_data[272 % IN_WIDTH];
                310 / IN_WIDTH: pong_storage_data_1047 <= (fillup_transition == 1'b1) ? i_input_data[310 % IN_WIDTH] : pong_storage_data_1047 ^ i_input_data[310 % IN_WIDTH];
                816 / IN_WIDTH: pong_storage_data_1047 <= (fillup_transition == 1'b1) ? i_input_data[816 % IN_WIDTH] : pong_storage_data_1047 ^ i_input_data[816 % IN_WIDTH];
                902 / IN_WIDTH: pong_storage_data_1047 <= (fillup_transition == 1'b1) ? i_input_data[902 % IN_WIDTH] : pong_storage_data_1047 ^ i_input_data[902 % IN_WIDTH];
                default: pong_storage_data_1047 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1047;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1047 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1047;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1047 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1047;
            end
        end
    end
end

logic ping_storage_data_1048;
logic pong_storage_data_1048;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1048 <= 1'b0;
        pong_storage_data_1048 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                273 / IN_WIDTH: ping_storage_data_1048 <= (fillup_transition == 1'b1) ? i_input_data[273 % IN_WIDTH] : ping_storage_data_1048 ^ i_input_data[273 % IN_WIDTH];
                311 / IN_WIDTH: ping_storage_data_1048 <= (fillup_transition == 1'b1) ? i_input_data[311 % IN_WIDTH] : ping_storage_data_1048 ^ i_input_data[311 % IN_WIDTH];
                817 / IN_WIDTH: ping_storage_data_1048 <= (fillup_transition == 1'b1) ? i_input_data[817 % IN_WIDTH] : ping_storage_data_1048 ^ i_input_data[817 % IN_WIDTH];
                903 / IN_WIDTH: ping_storage_data_1048 <= (fillup_transition == 1'b1) ? i_input_data[903 % IN_WIDTH] : ping_storage_data_1048 ^ i_input_data[903 % IN_WIDTH];
                default: ping_storage_data_1048 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1048;
                endcase
            end else begin
                case (input_count)
                273 / IN_WIDTH: pong_storage_data_1048 <= (fillup_transition == 1'b1) ? i_input_data[273 % IN_WIDTH] : pong_storage_data_1048 ^ i_input_data[273 % IN_WIDTH];
                311 / IN_WIDTH: pong_storage_data_1048 <= (fillup_transition == 1'b1) ? i_input_data[311 % IN_WIDTH] : pong_storage_data_1048 ^ i_input_data[311 % IN_WIDTH];
                817 / IN_WIDTH: pong_storage_data_1048 <= (fillup_transition == 1'b1) ? i_input_data[817 % IN_WIDTH] : pong_storage_data_1048 ^ i_input_data[817 % IN_WIDTH];
                903 / IN_WIDTH: pong_storage_data_1048 <= (fillup_transition == 1'b1) ? i_input_data[903 % IN_WIDTH] : pong_storage_data_1048 ^ i_input_data[903 % IN_WIDTH];
                default: pong_storage_data_1048 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1048;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1048 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1048;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1048 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1048;
            end
        end
    end
end

logic ping_storage_data_1049;
logic pong_storage_data_1049;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1049 <= 1'b0;
        pong_storage_data_1049 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                274 / IN_WIDTH: ping_storage_data_1049 <= (fillup_transition == 1'b1) ? i_input_data[274 % IN_WIDTH] : ping_storage_data_1049 ^ i_input_data[274 % IN_WIDTH];
                312 / IN_WIDTH: ping_storage_data_1049 <= (fillup_transition == 1'b1) ? i_input_data[312 % IN_WIDTH] : ping_storage_data_1049 ^ i_input_data[312 % IN_WIDTH];
                818 / IN_WIDTH: ping_storage_data_1049 <= (fillup_transition == 1'b1) ? i_input_data[818 % IN_WIDTH] : ping_storage_data_1049 ^ i_input_data[818 % IN_WIDTH];
                904 / IN_WIDTH: ping_storage_data_1049 <= (fillup_transition == 1'b1) ? i_input_data[904 % IN_WIDTH] : ping_storage_data_1049 ^ i_input_data[904 % IN_WIDTH];
                default: ping_storage_data_1049 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1049;
                endcase
            end else begin
                case (input_count)
                274 / IN_WIDTH: pong_storage_data_1049 <= (fillup_transition == 1'b1) ? i_input_data[274 % IN_WIDTH] : pong_storage_data_1049 ^ i_input_data[274 % IN_WIDTH];
                312 / IN_WIDTH: pong_storage_data_1049 <= (fillup_transition == 1'b1) ? i_input_data[312 % IN_WIDTH] : pong_storage_data_1049 ^ i_input_data[312 % IN_WIDTH];
                818 / IN_WIDTH: pong_storage_data_1049 <= (fillup_transition == 1'b1) ? i_input_data[818 % IN_WIDTH] : pong_storage_data_1049 ^ i_input_data[818 % IN_WIDTH];
                904 / IN_WIDTH: pong_storage_data_1049 <= (fillup_transition == 1'b1) ? i_input_data[904 % IN_WIDTH] : pong_storage_data_1049 ^ i_input_data[904 % IN_WIDTH];
                default: pong_storage_data_1049 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1049;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1049 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1049;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1049 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1049;
            end
        end
    end
end

logic ping_storage_data_1050;
logic pong_storage_data_1050;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1050 <= 1'b0;
        pong_storage_data_1050 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                275 / IN_WIDTH: ping_storage_data_1050 <= (fillup_transition == 1'b1) ? i_input_data[275 % IN_WIDTH] : ping_storage_data_1050 ^ i_input_data[275 % IN_WIDTH];
                313 / IN_WIDTH: ping_storage_data_1050 <= (fillup_transition == 1'b1) ? i_input_data[313 % IN_WIDTH] : ping_storage_data_1050 ^ i_input_data[313 % IN_WIDTH];
                819 / IN_WIDTH: ping_storage_data_1050 <= (fillup_transition == 1'b1) ? i_input_data[819 % IN_WIDTH] : ping_storage_data_1050 ^ i_input_data[819 % IN_WIDTH];
                905 / IN_WIDTH: ping_storage_data_1050 <= (fillup_transition == 1'b1) ? i_input_data[905 % IN_WIDTH] : ping_storage_data_1050 ^ i_input_data[905 % IN_WIDTH];
                default: ping_storage_data_1050 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1050;
                endcase
            end else begin
                case (input_count)
                275 / IN_WIDTH: pong_storage_data_1050 <= (fillup_transition == 1'b1) ? i_input_data[275 % IN_WIDTH] : pong_storage_data_1050 ^ i_input_data[275 % IN_WIDTH];
                313 / IN_WIDTH: pong_storage_data_1050 <= (fillup_transition == 1'b1) ? i_input_data[313 % IN_WIDTH] : pong_storage_data_1050 ^ i_input_data[313 % IN_WIDTH];
                819 / IN_WIDTH: pong_storage_data_1050 <= (fillup_transition == 1'b1) ? i_input_data[819 % IN_WIDTH] : pong_storage_data_1050 ^ i_input_data[819 % IN_WIDTH];
                905 / IN_WIDTH: pong_storage_data_1050 <= (fillup_transition == 1'b1) ? i_input_data[905 % IN_WIDTH] : pong_storage_data_1050 ^ i_input_data[905 % IN_WIDTH];
                default: pong_storage_data_1050 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1050;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1050 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1050;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1050 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1050;
            end
        end
    end
end

logic ping_storage_data_1051;
logic pong_storage_data_1051;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1051 <= 1'b0;
        pong_storage_data_1051 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                276 / IN_WIDTH: ping_storage_data_1051 <= (fillup_transition == 1'b1) ? i_input_data[276 % IN_WIDTH] : ping_storage_data_1051 ^ i_input_data[276 % IN_WIDTH];
                314 / IN_WIDTH: ping_storage_data_1051 <= (fillup_transition == 1'b1) ? i_input_data[314 % IN_WIDTH] : ping_storage_data_1051 ^ i_input_data[314 % IN_WIDTH];
                820 / IN_WIDTH: ping_storage_data_1051 <= (fillup_transition == 1'b1) ? i_input_data[820 % IN_WIDTH] : ping_storage_data_1051 ^ i_input_data[820 % IN_WIDTH];
                906 / IN_WIDTH: ping_storage_data_1051 <= (fillup_transition == 1'b1) ? i_input_data[906 % IN_WIDTH] : ping_storage_data_1051 ^ i_input_data[906 % IN_WIDTH];
                default: ping_storage_data_1051 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1051;
                endcase
            end else begin
                case (input_count)
                276 / IN_WIDTH: pong_storage_data_1051 <= (fillup_transition == 1'b1) ? i_input_data[276 % IN_WIDTH] : pong_storage_data_1051 ^ i_input_data[276 % IN_WIDTH];
                314 / IN_WIDTH: pong_storage_data_1051 <= (fillup_transition == 1'b1) ? i_input_data[314 % IN_WIDTH] : pong_storage_data_1051 ^ i_input_data[314 % IN_WIDTH];
                820 / IN_WIDTH: pong_storage_data_1051 <= (fillup_transition == 1'b1) ? i_input_data[820 % IN_WIDTH] : pong_storage_data_1051 ^ i_input_data[820 % IN_WIDTH];
                906 / IN_WIDTH: pong_storage_data_1051 <= (fillup_transition == 1'b1) ? i_input_data[906 % IN_WIDTH] : pong_storage_data_1051 ^ i_input_data[906 % IN_WIDTH];
                default: pong_storage_data_1051 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1051;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1051 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1051;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1051 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1051;
            end
        end
    end
end

logic ping_storage_data_1052;
logic pong_storage_data_1052;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1052 <= 1'b0;
        pong_storage_data_1052 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                277 / IN_WIDTH: ping_storage_data_1052 <= (fillup_transition == 1'b1) ? i_input_data[277 % IN_WIDTH] : ping_storage_data_1052 ^ i_input_data[277 % IN_WIDTH];
                315 / IN_WIDTH: ping_storage_data_1052 <= (fillup_transition == 1'b1) ? i_input_data[315 % IN_WIDTH] : ping_storage_data_1052 ^ i_input_data[315 % IN_WIDTH];
                821 / IN_WIDTH: ping_storage_data_1052 <= (fillup_transition == 1'b1) ? i_input_data[821 % IN_WIDTH] : ping_storage_data_1052 ^ i_input_data[821 % IN_WIDTH];
                907 / IN_WIDTH: ping_storage_data_1052 <= (fillup_transition == 1'b1) ? i_input_data[907 % IN_WIDTH] : ping_storage_data_1052 ^ i_input_data[907 % IN_WIDTH];
                default: ping_storage_data_1052 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1052;
                endcase
            end else begin
                case (input_count)
                277 / IN_WIDTH: pong_storage_data_1052 <= (fillup_transition == 1'b1) ? i_input_data[277 % IN_WIDTH] : pong_storage_data_1052 ^ i_input_data[277 % IN_WIDTH];
                315 / IN_WIDTH: pong_storage_data_1052 <= (fillup_transition == 1'b1) ? i_input_data[315 % IN_WIDTH] : pong_storage_data_1052 ^ i_input_data[315 % IN_WIDTH];
                821 / IN_WIDTH: pong_storage_data_1052 <= (fillup_transition == 1'b1) ? i_input_data[821 % IN_WIDTH] : pong_storage_data_1052 ^ i_input_data[821 % IN_WIDTH];
                907 / IN_WIDTH: pong_storage_data_1052 <= (fillup_transition == 1'b1) ? i_input_data[907 % IN_WIDTH] : pong_storage_data_1052 ^ i_input_data[907 % IN_WIDTH];
                default: pong_storage_data_1052 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1052;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1052 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1052;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1052 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1052;
            end
        end
    end
end

logic ping_storage_data_1053;
logic pong_storage_data_1053;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1053 <= 1'b0;
        pong_storage_data_1053 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                278 / IN_WIDTH: ping_storage_data_1053 <= (fillup_transition == 1'b1) ? i_input_data[278 % IN_WIDTH] : ping_storage_data_1053 ^ i_input_data[278 % IN_WIDTH];
                316 / IN_WIDTH: ping_storage_data_1053 <= (fillup_transition == 1'b1) ? i_input_data[316 % IN_WIDTH] : ping_storage_data_1053 ^ i_input_data[316 % IN_WIDTH];
                822 / IN_WIDTH: ping_storage_data_1053 <= (fillup_transition == 1'b1) ? i_input_data[822 % IN_WIDTH] : ping_storage_data_1053 ^ i_input_data[822 % IN_WIDTH];
                908 / IN_WIDTH: ping_storage_data_1053 <= (fillup_transition == 1'b1) ? i_input_data[908 % IN_WIDTH] : ping_storage_data_1053 ^ i_input_data[908 % IN_WIDTH];
                default: ping_storage_data_1053 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1053;
                endcase
            end else begin
                case (input_count)
                278 / IN_WIDTH: pong_storage_data_1053 <= (fillup_transition == 1'b1) ? i_input_data[278 % IN_WIDTH] : pong_storage_data_1053 ^ i_input_data[278 % IN_WIDTH];
                316 / IN_WIDTH: pong_storage_data_1053 <= (fillup_transition == 1'b1) ? i_input_data[316 % IN_WIDTH] : pong_storage_data_1053 ^ i_input_data[316 % IN_WIDTH];
                822 / IN_WIDTH: pong_storage_data_1053 <= (fillup_transition == 1'b1) ? i_input_data[822 % IN_WIDTH] : pong_storage_data_1053 ^ i_input_data[822 % IN_WIDTH];
                908 / IN_WIDTH: pong_storage_data_1053 <= (fillup_transition == 1'b1) ? i_input_data[908 % IN_WIDTH] : pong_storage_data_1053 ^ i_input_data[908 % IN_WIDTH];
                default: pong_storage_data_1053 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1053;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1053 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1053;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1053 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1053;
            end
        end
    end
end

logic ping_storage_data_1054;
logic pong_storage_data_1054;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1054 <= 1'b0;
        pong_storage_data_1054 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                279 / IN_WIDTH: ping_storage_data_1054 <= (fillup_transition == 1'b1) ? i_input_data[279 % IN_WIDTH] : ping_storage_data_1054 ^ i_input_data[279 % IN_WIDTH];
                317 / IN_WIDTH: ping_storage_data_1054 <= (fillup_transition == 1'b1) ? i_input_data[317 % IN_WIDTH] : ping_storage_data_1054 ^ i_input_data[317 % IN_WIDTH];
                823 / IN_WIDTH: ping_storage_data_1054 <= (fillup_transition == 1'b1) ? i_input_data[823 % IN_WIDTH] : ping_storage_data_1054 ^ i_input_data[823 % IN_WIDTH];
                909 / IN_WIDTH: ping_storage_data_1054 <= (fillup_transition == 1'b1) ? i_input_data[909 % IN_WIDTH] : ping_storage_data_1054 ^ i_input_data[909 % IN_WIDTH];
                default: ping_storage_data_1054 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1054;
                endcase
            end else begin
                case (input_count)
                279 / IN_WIDTH: pong_storage_data_1054 <= (fillup_transition == 1'b1) ? i_input_data[279 % IN_WIDTH] : pong_storage_data_1054 ^ i_input_data[279 % IN_WIDTH];
                317 / IN_WIDTH: pong_storage_data_1054 <= (fillup_transition == 1'b1) ? i_input_data[317 % IN_WIDTH] : pong_storage_data_1054 ^ i_input_data[317 % IN_WIDTH];
                823 / IN_WIDTH: pong_storage_data_1054 <= (fillup_transition == 1'b1) ? i_input_data[823 % IN_WIDTH] : pong_storage_data_1054 ^ i_input_data[823 % IN_WIDTH];
                909 / IN_WIDTH: pong_storage_data_1054 <= (fillup_transition == 1'b1) ? i_input_data[909 % IN_WIDTH] : pong_storage_data_1054 ^ i_input_data[909 % IN_WIDTH];
                default: pong_storage_data_1054 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1054;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1054 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1054;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1054 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1054;
            end
        end
    end
end

logic ping_storage_data_1055;
logic pong_storage_data_1055;

always_ff @ (posedge i_clock) begin
    if (i_reset == 1'b1) begin
        ping_storage_data_1055 <= 1'b0;
        pong_storage_data_1055 <= 1'b0;
    end else begin
        if ((i_input_valid & o_input_ready) == 1'b1) begin
            if (fillup_state == ST_PING) begin
                case (input_count)
                280 / IN_WIDTH: ping_storage_data_1055 <= (fillup_transition == 1'b1) ? i_input_data[280 % IN_WIDTH] : ping_storage_data_1055 ^ i_input_data[280 % IN_WIDTH];
                318 / IN_WIDTH: ping_storage_data_1055 <= (fillup_transition == 1'b1) ? i_input_data[318 % IN_WIDTH] : ping_storage_data_1055 ^ i_input_data[318 % IN_WIDTH];
                824 / IN_WIDTH: ping_storage_data_1055 <= (fillup_transition == 1'b1) ? i_input_data[824 % IN_WIDTH] : ping_storage_data_1055 ^ i_input_data[824 % IN_WIDTH];
                910 / IN_WIDTH: ping_storage_data_1055 <= (fillup_transition == 1'b1) ? i_input_data[910 % IN_WIDTH] : ping_storage_data_1055 ^ i_input_data[910 % IN_WIDTH];
                default: ping_storage_data_1055 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1055;
                endcase
            end else begin
                case (input_count)
                280 / IN_WIDTH: pong_storage_data_1055 <= (fillup_transition == 1'b1) ? i_input_data[280 % IN_WIDTH] : pong_storage_data_1055 ^ i_input_data[280 % IN_WIDTH];
                318 / IN_WIDTH: pong_storage_data_1055 <= (fillup_transition == 1'b1) ? i_input_data[318 % IN_WIDTH] : pong_storage_data_1055 ^ i_input_data[318 % IN_WIDTH];
                824 / IN_WIDTH: pong_storage_data_1055 <= (fillup_transition == 1'b1) ? i_input_data[824 % IN_WIDTH] : pong_storage_data_1055 ^ i_input_data[824 % IN_WIDTH];
                910 / IN_WIDTH: pong_storage_data_1055 <= (fillup_transition == 1'b1) ? i_input_data[910 % IN_WIDTH] : pong_storage_data_1055 ^ i_input_data[910 % IN_WIDTH];
                default: pong_storage_data_1055 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1055;
                endcase
            end
        end else begin
            if ((fillup_state == ST_PING)) begin
                ping_storage_data_1055 <= (fillup_transition == 1'b1) ? 1'b0 : ping_storage_data_1055;
            end
            if ((fillup_state == ST_PONG) && (fillup_transition == 1'b1)) begin
                pong_storage_data_1055 <= (fillup_transition == 1'b1) ? 1'b0 : pong_storage_data_1055;
            end
        end
    end
end


endmodule: sparse_mult_by_A

`default_nettype wire
