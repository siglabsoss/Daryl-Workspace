`timescale 10ps / 10ps

`default_nettype none

module chmod_dds (
    input  wire logic [32-1:0] i_phase_inc,
    input  wire logic          i_phase_inc_valid,
    output      logic [36-1:0] o_cosine_data,
    output      logic [36-1:0] o_sine_data,
    input       logic          i_ready,
    input  wire logic          i_clock,
    input  wire logic          i_reset
);

// Phase increment
logic [32-1:0] phase_inc_reg;
logic [32-1:0] phase_accum;

always_ff @ (posedge i_clock) begin
    // Read input phase increment
    if (i_phase_inc_valid == 1'b1) begin
        phase_inc_reg <= i_phase_inc;
    end
    // Increment phase whenever an output is requested
    if (i_reset == 1'b1) begin
        phase_accum <= '0;
    end else if (i_ready == 1'b1) begin
        phase_accum <= phase_accum + phase_inc_reg;
    end
end

// Sine/Cosine Look Up Table
localparam integer WIDTH = 36;
localparam integer RESIDUAL_WIDTH = WIDTH-12;

logic signed [WIDTH-1:0]      cosine_reg0 /* synthesis syn_ramstyle="block_ram" */;
logic signed [WIDTH-1:0]      sine_reg0 /* synthesis syn_ramstyle="block_ram" */;
// logic [16+RESIDUAL_WIDTH-1:0] residual_reg0;

// Pipeline Stage 0
always_ff @ (posedge i_clock) begin
    if (i_ready == 1'b1) begin
        // Perform table look up
        case(phase_accum[32-1:32-12])
        0: begin
            cosine_reg0 <= 36'sb11111111111111111111111111111111111;
            sine_reg0   <= 36'sb0;
        end
        1: begin
            cosine_reg0 <= 36'sb11111111111111111110110001000010101;
            sine_reg0   <= 36'sb11001001000011111101010110;
        end
        2: begin
            cosine_reg0 <= 36'sb11111111111111111011000100001011000;
            sine_reg0   <= 36'sb110010010000111111000110000;
        end
        3: begin
            cosine_reg0 <= 36'sb11111111111111110100111001011000111;
            sine_reg0   <= 36'sb1001011011001011110000010001;
        end
        4: begin
            cosine_reg0 <= 36'sb11111111111111101100010000101100011;
            sine_reg0   <= 36'sb1100100100001111100001111111;
        end
        5: begin
            cosine_reg0 <= 36'sb11111111111111100001001010000101100;
            sine_reg0   <= 36'sb1111101101010011001011111101;
        end
        6: begin
            cosine_reg0 <= 36'sb11111111111111010011100101100100101;
            sine_reg0   <= 36'sb10010110110010110101100001110;
        end
        7: begin
            cosine_reg0 <= 36'sb11111111111111000011100011001001101;
            sine_reg0   <= 36'sb10101111111011010000000111000;
        end
        8: begin
            cosine_reg0 <= 36'sb11111111111110110001000010110100110;
            sine_reg0   <= 36'sb11001001000011101000111111101;
        end
        9: begin
            cosine_reg0 <= 36'sb11111111111110011100000100100110001;
            sine_reg0   <= 36'sb11100010001011111111111100010;
        end
        10: begin
            cosine_reg0 <= 36'sb11111111111110000100101000011110000;
            sine_reg0   <= 36'sb11111011010100010100101101011;
        end
        11: begin
            cosine_reg0 <= 36'sb11111111111101101010101110011100101;
            sine_reg0   <= 36'sb100010100011100100111000011011;
        end
        12: begin
            cosine_reg0 <= 36'sb11111111111101001110010110100010010;
            sine_reg0   <= 36'sb100101101100100110110101111000;
        end
        13: begin
            cosine_reg0 <= 36'sb11111111111100101111100000101111000;
            sine_reg0   <= 36'sb101000110101101000011100000100;
        end
        14: begin
            cosine_reg0 <= 36'sb11111111111100001110001101000011011;
            sine_reg0   <= 36'sb101011111110101001101001000100;
        end
        15: begin
            cosine_reg0 <= 36'sb11111111111011101010011011011111101;
            sine_reg0   <= 36'sb101111000111101010011010111100;
        end
        16: begin
            cosine_reg0 <= 36'sb11111111111011000100001100000100000;
            sine_reg0   <= 36'sb110010010000101010101111101111;
        end
        17: begin
            cosine_reg0 <= 36'sb11111111111010011011011110110001000;
            sine_reg0   <= 36'sb110101011001101010100101100011;
        end
        18: begin
            cosine_reg0 <= 36'sb11111111111001110000010011100111000;
            sine_reg0   <= 36'sb111000100010101001111010011010;
        end
        19: begin
            cosine_reg0 <= 36'sb11111111111001000010101010100110010;
            sine_reg0   <= 36'sb111011101011101000101100011001;
        end
        20: begin
            cosine_reg0 <= 36'sb11111111111000010010100011101111011;
            sine_reg0   <= 36'sb111110110100100110111001100100;
        end
        21: begin
            cosine_reg0 <= 36'sb11111111110111011111111111000010111;
            sine_reg0   <= 36'sb1000001111101100100011111111110;
        end
        22: begin
            cosine_reg0 <= 36'sb11111111110110101010111100100001000;
            sine_reg0   <= 36'sb1000101000110100001011101101101;
        end
        23: begin
            cosine_reg0 <= 36'sb11111111110101110011011100001010100;
            sine_reg0   <= 36'sb1001000001111011101110000110100;
        end
        24: begin
            cosine_reg0 <= 36'sb11111111110100111001011101111111111;
            sine_reg0   <= 36'sb1001011011000011001010111010110;
        end
        25: begin
            cosine_reg0 <= 36'sb11111111110011111101000010000001100;
            sine_reg0   <= 36'sb1001110100001010100001111011001;
        end
        26: begin
            cosine_reg0 <= 36'sb11111111110010111110001000010000001;
            sine_reg0   <= 36'sb1010001101010001110010111000000;
        end
        27: begin
            cosine_reg0 <= 36'sb11111111110001111100110000101100011;
            sine_reg0   <= 36'sb1010100110011000111101100001111;
        end
        28: begin
            cosine_reg0 <= 36'sb11111111110000111000111011010110110;
            sine_reg0   <= 36'sb1010111111100000000001101001010;
        end
        29: begin
            cosine_reg0 <= 36'sb11111111101111110010101000010000000;
            sine_reg0   <= 36'sb1011011000100110111110111110110;
        end
        30: begin
            cosine_reg0 <= 36'sb11111111101110101001110111011000110;
            sine_reg0   <= 36'sb1011110001101101110101010010110;
        end
        31: begin
            cosine_reg0 <= 36'sb11111111101101011110101000110001110;
            sine_reg0   <= 36'sb1100001010110100100100010101111;
        end
        32: begin
            cosine_reg0 <= 36'sb11111111101100010000111100011011101;
            sine_reg0   <= 36'sb1100100011111011001011111000100;
        end
        33: begin
            cosine_reg0 <= 36'sb11111111101011000000110010010111011;
            sine_reg0   <= 36'sb1100111101000001101011101011010;
        end
        34: begin
            cosine_reg0 <= 36'sb11111111101001101110001010100101011;
            sine_reg0   <= 36'sb1101010110001000000011011110101;
        end
        35: begin
            cosine_reg0 <= 36'sb11111111101000011001000101000110111;
            sine_reg0   <= 36'sb1101101111001110010011000011010;
        end
        36: begin
            cosine_reg0 <= 36'sb11111111100111000001100001111100010;
            sine_reg0   <= 36'sb1110001000010100011010001001011;
        end
        37: begin
            cosine_reg0 <= 36'sb11111111100101100111100001000110110;
            sine_reg0   <= 36'sb1110100001011010011000100001110;
        end
        38: begin
            cosine_reg0 <= 36'sb11111111100100001011000010100110111;
            sine_reg0   <= 36'sb1110111010100000001101111100110;
        end
        39: begin
            cosine_reg0 <= 36'sb11111111100010101100000110011101111;
            sine_reg0   <= 36'sb1111010011100101111010001011000;
        end
        40: begin
            cosine_reg0 <= 36'sb11111111100001001010101100101100011;
            sine_reg0   <= 36'sb1111101100101011011100111101000;
        end
        41: begin
            cosine_reg0 <= 36'sb11111111011111100110110101010011011;
            sine_reg0   <= 36'sb10000000101110000110110000011010;
        end
        42: begin
            cosine_reg0 <= 36'sb11111111011110000000100000010100000;
            sine_reg0   <= 36'sb10000011110110110000101001110010;
        end
        43: begin
            cosine_reg0 <= 36'sb11111111011100010111101101101111000;
            sine_reg0   <= 36'sb10000110111111011001010001110101;
        end
        44: begin
            cosine_reg0 <= 36'sb11111111011010101100011101100101101;
            sine_reg0   <= 36'sb10001010001000000000100110100111;
        end
        45: begin
            cosine_reg0 <= 36'sb11111111011000111110101111111000101;
            sine_reg0   <= 36'sb10001101010000100110100110001011;
        end
        46: begin
            cosine_reg0 <= 36'sb11111111010111001110100100101001011;
            sine_reg0   <= 36'sb10010000011001001011001110100111;
        end
        47: begin
            cosine_reg0 <= 36'sb11111111010101011011111011111000110;
            sine_reg0   <= 36'sb10010011100001101110011101111111;
        end
        48: begin
            cosine_reg0 <= 36'sb11111111010011100110110101100111111;
            sine_reg0   <= 36'sb10010110101010010000010010010110;
        end
        49: begin
            cosine_reg0 <= 36'sb11111111010001101111010001111000000;
            sine_reg0   <= 36'sb10011001110010110000101001110010;
        end
        50: begin
            cosine_reg0 <= 36'sb11111111001111110101010000101010001;
            sine_reg0   <= 36'sb10011100111011001111100010010110;
        end
        51: begin
            cosine_reg0 <= 36'sb11111111001101111000110001111111100;
            sine_reg0   <= 36'sb10100000000011101100111010000111;
        end
        52: begin
            cosine_reg0 <= 36'sb11111111001011111001110101111001011;
            sine_reg0   <= 36'sb10100011001100001000101111001001;
        end
        53: begin
            cosine_reg0 <= 36'sb11111111001001111000011100011000110;
            sine_reg0   <= 36'sb10100110010100100010111111100001;
        end
        54: begin
            cosine_reg0 <= 36'sb11111111000111110100100101011111001;
            sine_reg0   <= 36'sb10101001011100111011101001010010;
        end
        55: begin
            cosine_reg0 <= 36'sb11111111000101101110010001001101110;
            sine_reg0   <= 36'sb10101100100101010010101010100010;
        end
        56: begin
            cosine_reg0 <= 36'sb11111111000011100101011111100101110;
            sine_reg0   <= 36'sb10101111101101101000000001010101;
        end
        57: begin
            cosine_reg0 <= 36'sb11111111000001011010010000101000101;
            sine_reg0   <= 36'sb10110010110101111011101011101110;
        end
        58: begin
            cosine_reg0 <= 36'sb11111110111111001100100100010111101;
            sine_reg0   <= 36'sb10110101111110001101100111110100;
        end
        59: begin
            cosine_reg0 <= 36'sb11111110111100111100011010110100001;
            sine_reg0   <= 36'sb10111001000110011101110011101001;
        end
        60: begin
            cosine_reg0 <= 36'sb11111110111010101001110011111111011;
            sine_reg0   <= 36'sb10111100001110101100001101010011;
        end
        61: begin
            cosine_reg0 <= 36'sb11111110111000010100101111111011001;
            sine_reg0   <= 36'sb10111111010110111000110010110110;
        end
        62: begin
            cosine_reg0 <= 36'sb11111110110101111101001110101000100;
            sine_reg0   <= 36'sb11000010011111000011100010010110;
        end
        63: begin
            cosine_reg0 <= 36'sb11111110110011100011010000001001001;
            sine_reg0   <= 36'sb11000101100111001100011001111000;
        end
        64: begin
            cosine_reg0 <= 36'sb11111110110001000110110100011110011;
            sine_reg0   <= 36'sb11001000101111010011010111100001;
        end
        65: begin
            cosine_reg0 <= 36'sb11111110101110100111111011101001111;
            sine_reg0   <= 36'sb11001011110111011000011001010101;
        end
        66: begin
            cosine_reg0 <= 36'sb11111110101100000110100101101101001;
            sine_reg0   <= 36'sb11001110111111011011011101011001;
        end
        67: begin
            cosine_reg0 <= 36'sb11111110101001100010110010101001101;
            sine_reg0   <= 36'sb11010010000111011100100001110001;
        end
        68: begin
            cosine_reg0 <= 36'sb11111110100110111100100010100001000;
            sine_reg0   <= 36'sb11010101001111011011100100100010;
        end
        69: begin
            cosine_reg0 <= 36'sb11111110100100010011110101010100110;
            sine_reg0   <= 36'sb11011000010111011000100011110001;
        end
        70: begin
            cosine_reg0 <= 36'sb11111110100001101000101011000110101;
            sine_reg0   <= 36'sb11011011011111010011011101100010;
        end
        71: begin
            cosine_reg0 <= 36'sb11111110011110111011000011111000010;
            sine_reg0   <= 36'sb11011110100111001100001111111001;
        end
        72: begin
            cosine_reg0 <= 36'sb11111110011100001010111111101011010;
            sine_reg0   <= 36'sb11100001101111000010111000111101;
        end
        73: begin
            cosine_reg0 <= 36'sb11111110011001011000011110100001100;
            sine_reg0   <= 36'sb11100100110110110111010110110001;
        end
        74: begin
            cosine_reg0 <= 36'sb11111110010110100011100000011100011;
            sine_reg0   <= 36'sb11100111111110101001100111011001;
        end
        75: begin
            cosine_reg0 <= 36'sb11111110010011101100000101011110000;
            sine_reg0   <= 36'sb11101011000110011001101000111100;
        end
        76: begin
            cosine_reg0 <= 36'sb11111110010000110010001101100111111;
            sine_reg0   <= 36'sb11101110001110000111011001011101;
        end
        77: begin
            cosine_reg0 <= 36'sb11111110001101110101111000111011111;
            sine_reg0   <= 36'sb11110001010101110010110111000010;
        end
        78: begin
            cosine_reg0 <= 36'sb11111110001010110111000111011011110;
            sine_reg0   <= 36'sb11110100011101011011111111101111;
        end
        79: begin
            cosine_reg0 <= 36'sb11111110000111110101111001001001100;
            sine_reg0   <= 36'sb11110111100101000010110001101001;
        end
        80: begin
            cosine_reg0 <= 36'sb11111110000100110010001110000110111;
            sine_reg0   <= 36'sb11111010101100100111001010110101;
        end
        81: begin
            cosine_reg0 <= 36'sb11111110000001101100000110010101111;
            sine_reg0   <= 36'sb11111101110100001001001001011000;
        end
        82: begin
            cosine_reg0 <= 36'sb11111101111110100011100001111000010;
            sine_reg0   <= 36'sb100000000111011101000101011010111;
        end
        83: begin
            cosine_reg0 <= 36'sb11111101111011011000100000110000000;
            sine_reg0   <= 36'sb100000100000011000101101110110110;
        end
        84: begin
            cosine_reg0 <= 36'sb11111101111000001011000010111111000;
            sine_reg0   <= 36'sb100000111001010100000010001111100;
        end
        85: begin
            cosine_reg0 <= 36'sb11111101110100111011001000100111011;
            sine_reg0   <= 36'sb100001010010001111000010010101011;
        end
        86: begin
            cosine_reg0 <= 36'sb11111101110001101000110001101011001;
            sine_reg0   <= 36'sb100001101011001001101101111001011;
        end
        87: begin
            cosine_reg0 <= 36'sb11111101101110010011111110001100001;
            sine_reg0   <= 36'sb100010000100000100000100101011111;
        end
        88: begin
            cosine_reg0 <= 36'sb11111101101010111100101110001100100;
            sine_reg0   <= 36'sb100010011100111110000110011101110;
        end
        89: begin
            cosine_reg0 <= 36'sb11111101100111100011000001101110100;
            sine_reg0   <= 36'sb100010110101110111110010111111011;
        end
        90: begin
            cosine_reg0 <= 36'sb11111101100100000110111000110011111;
            sine_reg0   <= 36'sb100011001110110001001010000001100;
        end
        91: begin
            cosine_reg0 <= 36'sb11111101100000101000010011011111001;
            sine_reg0   <= 36'sb100011100111101010001011010100110;
        end
        92: begin
            cosine_reg0 <= 36'sb11111101011101000111010001110010001;
            sine_reg0   <= 36'sb100100000000100010110110101001111;
        end
        93: begin
            cosine_reg0 <= 36'sb11111101011001100011110011101111001;
            sine_reg0   <= 36'sb100100011001011011001011110001011;
        end
        94: begin
            cosine_reg0 <= 36'sb11111101010101111101111001011000010;
            sine_reg0   <= 36'sb100100110010010011001010011100000;
        end
        95: begin
            cosine_reg0 <= 36'sb11111101010010010101100010101111111;
            sine_reg0   <= 36'sb100101001011001010110010011010011;
        end
        96: begin
            cosine_reg0 <= 36'sb11111101001110101010101111111000001;
            sine_reg0   <= 36'sb100101100100000010000011011101001;
        end
        97: begin
            cosine_reg0 <= 36'sb11111101001010111101100000110011011;
            sine_reg0   <= 36'sb100101111100111000111101010101000;
        end
        98: begin
            cosine_reg0 <= 36'sb11111101000111001101110101100011110;
            sine_reg0   <= 36'sb100110010101101111011111110010100;
        end
        99: begin
            cosine_reg0 <= 36'sb11111101000011011011101110001011101;
            sine_reg0   <= 36'sb100110101110100101101010100110100;
        end
        100: begin
            cosine_reg0 <= 36'sb11111100111111100111001010101101010;
            sine_reg0   <= 36'sb100111000111011011011101100001101;
        end
        101: begin
            cosine_reg0 <= 36'sb11111100111011110000001011001011010;
            sine_reg0   <= 36'sb100111100000010000111000010100011;
        end
        102: begin
            cosine_reg0 <= 36'sb11111100110111110110101111100111110;
            sine_reg0   <= 36'sb100111111001000101111010101111110;
        end
        103: begin
            cosine_reg0 <= 36'sb11111100110011111010111000000101010;
            sine_reg0   <= 36'sb101000010001111010100100100100001;
        end
        104: begin
            cosine_reg0 <= 36'sb11111100101111111100100100100110001;
            sine_reg0   <= 36'sb101000101010101110110101100010010;
        end
        105: begin
            cosine_reg0 <= 36'sb11111100101011111011110101001100111;
            sine_reg0   <= 36'sb101001000011100010101101011011000;
        end
        106: begin
            cosine_reg0 <= 36'sb11111100100111111000101001111100000;
            sine_reg0   <= 36'sb101001011100010110001011111110111;
        end
        107: begin
            cosine_reg0 <= 36'sb11111100100011110011000010110110000;
            sine_reg0   <= 36'sb101001110101001001010000111110110;
        end
        108: begin
            cosine_reg0 <= 36'sb11111100011111101010111111111101011;
            sine_reg0   <= 36'sb101010001101111011111100001011001;
        end
        109: begin
            cosine_reg0 <= 36'sb11111100011011100000100001010100100;
            sine_reg0   <= 36'sb101010100110101110001101010100111;
        end
        110: begin
            cosine_reg0 <= 36'sb11111100010111010011100110111110010;
            sine_reg0   <= 36'sb101010111111100000000100001100101;
        end
        111: begin
            cosine_reg0 <= 36'sb11111100010011000100010000111101000;
            sine_reg0   <= 36'sb101011011000010001100000100011001;
        end
        112: begin
            cosine_reg0 <= 36'sb11111100001110110010011111010011011;
            sine_reg0   <= 36'sb101011110001000010100010001001001;
        end
        113: begin
            cosine_reg0 <= 36'sb11111100001010011110010010000100001;
            sine_reg0   <= 36'sb101100001001110011001000101111001;
        end
        114: begin
            cosine_reg0 <= 36'sb11111100000110000111101001010001111;
            sine_reg0   <= 36'sb101100100010100011010100000110010;
        end
        115: begin
            cosine_reg0 <= 36'sb11111100000001101110100100111111010;
            sine_reg0   <= 36'sb101100111011010011000011111110111;
        end
        116: begin
            cosine_reg0 <= 36'sb11111011111101010011000101001111001;
            sine_reg0   <= 36'sb101101010100000010011000001001111;
        end
        117: begin
            cosine_reg0 <= 36'sb11111011111000110101001010000100000;
            sine_reg0   <= 36'sb101101101100110001010000011000000;
        end
        118: begin
            cosine_reg0 <= 36'sb11111011110100010100110011100000110;
            sine_reg0   <= 36'sb101110000101011111101100011010000;
        end
        119: begin
            cosine_reg0 <= 36'sb11111011101111110010000001101000001;
            sine_reg0   <= 36'sb101110011110001101101100000000101;
        end
        120: begin
            cosine_reg0 <= 36'sb11111011101011001100110100011100111;
            sine_reg0   <= 36'sb101110110110111011001110111100101;
        end
        121: begin
            cosine_reg0 <= 36'sb11111011100110100101001100000010000;
            sine_reg0   <= 36'sb101111001111101000010100111110101;
        end
        122: begin
            cosine_reg0 <= 36'sb11111011100001111011001000011010010;
            sine_reg0   <= 36'sb101111101000010100111101110111101;
        end
        123: begin
            cosine_reg0 <= 36'sb11111011011101001110101001101000100;
            sine_reg0   <= 36'sb110000000001000001001001011000010;
        end
        124: begin
            cosine_reg0 <= 36'sb11111011011000011111101111101111100;
            sine_reg0   <= 36'sb110000011001101100110111010001010;
        end
        125: begin
            cosine_reg0 <= 36'sb11111011010011101110011010110010100;
            sine_reg0   <= 36'sb110000110010011000000111010011011;
        end
        126: begin
            cosine_reg0 <= 36'sb11111011001110111010101010110100001;
            sine_reg0   <= 36'sb110001001011000010111001001111100;
        end
        127: begin
            cosine_reg0 <= 36'sb11111011001010000100011111110111100;
            sine_reg0   <= 36'sb110001100011101101001100110110011;
        end
        128: begin
            cosine_reg0 <= 36'sb11111011000101001011111001111111101;
            sine_reg0   <= 36'sb110001111100010111000001111000110;
        end
        129: begin
            cosine_reg0 <= 36'sb11111011000000010000111001001111011;
            sine_reg0   <= 36'sb110010010101000000011000000111100;
        end
        130: begin
            cosine_reg0 <= 36'sb11111010111011010011011101101010000;
            sine_reg0   <= 36'sb110010101101101001001111010011011;
        end
        131: begin
            cosine_reg0 <= 36'sb11111010110110010011100111010010011;
            sine_reg0   <= 36'sb110011000110010001100111001101001;
        end
        132: begin
            cosine_reg0 <= 36'sb11111010110001010001010110001011101;
            sine_reg0   <= 36'sb110011011110111001011111100101110;
        end
        133: begin
            cosine_reg0 <= 36'sb11111010101100001100101010011000111;
            sine_reg0   <= 36'sb110011110111100000111000001101110;
        end
        134: begin
            cosine_reg0 <= 36'sb11111010100111000101100011111101011;
            sine_reg0   <= 36'sb110100010000000111110000110110001;
        end
        135: begin
            cosine_reg0 <= 36'sb11111010100001111100000010111100000;
            sine_reg0   <= 36'sb110100101000101110001001001111110;
        end
        136: begin
            cosine_reg0 <= 36'sb11111010011100110000000111011000010;
            sine_reg0   <= 36'sb110101000001010100000001001011011;
        end
        137: begin
            cosine_reg0 <= 36'sb11111010010111100001110001010101000;
            sine_reg0   <= 36'sb110101011001111001011000011001110;
        end
        138: begin
            cosine_reg0 <= 36'sb11111010010010010001000000110101110;
            sine_reg0   <= 36'sb110101110010011110001110101011111;
        end
        139: begin
            cosine_reg0 <= 36'sb11111010001100111101110101111101101;
            sine_reg0   <= 36'sb110110001011000010100011110010100;
        end
        140: begin
            cosine_reg0 <= 36'sb11111010000111101000010000101111111;
            sine_reg0   <= 36'sb110110100011100110010111011110100;
        end
        141: begin
            cosine_reg0 <= 36'sb11111010000010010000010001001111110;
            sine_reg0   <= 36'sb110110111100001001101001100000101;
        end
        142: begin
            cosine_reg0 <= 36'sb11111001111100110101110111100000110;
            sine_reg0   <= 36'sb110111010100101100011001101001111;
        end
        143: begin
            cosine_reg0 <= 36'sb11111001110111011001000011100110000;
            sine_reg0   <= 36'sb110111101101001110100111101011000;
        end
        144: begin
            cosine_reg0 <= 36'sb11111001110001111001110101100011000;
            sine_reg0   <= 36'sb111000000101110000010011010101000;
        end
        145: begin
            cosine_reg0 <= 36'sb11111001101100011000001101011011001;
            sine_reg0   <= 36'sb111000011110010001011100011000101;
        end
        146: begin
            cosine_reg0 <= 36'sb11111001100110110100001011010001110;
            sine_reg0   <= 36'sb111000110110110010000010100110110;
        end
        147: begin
            cosine_reg0 <= 36'sb11111001100001001101101111001010010;
            sine_reg0   <= 36'sb111001001111010010000101110000010;
        end
        148: begin
            cosine_reg0 <= 36'sb11111001011011100100111001001000001;
            sine_reg0   <= 36'sb111001100111110001100101100110001;
        end
        149: begin
            cosine_reg0 <= 36'sb11111001010101111001101001001110111;
            sine_reg0   <= 36'sb111010000000010000100001111001001;
        end
        150: begin
            cosine_reg0 <= 36'sb11111001010000001011111111100010001;
            sine_reg0   <= 36'sb111010011000101110111010011010011;
        end
        151: begin
            cosine_reg0 <= 36'sb11111001001010011011111100000101001;
            sine_reg0   <= 36'sb111010110001001100101110111010100;
        end
        152: begin
            cosine_reg0 <= 36'sb11111001000100101001011110111011101;
            sine_reg0   <= 36'sb111011001001101001111111001010100;
        end
        153: begin
            cosine_reg0 <= 36'sb11111000111110110100101000001001000;
            sine_reg0   <= 36'sb111011100010000110101010111011011;
        end
        154: begin
            cosine_reg0 <= 36'sb11111000111000111101010111110001001;
            sine_reg0   <= 36'sb111011111010100010110001111110000;
        end
        155: begin
            cosine_reg0 <= 36'sb11111000110011000011101101110111100;
            sine_reg0   <= 36'sb111100010010111110010100000011010;
        end
        156: begin
            cosine_reg0 <= 36'sb11111000101101000111101010011111101;
            sine_reg0   <= 36'sb111100101011011001010000111100001;
        end
        157: begin
            cosine_reg0 <= 36'sb11111000100111001001001101101101010;
            sine_reg0   <= 36'sb111101000011110011101000011001100;
        end
        158: begin
            cosine_reg0 <= 36'sb11111000100001001000010111100100001;
            sine_reg0   <= 36'sb111101011100001101011010001100011;
        end
        159: begin
            cosine_reg0 <= 36'sb11111000011011000101001000001000000;
            sine_reg0   <= 36'sb111101110100100110100110000101101;
        end
        160: begin
            cosine_reg0 <= 36'sb11111000010100111111011111011100100;
            sine_reg0   <= 36'sb111110001100111111001011110110010;
        end
        161: begin
            cosine_reg0 <= 36'sb11111000001110110111011101100101011;
            sine_reg0   <= 36'sb111110100101010111001011001111010;
        end
        162: begin
            cosine_reg0 <= 36'sb11111000001000101101000010100110011;
            sine_reg0   <= 36'sb111110111101101110100100000001100;
        end
        163: begin
            cosine_reg0 <= 36'sb11111000000010100000001110100011011;
            sine_reg0   <= 36'sb111111010110000101010101111110000;
        end
        164: begin
            cosine_reg0 <= 36'sb11110111111100010001000001100000010;
            sine_reg0   <= 36'sb111111101110011011100000110101110;
        end
        165: begin
            cosine_reg0 <= 36'sb11110111110101111111011011100000110;
            sine_reg0   <= 36'sb1000000000110110001000100011001110;
        end
        166: begin
            cosine_reg0 <= 36'sb11110111101111101011011100101000110;
            sine_reg0   <= 36'sb1000000011111000110000000011010111;
        end
        167: begin
            cosine_reg0 <= 36'sb11110111101001010101000100111100010;
            sine_reg0   <= 36'sb1000000110111011010010100101010010;
        end
        168: begin
            cosine_reg0 <= 36'sb11110111100010111100010100011111000;
            sine_reg0   <= 36'sb1000001001111101110000000111000111;
        end
        169: begin
            cosine_reg0 <= 36'sb11110111011100100001001011010101001;
            sine_reg0   <= 36'sb1000001101000000001000100110111101;
        end
        170: begin
            cosine_reg0 <= 36'sb11110111010110000011101001100010011;
            sine_reg0   <= 36'sb1000010000000010011100000010111101;
        end
        171: begin
            cosine_reg0 <= 36'sb11110111001111100011101111001010111;
            sine_reg0   <= 36'sb1000010011000100101010011001001111;
        end
        172: begin
            cosine_reg0 <= 36'sb11110111001001000001011100010010110;
            sine_reg0   <= 36'sb1000010110000110110011100111111011;
        end
        173: begin
            cosine_reg0 <= 36'sb11110111000010011100110000111101110;
            sine_reg0   <= 36'sb1000011001001000110111101101001010;
        end
        174: begin
            cosine_reg0 <= 36'sb11110110111011110101101101010000001;
            sine_reg0   <= 36'sb1000011100001010110110100111000011;
        end
        175: begin
            cosine_reg0 <= 36'sb11110110110101001100010001001101111;
            sine_reg0   <= 36'sb1000011111001100110000010011101111;
        end
        176: begin
            cosine_reg0 <= 36'sb11110110101110100000011100111011001;
            sine_reg0   <= 36'sb1000100010001110100100110001010110;
        end
        177: begin
            cosine_reg0 <= 36'sb11110110100111110010010000011100000;
            sine_reg0   <= 36'sb1000100101010000010011111110000001;
        end
        178: begin
            cosine_reg0 <= 36'sb11110110100001000001101011110100101;
            sine_reg0   <= 36'sb1000101000010001111101110111111001;
        end
        179: begin
            cosine_reg0 <= 36'sb11110110011010001110101111001001010;
            sine_reg0   <= 36'sb1000101011010011100010011101000101;
        end
        180: begin
            cosine_reg0 <= 36'sb11110110010011011001011010011110000;
            sine_reg0   <= 36'sb1000101110010101000001101011101111;
        end
        181: begin
            cosine_reg0 <= 36'sb11110110001100100001101101110111001;
            sine_reg0   <= 36'sb1000110001010110011011100001111110;
        end
        182: begin
            cosine_reg0 <= 36'sb11110110000101100111101001011000110;
            sine_reg0   <= 36'sb1000110100010111101111111101111101;
        end
        183: begin
            cosine_reg0 <= 36'sb11110101111110101011001101000111010;
            sine_reg0   <= 36'sb1000110111011000111110111101110011;
        end
        184: begin
            cosine_reg0 <= 36'sb11110101110111101100011001000110111;
            sine_reg0   <= 36'sb1000111010011010001000011111101001;
        end
        185: begin
            cosine_reg0 <= 36'sb11110101110000101011001101011011111;
            sine_reg0   <= 36'sb1000111101011011001100100001101001;
        end
        186: begin
            cosine_reg0 <= 36'sb11110101101001100111101010001010110;
            sine_reg0   <= 36'sb1001000000011100001011000001111011;
        end
        187: begin
            cosine_reg0 <= 36'sb11110101100010100001101111010111101;
            sine_reg0   <= 36'sb1001000011011101000011111110100111;
        end
        188: begin
            cosine_reg0 <= 36'sb11110101011011011001011101000111001;
            sine_reg0   <= 36'sb1001000110011101110111010101111000;
        end
        189: begin
            cosine_reg0 <= 36'sb11110101010100001110110011011101100;
            sine_reg0   <= 36'sb1001001001011110100101000101110110;
        end
        190: begin
            cosine_reg0 <= 36'sb11110101001101000001110010011111001;
            sine_reg0   <= 36'sb1001001100011111001101001100101010;
        end
        191: begin
            cosine_reg0 <= 36'sb11110101000101110010011010010000100;
            sine_reg0   <= 36'sb1001001111011111101111101000011110;
        end
        192: begin
            cosine_reg0 <= 36'sb11110100111110100000101010110110001;
            sine_reg0   <= 36'sb1001010010100000001100010111011010;
        end
        193: begin
            cosine_reg0 <= 36'sb11110100110111001100100100010100011;
            sine_reg0   <= 36'sb1001010101100000100011010111101001;
        end
        194: begin
            cosine_reg0 <= 36'sb11110100101111110110000110101111111;
            sine_reg0   <= 36'sb1001011000100000110100100111010010;
        end
        195: begin
            cosine_reg0 <= 36'sb11110100101000011101010010001101010;
            sine_reg0   <= 36'sb1001011011100001000000000100100001;
        end
        196: begin
            cosine_reg0 <= 36'sb11110100100001000010000110110000111;
            sine_reg0   <= 36'sb1001011110100001000101101101011101;
        end
        197: begin
            cosine_reg0 <= 36'sb11110100011001100100100100011111010;
            sine_reg0   <= 36'sb1001100001100001000101100000010001;
        end
        198: begin
            cosine_reg0 <= 36'sb11110100010010000100101011011101010;
            sine_reg0   <= 36'sb1001100100100000111111011011000111;
        end
        199: begin
            cosine_reg0 <= 36'sb11110100001010100010011011101111011;
            sine_reg0   <= 36'sb1001100111100000110011011100000111;
        end
        200: begin
            cosine_reg0 <= 36'sb11110100000010111101110101011010010;
            sine_reg0   <= 36'sb1001101010100000100001100001011100;
        end
        201: begin
            cosine_reg0 <= 36'sb11110011111011010110111000100010101;
            sine_reg0   <= 36'sb1001101101100000001001101001001111;
        end
        202: begin
            cosine_reg0 <= 36'sb11110011110011101101100101001101000;
            sine_reg0   <= 36'sb1001110000011111101011110001101010;
        end
        203: begin
            cosine_reg0 <= 36'sb11110011101100000001111011011110011;
            sine_reg0   <= 36'sb1001110011011111000111111000110111;
        end
        204: begin
            cosine_reg0 <= 36'sb11110011100100010011111011011011010;
            sine_reg0   <= 36'sb1001110110011110011101111101000000;
        end
        205: begin
            cosine_reg0 <= 36'sb11110011011100100011100101001000100;
            sine_reg0   <= 36'sb1001111001011101101101111100001111;
        end
        206: begin
            cosine_reg0 <= 36'sb11110011010100110000111000101010110;
            sine_reg0   <= 36'sb1001111100011100110111110100101110;
        end
        207: begin
            cosine_reg0 <= 36'sb11110011001100111011110110000111001;
            sine_reg0   <= 36'sb1001111111011011111011100100100110;
        end
        208: begin
            cosine_reg0 <= 36'sb11110011000101000100011101100010001;
            sine_reg0   <= 36'sb1010000010011010111001001010000011;
        end
        209: begin
            cosine_reg0 <= 36'sb11110010111101001010101111000000111;
            sine_reg0   <= 36'sb1010000101011001110000100011001101;
        end
        210: begin
            cosine_reg0 <= 36'sb11110010110101001110101010101000000;
            sine_reg0   <= 36'sb1010001000011000100001101110010001;
        end
        211: begin
            cosine_reg0 <= 36'sb11110010101101010000010000011100101;
            sine_reg0   <= 36'sb1010001011010111001100101001010111;
        end
        212: begin
            cosine_reg0 <= 36'sb11110010100101001111100000100011100;
            sine_reg0   <= 36'sb1010001110010101110001010010101011;
        end
        213: begin
            cosine_reg0 <= 36'sb11110010011101001100011011000001101;
            sine_reg0   <= 36'sb1010010001010100001111101000010110;
        end
        214: begin
            cosine_reg0 <= 36'sb11110010010101000110111111111100000;
            sine_reg0   <= 36'sb1010010100010010100111101000100011;
        end
        215: begin
            cosine_reg0 <= 36'sb11110010001100111111001111010111100;
            sine_reg0   <= 36'sb1010010111010000111001010001011101;
        end
        216: begin
            cosine_reg0 <= 36'sb11110010000100110101001001011001010;
            sine_reg0   <= 36'sb1010011010001111000100100001001111;
        end
        217: begin
            cosine_reg0 <= 36'sb11110001111100101000101110000110010;
            sine_reg0   <= 36'sb1010011101001101001001010110000010;
        end
        218: begin
            cosine_reg0 <= 36'sb11110001110100011001111101100011101;
            sine_reg0   <= 36'sb1010100000001011000111101110000011;
        end
        219: begin
            cosine_reg0 <= 36'sb11110001101100001000110111110110010;
            sine_reg0   <= 36'sb1010100011001000111111100111011011;
        end
        220: begin
            cosine_reg0 <= 36'sb11110001100011110101011101000011011;
            sine_reg0   <= 36'sb1010100110000110110001000000010110;
        end
        221: begin
            cosine_reg0 <= 36'sb11110001011011011111101101010000001;
            sine_reg0   <= 36'sb1010101001000100011011110110111110;
        end
        222: begin
            cosine_reg0 <= 36'sb11110001010011000111101000100001101;
            sine_reg0   <= 36'sb1010101100000010000000001001011110;
        end
        223: begin
            cosine_reg0 <= 36'sb11110001001010101101001110111101001;
            sine_reg0   <= 36'sb1010101110111111011101110110000010;
        end
        224: begin
            cosine_reg0 <= 36'sb11110001000010010000100000100111101;
            sine_reg0   <= 36'sb1010110001111100110100111010110101;
        end
        225: begin
            cosine_reg0 <= 36'sb11110000111001110001011101100110011;
            sine_reg0   <= 36'sb1010110100111010000101010110000010;
        end
        226: begin
            cosine_reg0 <= 36'sb11110000110001010000000101111110110;
            sine_reg0   <= 36'sb1010110111110111001111000101110011;
        end
        227: begin
            cosine_reg0 <= 36'sb11110000101000101100011001110101111;
            sine_reg0   <= 36'sb1010111010110100010010001000010110;
        end
        228: begin
            cosine_reg0 <= 36'sb11110000100000000110011001010001001;
            sine_reg0   <= 36'sb1010111101110001001110011011110011;
        end
        229: begin
            cosine_reg0 <= 36'sb11110000010111011110000100010101110;
            sine_reg0   <= 36'sb1011000000101110000011111110011001;
        end
        230: begin
            cosine_reg0 <= 36'sb11110000001110110011011011001001001;
            sine_reg0   <= 36'sb1011000011101010110010101110010001;
        end
        231: begin
            cosine_reg0 <= 36'sb11110000000110000110011101110000100;
            sine_reg0   <= 36'sb1011000110100111011010101001100111;
        end
        232: begin
            cosine_reg0 <= 36'sb11101111111101010111001100010001010;
            sine_reg0   <= 36'sb1011001001100011111011101110101000;
        end
        233: begin
            cosine_reg0 <= 36'sb11101111110100100101100110110000111;
            sine_reg0   <= 36'sb1011001100100000010101111011011110;
        end
        234: begin
            cosine_reg0 <= 36'sb11101111101011110001101101010100110;
            sine_reg0   <= 36'sb1011001111011100101001001110010101;
        end
        235: begin
            cosine_reg0 <= 36'sb11101111100010111011100000000010010;
            sine_reg0   <= 36'sb1011010010011000110101100101011010;
        end
        236: begin
            cosine_reg0 <= 36'sb11101111011010000010111110111110111;
            sine_reg0   <= 36'sb1011010101010100111010111110111001;
        end
        237: begin
            cosine_reg0 <= 36'sb11101111010001001000001010010000000;
            sine_reg0   <= 36'sb1011011000010000111001011000111100;
        end
        238: begin
            cosine_reg0 <= 36'sb11101111001000001011000001111011010;
            sine_reg0   <= 36'sb1011011011001100110000110001110001;
        end
        239: begin
            cosine_reg0 <= 36'sb11101110111111001011100110000110010;
            sine_reg0   <= 36'sb1011011110001000100001000111100011;
        end
        240: begin
            cosine_reg0 <= 36'sb11101110110110001001110110110110010;
            sine_reg0   <= 36'sb1011100001000100001010011000011111;
        end
        241: begin
            cosine_reg0 <= 36'sb11101110101101000101110100010001001;
            sine_reg0   <= 36'sb1011100011111111101100100010110001;
        end
        242: begin
            cosine_reg0 <= 36'sb11101110100011111111011110011100010;
            sine_reg0   <= 36'sb1011100110111011000111100100100100;
        end
        243: begin
            cosine_reg0 <= 36'sb11101110011010110110110101011101010;
            sine_reg0   <= 36'sb1011101001110110011011011100000111;
        end
        244: begin
            cosine_reg0 <= 36'sb11101110010001101011111001011001111;
            sine_reg0   <= 36'sb1011101100110001101000000111100100;
        end
        245: begin
            cosine_reg0 <= 36'sb11101110001000011110101010010111110;
            sine_reg0   <= 36'sb1011101111101100101101100101001001;
        end
        246: begin
            cosine_reg0 <= 36'sb11101101111111001111001000011100100;
            sine_reg0   <= 36'sb1011110010100111101011110011000010;
        end
        247: begin
            cosine_reg0 <= 36'sb11101101110101111101010011101110000;
            sine_reg0   <= 36'sb1011110101100010100010101111011100;
        end
        248: begin
            cosine_reg0 <= 36'sb11101101101100101001001100010001101;
            sine_reg0   <= 36'sb1011111000011101010010011000100011;
        end
        249: begin
            cosine_reg0 <= 36'sb11101101100011010010110010001101100;
            sine_reg0   <= 36'sb1011111011010111111010101100100101;
        end
        250: begin
            cosine_reg0 <= 36'sb11101101011001111010000101100111001;
            sine_reg0   <= 36'sb1011111110010010011011101001101110;
        end
        251: begin
            cosine_reg0 <= 36'sb11101101010000011111000110100100011;
            sine_reg0   <= 36'sb1100000001001100110101001110001011;
        end
        252: begin
            cosine_reg0 <= 36'sb11101101000111000001110101001011001;
            sine_reg0   <= 36'sb1100000100000111000111011000001001;
        end
        253: begin
            cosine_reg0 <= 36'sb11101100111101100010010001100001001;
            sine_reg0   <= 36'sb1100000111000001010010000101110110;
        end
        254: begin
            cosine_reg0 <= 36'sb11101100110100000000011011101100010;
            sine_reg0   <= 36'sb1100001001111011010101010101011110;
        end
        255: begin
            cosine_reg0 <= 36'sb11101100101010011100010011110010011;
            sine_reg0   <= 36'sb1100001100110101010001000101001111;
        end
        256: begin
            cosine_reg0 <= 36'sb11101100100000110101111001111001100;
            sine_reg0   <= 36'sb1100001111101111000101010011010101;
        end
        257: begin
            cosine_reg0 <= 36'sb11101100010111001101001110000111011;
            sine_reg0   <= 36'sb1100010010101000110001111101111111;
        end
        258: begin
            cosine_reg0 <= 36'sb11101100001101100010010000100010000;
            sine_reg0   <= 36'sb1100010101100010010111000011011010;
        end
        259: begin
            cosine_reg0 <= 36'sb11101100000011110101000001001111100;
            sine_reg0   <= 36'sb1100011000011011110100100001110100;
        end
        260: begin
            cosine_reg0 <= 36'sb11101011111010000101100000010101101;
            sine_reg0   <= 36'sb1100011011010101001010010111011001;
        end
        261: begin
            cosine_reg0 <= 36'sb11101011110000010011101101111010101;
            sine_reg0   <= 36'sb1100011110001110011000100010010111;
        end
        262: begin
            cosine_reg0 <= 36'sb11101011100110011111101010000100010;
            sine_reg0   <= 36'sb1100100001000111011111000000111110;
        end
        263: begin
            cosine_reg0 <= 36'sb11101011011100101001010100111000110;
            sine_reg0   <= 36'sb1100100100000000011101110001011001;
        end
        264: begin
            cosine_reg0 <= 36'sb11101011010010110000101110011110010;
            sine_reg0   <= 36'sb1100100110111001010100110001110111;
        end
        265: begin
            cosine_reg0 <= 36'sb11101011001000110101110110111010101;
            sine_reg0   <= 36'sb1100101001110010000100000000100111;
        end
        266: begin
            cosine_reg0 <= 36'sb11101010111110111000101110010100001;
            sine_reg0   <= 36'sb1100101100101010101011011011110101;
        end
        267: begin
            cosine_reg0 <= 36'sb11101010110100111001010100110001000;
            sine_reg0   <= 36'sb1100101111100011001011000001110001;
        end
        268: begin
            cosine_reg0 <= 36'sb11101010101010110111101010010111001;
            sine_reg0   <= 36'sb1100110010011011100010110000101000;
        end
        269: begin
            cosine_reg0 <= 36'sb11101010100000110011101111001101000;
            sine_reg0   <= 36'sb1100110101010011110010100110101001;
        end
        270: begin
            cosine_reg0 <= 36'sb11101010010110101101100011011000101;
            sine_reg0   <= 36'sb1100111000001011111010100010000001;
        end
        271: begin
            cosine_reg0 <= 36'sb11101010001100100101000111000000011;
            sine_reg0   <= 36'sb1100111011000011111010100001000001;
        end
        272: begin
            cosine_reg0 <= 36'sb11101010000010011010011010001010011;
            sine_reg0   <= 36'sb1100111101111011110010100001110101;
        end
        273: begin
            cosine_reg0 <= 36'sb11101001111000001101011100111100111;
            sine_reg0   <= 36'sb1101000000110011100010100010101100;
        end
        274: begin
            cosine_reg0 <= 36'sb11101001101101111110001111011110010;
            sine_reg0   <= 36'sb1101000011101011001010100001110110;
        end
        275: begin
            cosine_reg0 <= 36'sb11101001100011101100110001110100111;
            sine_reg0   <= 36'sb1101000110100010101010011101100001;
        end
        276: begin
            cosine_reg0 <= 36'sb11101001011001011001000100000110111;
            sine_reg0   <= 36'sb1101001001011010000010010011111011;
        end
        277: begin
            cosine_reg0 <= 36'sb11101001001111000011000110011010111;
            sine_reg0   <= 36'sb1101001100010001010010000011010100;
        end
        278: begin
            cosine_reg0 <= 36'sb11101001000100101010111000110111001;
            sine_reg0   <= 36'sb1101001111001000011001101001111011;
        end
        279: begin
            cosine_reg0 <= 36'sb11101000111010010000011011100001111;
            sine_reg0   <= 36'sb1101010001111111011001000101111110;
        end
        280: begin
            cosine_reg0 <= 36'sb11101000101111110011101110100001111;
            sine_reg0   <= 36'sb1101010100110110010000010101101101;
        end
        281: begin
            cosine_reg0 <= 36'sb11101000100101010100110001111101010;
            sine_reg0   <= 36'sb1101010111101100111111010111010111;
        end
        282: begin
            cosine_reg0 <= 36'sb11101000011010110011100101111010110;
            sine_reg0   <= 36'sb1101011010100011100110001001001011;
        end
        283: begin
            cosine_reg0 <= 36'sb11101000010000010000001010100000101;
            sine_reg0   <= 36'sb1101011101011010000100101001011001;
        end
        284: begin
            cosine_reg0 <= 36'sb11101000000101101010011111110101100;
            sine_reg0   <= 36'sb1101100000010000011010110110001111;
        end
        285: begin
            cosine_reg0 <= 36'sb11100111111011000010100101111111111;
            sine_reg0   <= 36'sb1101100011000110101000101101111111;
        end
        286: begin
            cosine_reg0 <= 36'sb11100111110000011000011101000110011;
            sine_reg0   <= 36'sb1101100101111100101110001110110110;
        end
        287: begin
            cosine_reg0 <= 36'sb11100111100101101100000101001111100;
            sine_reg0   <= 36'sb1101101000110010101011010111000101;
        end
        288: begin
            cosine_reg0 <= 36'sb11100111011010111101011110100001110;
            sine_reg0   <= 36'sb1101101011101000100000000100111100;
        end
        289: begin
            cosine_reg0 <= 36'sb11100111010000001100101001000100000;
            sine_reg0   <= 36'sb1101101110011110001100010110101010;
        end
        290: begin
            cosine_reg0 <= 36'sb11100111000101011001100100111100110;
            sine_reg0   <= 36'sb1101110001010011110000001010011111;
        end
        291: begin
            cosine_reg0 <= 36'sb11100110111010100100010010010010100;
            sine_reg0   <= 36'sb1101110100001001001011011110101100;
        end
        292: begin
            cosine_reg0 <= 36'sb11100110101111101100110001001100010;
            sine_reg0   <= 36'sb1101110110111110011110010001100000;
        end
        293: begin
            cosine_reg0 <= 36'sb11100110100100110011000001110000100;
            sine_reg0   <= 36'sb1101111001110011101000100001001100;
        end
        294: begin
            cosine_reg0 <= 36'sb11100110011001110111000100000110000;
            sine_reg0   <= 36'sb1101111100101000101010001100000000;
        end
        295: begin
            cosine_reg0 <= 36'sb11100110001110111000111000010011100;
            sine_reg0   <= 36'sb1101111111011101100011010000001011;
        end
        296: begin
            cosine_reg0 <= 36'sb11100110000011111000011110011111110;
            sine_reg0   <= 36'sb1110000010010010010011101100000000;
        end
        297: begin
            cosine_reg0 <= 36'sb11100101111000110101110110110001101;
            sine_reg0   <= 36'sb1110000101000110111011011101101101;
        end
        298: begin
            cosine_reg0 <= 36'sb11100101101101110001000001001111111;
            sine_reg0   <= 36'sb1110000111111011011010100011100100;
        end
        299: begin
            cosine_reg0 <= 36'sb11100101100010101001111110000001011;
            sine_reg0   <= 36'sb1110001010101111110000111011110110;
        end
        300: begin
            cosine_reg0 <= 36'sb11100101010111100000101101001100111;
            sine_reg0   <= 36'sb1110001101100011111110100100110010;
        end
        301: begin
            cosine_reg0 <= 36'sb11100101001100010101001110111001011;
            sine_reg0   <= 36'sb1110010000011000000011011100101011;
        end
        302: begin
            cosine_reg0 <= 36'sb11100101000001000111100011001101110;
            sine_reg0   <= 36'sb1110010011001011111111100001110000;
        end
        303: begin
            cosine_reg0 <= 36'sb11100100110101110111101010010000110;
            sine_reg0   <= 36'sb1110010101111111110010110010010100;
        end
        304: begin
            cosine_reg0 <= 36'sb11100100101010100101100100001001100;
            sine_reg0   <= 36'sb1110011000110011011101001100100110;
        end
        305: begin
            cosine_reg0 <= 36'sb11100100011111010001010000111110111;
            sine_reg0   <= 36'sb1110011011100110111110101110111000;
        end
        306: begin
            cosine_reg0 <= 36'sb11100100010011111010110000111000000;
            sine_reg0   <= 36'sb1110011110011010010111010111011100;
        end
        307: begin
            cosine_reg0 <= 36'sb11100100001000100010000011111011101;
            sine_reg0   <= 36'sb1110100001001101100111000100100010;
        end
        308: begin
            cosine_reg0 <= 36'sb11100011111101000111001010010001000;
            sine_reg0   <= 36'sb1110100100000000101101110100011101;
        end
        309: begin
            cosine_reg0 <= 36'sb11100011110001101010000011111111000;
            sine_reg0   <= 36'sb1110100110110011101011100101011101;
        end
        310: begin
            cosine_reg0 <= 36'sb11100011100110001010110001001100111;
            sine_reg0   <= 36'sb1110101001100110100000010101110101;
        end
        311: begin
            cosine_reg0 <= 36'sb11100011011010101001010010000001100;
            sine_reg0   <= 36'sb1110101100011001001100000011110101;
        end
        312: begin
            cosine_reg0 <= 36'sb11100011001111000101100110100100001;
            sine_reg0   <= 36'sb1110101111001011101110101101110000;
        end
        313: begin
            cosine_reg0 <= 36'sb11100011000011011111101110111011111;
            sine_reg0   <= 36'sb1110110001111110001000010001111000;
        end
        314: begin
            cosine_reg0 <= 36'sb11100010110111110111101011001111111;
            sine_reg0   <= 36'sb1110110100110000011000101110011111;
        end
        315: begin
            cosine_reg0 <= 36'sb11100010101100001101011011100111010;
            sine_reg0   <= 36'sb1110110111100010100000000001110110;
        end
        316: begin
            cosine_reg0 <= 36'sb11100010100000100001000000001001010;
            sine_reg0   <= 36'sb1110111010010100011110001010010000;
        end
        317: begin
            cosine_reg0 <= 36'sb11100010010100110010011000111101001;
            sine_reg0   <= 36'sb1110111101000110010011000101111111;
        end
        318: begin
            cosine_reg0 <= 36'sb11100010001001000001100110001010000;
            sine_reg0   <= 36'sb1110111111110111111110110011010101;
        end
        319: begin
            cosine_reg0 <= 36'sb11100001111101001110100111110111001;
            sine_reg0   <= 36'sb1111000010101001100001010000100100;
        end
        320: begin
            cosine_reg0 <= 36'sb11100001110001011001011110001011111;
            sine_reg0   <= 36'sb1111000101011010111010011100000000;
        end
        321: begin
            cosine_reg0 <= 36'sb11100001100101100010001001001111101;
            sine_reg0   <= 36'sb1111001000001100001010010011111011;
        end
        322: begin
            cosine_reg0 <= 36'sb11100001011001101000101001001001100;
            sine_reg0   <= 36'sb1111001010111101010000110110100111;
        end
        323: begin
            cosine_reg0 <= 36'sb11100001001101101100111110000000111;
            sine_reg0   <= 36'sb1111001101101110001110000010010111;
        end
        324: begin
            cosine_reg0 <= 36'sb11100001000001101111000111111101001;
            sine_reg0   <= 36'sb1111010000011111000001110101011111;
        end
        325: begin
            cosine_reg0 <= 36'sb11100000110101101111000111000101110;
            sine_reg0   <= 36'sb1111010011001111101100001110010000;
        end
        326: begin
            cosine_reg0 <= 36'sb11100000101001101100111011100010001;
            sine_reg0   <= 36'sb1111010110000000001101001010111110;
        end
        327: begin
            cosine_reg0 <= 36'sb11100000011101101000100101011001100;
            sine_reg0   <= 36'sb1111011000110000100100101001111100;
        end
        328: begin
            cosine_reg0 <= 36'sb11100000010001100010000100110011100;
            sine_reg0   <= 36'sb1111011011100000110010101001011101;
        end
        329: begin
            cosine_reg0 <= 36'sb11100000000101011001011001110111100;
            sine_reg0   <= 36'sb1111011110010000110111000111110101;
        end
        330: begin
            cosine_reg0 <= 36'sb11011111111001001110100100101101000;
            sine_reg0   <= 36'sb1111100001000000110010000011011000;
        end
        331: begin
            cosine_reg0 <= 36'sb11011111101101000001100101011011100;
            sine_reg0   <= 36'sb1111100011110000100011011010010111;
        end
        332: begin
            cosine_reg0 <= 36'sb11011111100000110010011100001010100;
            sine_reg0   <= 36'sb1111100110100000001011001011000111;
        end
        333: begin
            cosine_reg0 <= 36'sb11011111010100100001001001000001101;
            sine_reg0   <= 36'sb1111101001001111101001010011111101;
        end
        334: begin
            cosine_reg0 <= 36'sb11011111001000001101101100001000011;
            sine_reg0   <= 36'sb1111101011111110111101110011001010;
        end
        335: begin
            cosine_reg0 <= 36'sb11011110111011111000000101100110100;
            sine_reg0   <= 36'sb1111101110101110001000100111000100;
        end
        336: begin
            cosine_reg0 <= 36'sb11011110101111100000010101100011011;
            sine_reg0   <= 36'sb1111110001011101001001101101111111;
        end
        337: begin
            cosine_reg0 <= 36'sb11011110100011000110011100000110110;
            sine_reg0   <= 36'sb1111110100001100000001000110001101;
        end
        338: begin
            cosine_reg0 <= 36'sb11011110010110101010011001011000010;
            sine_reg0   <= 36'sb1111110110111010101110101110000100;
        end
        339: begin
            cosine_reg0 <= 36'sb11011110001010001100001101011111101;
            sine_reg0   <= 36'sb1111111001101001010010100011111000;
        end
        340: begin
            cosine_reg0 <= 36'sb11011101111101101011111000100100100;
            sine_reg0   <= 36'sb1111111100010111101100100101111100;
        end
        341: begin
            cosine_reg0 <= 36'sb11011101110001001001011010101110101;
            sine_reg0   <= 36'sb1111111111000101111100110010100110;
        end
        342: begin
            cosine_reg0 <= 36'sb11011101100100100100110100000101101;
            sine_reg0   <= 36'sb10000000001110100000011001000001010;
        end
        343: begin
            cosine_reg0 <= 36'sb11011101010111111110000100110001011;
            sine_reg0   <= 36'sb10000000100100001111111100100111101;
        end
        344: begin
            cosine_reg0 <= 36'sb11011101001011010101001100111001101;
            sine_reg0   <= 36'sb10000000111001111110010000111010011;
        end
        345: begin
            cosine_reg0 <= 36'sb11011100111110101010001100100110001;
            sine_reg0   <= 36'sb10000001001111101011010101101100000;
        end
        346: begin
            cosine_reg0 <= 36'sb11011100110001111101000011111110101;
            sine_reg0   <= 36'sb10000001100101010111001010101111011;
        end
        347: begin
            cosine_reg0 <= 36'sb11011100100101001101110011001011010;
            sine_reg0   <= 36'sb10000001111011000001101111110110111;
        end
        348: begin
            cosine_reg0 <= 36'sb11011100011000011100011010010011100;
            sine_reg0   <= 36'sb10000010010000101011000100110101011;
        end
        349: begin
            cosine_reg0 <= 36'sb11011100001011101000111001011111100;
            sine_reg0   <= 36'sb10000010100110010011001001011101011;
        end
        350: begin
            cosine_reg0 <= 36'sb11011011111110110011010000110111001;
            sine_reg0   <= 36'sb10000010111011111001111101100001100;
        end
        351: begin
            cosine_reg0 <= 36'sb11011011110001111011100000100010010;
            sine_reg0   <= 36'sb10000011010001011111100000110100100;
        end
        352: begin
            cosine_reg0 <= 36'sb11011011100101000001101000101000101;
            sine_reg0   <= 36'sb10000011100111000011110011001001000;
        end
        353: begin
            cosine_reg0 <= 36'sb11011011011000000101101001010010101;
            sine_reg0   <= 36'sb10000011111100100110110100010001110;
        end
        354: begin
            cosine_reg0 <= 36'sb11011011001011000111100010100111111;
            sine_reg0   <= 36'sb10000100010010001000100100000001100;
        end
        355: begin
            cosine_reg0 <= 36'sb11011010111110000111010100110000100;
            sine_reg0   <= 36'sb10000100100111101001000010001010111;
        end
        356: begin
            cosine_reg0 <= 36'sb11011010110001000100111111110100100;
            sine_reg0   <= 36'sb10000100111101001000001110100000101;
        end
        357: begin
            cosine_reg0 <= 36'sb11011010100100000000100011111011111;
            sine_reg0   <= 36'sb10000101010010100110001000110101101;
        end
        358: begin
            cosine_reg0 <= 36'sb11011010010110111010000001001110111;
            sine_reg0   <= 36'sb10000101101000000010110000111100011;
        end
        359: begin
            cosine_reg0 <= 36'sb11011010001001110001010111110101011;
            sine_reg0   <= 36'sb10000101111101011110000110100111111;
        end
        360: begin
            cosine_reg0 <= 36'sb11011001111100100110100111110111100;
            sine_reg0   <= 36'sb10000110010010111000001001101010111;
        end
        361: begin
            cosine_reg0 <= 36'sb11011001101111011001110001011101100;
            sine_reg0   <= 36'sb10000110101000010000111001111000000;
        end
        362: begin
            cosine_reg0 <= 36'sb11011001100010001010110100101111100;
            sine_reg0   <= 36'sb10000110111101101000010111000010010;
        end
        363: begin
            cosine_reg0 <= 36'sb11011001010100111001110001110101100;
            sine_reg0   <= 36'sb10000111010010111110100000111100011;
        end
        364: begin
            cosine_reg0 <= 36'sb11011001000111100110101000110111111;
            sine_reg0   <= 36'sb10000111101000010011010111011001010;
        end
        365: begin
            cosine_reg0 <= 36'sb11011000111010010001011001111110110;
            sine_reg0   <= 36'sb10000111111101100110111010001011101;
        end
        366: begin
            cosine_reg0 <= 36'sb11011000101100111010000101010010010;
            sine_reg0   <= 36'sb10001000010010111001001001000110100;
        end
        367: begin
            cosine_reg0 <= 36'sb11011000011111100000101010111010110;
            sine_reg0   <= 36'sb10001000101000001010000011111100100;
        end
        368: begin
            cosine_reg0 <= 36'sb11011000010010000101001011000000100;
            sine_reg0   <= 36'sb10001000111101011001101010100000110;
        end
        369: begin
            cosine_reg0 <= 36'sb11011000000100100111100101101011110;
            sine_reg0   <= 36'sb10001001010010100111111100100110001;
        end
        370: begin
            cosine_reg0 <= 36'sb11010111110111000111111011000100111;
            sine_reg0   <= 36'sb10001001100111110100111001111111011;
        end
        371: begin
            cosine_reg0 <= 36'sb11010111101001100110001011010100001;
            sine_reg0   <= 36'sb10001001111101000000100010011111100;
        end
        372: begin
            cosine_reg0 <= 36'sb11010111011100000010010110100001110;
            sine_reg0   <= 36'sb10001010010010001010110101111001100;
        end
        373: begin
            cosine_reg0 <= 36'sb11010111001110011100011100110110010;
            sine_reg0   <= 36'sb10001010100111010011110100000000010;
        end
        374: begin
            cosine_reg0 <= 36'sb11010111000000110100011110011010001;
            sine_reg0   <= 36'sb10001010111100011011011100100110110;
        end
        375: begin
            cosine_reg0 <= 36'sb11010110110011001010011011010101100;
            sine_reg0   <= 36'sb10001011010001100001101111100000000;
        end
        376: begin
            cosine_reg0 <= 36'sb11010110100101011110010011110001000;
            sine_reg0   <= 36'sb10001011100110100110101100011110111;
        end
        377: begin
            cosine_reg0 <= 36'sb11010110010111110000000111110100111;
            sine_reg0   <= 36'sb10001011111011101010010011010110100;
        end
        378: begin
            cosine_reg0 <= 36'sb11010110001001111111110111101001111;
            sine_reg0   <= 36'sb10001100010000101100100011111001110;
        end
        379: begin
            cosine_reg0 <= 36'sb11010101111100001101100011011000010;
            sine_reg0   <= 36'sb10001100100101101101011101111011110;
        end
        380: begin
            cosine_reg0 <= 36'sb11010101101110011001001011001000101;
            sine_reg0   <= 36'sb10001100111010101101000001001111100;
        end
        381: begin
            cosine_reg0 <= 36'sb11010101100000100010101111000011100;
            sine_reg0   <= 36'sb10001101001111101011001101101000001;
        end
        382: begin
            cosine_reg0 <= 36'sb11010101010010101010001111010001010;
            sine_reg0   <= 36'sb10001101100100101000000010111000100;
        end
        383: begin
            cosine_reg0 <= 36'sb11010101000100101111101011111010110;
            sine_reg0   <= 36'sb10001101111001100011100000110100000;
        end
        384: begin
            cosine_reg0 <= 36'sb11010100110110110011000101001000011;
            sine_reg0   <= 36'sb10001110001110011101100111001101011;
        end
        385: begin
            cosine_reg0 <= 36'sb11010100101000110100011011000010110;
            sine_reg0   <= 36'sb10001110100011010110010101111000000;
        end
        386: begin
            cosine_reg0 <= 36'sb11010100011010110011101101110010100;
            sine_reg0   <= 36'sb10001110111000001101101100100110111;
        end
        387: begin
            cosine_reg0 <= 36'sb11010100001100110000111101100000011;
            sine_reg0   <= 36'sb10001111001101000011101011001101000;
        end
        388: begin
            cosine_reg0 <= 36'sb11010011111110101100001010010100111;
            sine_reg0   <= 36'sb10001111100001111000010001011101111;
        end
        389: begin
            cosine_reg0 <= 36'sb11010011110000100101010100011000110;
            sine_reg0   <= 36'sb10001111110110101011011111001100010;
        end
        390: begin
            cosine_reg0 <= 36'sb11010011100010011100011011110100111;
            sine_reg0   <= 36'sb10010000001011011101010100001011101;
        end
        391: begin
            cosine_reg0 <= 36'sb11010011010100010001100000110001101;
            sine_reg0   <= 36'sb10010000100000001101110000001111000;
        end
        392: begin
            cosine_reg0 <= 36'sb11010011000110000100100011011000000;
            sine_reg0   <= 36'sb10010000110100111100110011001001100;
        end
        393: begin
            cosine_reg0 <= 36'sb11010010110111110101100011110000101;
            sine_reg0   <= 36'sb10010001001001101010011100101110101;
        end
        394: begin
            cosine_reg0 <= 36'sb11010010101001100100100010000100011;
            sine_reg0   <= 36'sb10010001011110010110101100110001010;
        end
        395: begin
            cosine_reg0 <= 36'sb11010010011011010001011110011100001;
            sine_reg0   <= 36'sb10010001110011000001100011000100111;
        end
        396: begin
            cosine_reg0 <= 36'sb11010010001100111100011001000000100;
            sine_reg0   <= 36'sb10010010000111101010111111011100110;
        end
        397: begin
            cosine_reg0 <= 36'sb11010001111110100101010001111010011;
            sine_reg0   <= 36'sb10010010011100010011000001101011111;
        end
        398: begin
            cosine_reg0 <= 36'sb11010001110000001100001001010010101;
            sine_reg0   <= 36'sb10010010110000111001101001100101110;
        end
        399: begin
            cosine_reg0 <= 36'sb11010001100001110000111111010010010;
            sine_reg0   <= 36'sb10010011000101011110110110111101101;
        end
        400: begin
            cosine_reg0 <= 36'sb11010001010011010011110100000010001;
            sine_reg0   <= 36'sb10010011011010000010101001100110111;
        end
        401: begin
            cosine_reg0 <= 36'sb11010001000100110100100111101011000;
            sine_reg0   <= 36'sb10010011101110100101000001010100101;
        end
        402: begin
            cosine_reg0 <= 36'sb11010000110110010011011010010101111;
            sine_reg0   <= 36'sb10010100000011000101111101111010011;
        end
        403: begin
            cosine_reg0 <= 36'sb11010000100111110000001100001011111;
            sine_reg0   <= 36'sb10010100010111100101011111001011011;
        end
        404: begin
            cosine_reg0 <= 36'sb11010000011001001010111101010101110;
            sine_reg0   <= 36'sb10010100101100000011100100111011000;
        end
        405: begin
            cosine_reg0 <= 36'sb11010000001010100011101101111100101;
            sine_reg0   <= 36'sb10010101000000100000001110111100101;
        end
        406: begin
            cosine_reg0 <= 36'sb11001111111011111010011110001001100;
            sine_reg0   <= 36'sb10010101010100111011011101000011110;
        end
        407: begin
            cosine_reg0 <= 36'sb11001111101101001111001110000101010;
            sine_reg0   <= 36'sb10010101101001010101001111000011101;
        end
        408: begin
            cosine_reg0 <= 36'sb11001111011110100001111101111001010;
            sine_reg0   <= 36'sb10010101111101101101100100101111110;
        end
        409: begin
            cosine_reg0 <= 36'sb11001111001111110010101101101110010;
            sine_reg0   <= 36'sb10010110010010000100011101111011100;
        end
        410: begin
            cosine_reg0 <= 36'sb11001111000001000001011101101101100;
            sine_reg0   <= 36'sb10010110100110011001111010011010011;
        end
        411: begin
            cosine_reg0 <= 36'sb11001110110010001110001110000000001;
            sine_reg0   <= 36'sb10010110111010101101111001111111110;
        end
        412: begin
            cosine_reg0 <= 36'sb11001110100011011000111110101111010;
            sine_reg0   <= 36'sb10010111001111000000011100011111010;
        end
        413: begin
            cosine_reg0 <= 36'sb11001110010100100001110000000011111;
            sine_reg0   <= 36'sb10010111100011010001100001101100001;
        end
        414: begin
            cosine_reg0 <= 36'sb11001110000101101000100010000111011;
            sine_reg0   <= 36'sb10010111110111100001001001011010000;
        end
        415: begin
            cosine_reg0 <= 36'sb11001101110110101101010101000010111;
            sine_reg0   <= 36'sb10011000001011101111010011011100100;
        end
        416: begin
            cosine_reg0 <= 36'sb11001101100111110000001000111111100;
            sine_reg0   <= 36'sb10011000011111111011111111100111000;
        end
        417: begin
            cosine_reg0 <= 36'sb11001101011000110000111110000110100;
            sine_reg0   <= 36'sb10011000110100000111001101101101000;
        end
        418: begin
            cosine_reg0 <= 36'sb11001101001001101111110100100001010;
            sine_reg0   <= 36'sb10011001001000010000111101100010010;
        end
        419: begin
            cosine_reg0 <= 36'sb11001100111010101100101100011000111;
            sine_reg0   <= 36'sb10011001011100011001001110111010001;
        end
        420: begin
            cosine_reg0 <= 36'sb11001100101011100111100101110110101;
            sine_reg0   <= 36'sb10011001110000100000000001101000011;
        end
        421: begin
            cosine_reg0 <= 36'sb11001100011100100000100001000100000;
            sine_reg0   <= 36'sb10011010000100100101010101100000011;
        end
        422: begin
            cosine_reg0 <= 36'sb11001100001101010111011110001010001;
            sine_reg0   <= 36'sb10011010011000101001001010010110000;
        end
        423: begin
            cosine_reg0 <= 36'sb11001011111110001100011101010010011;
            sine_reg0   <= 36'sb10011010101100101011011111111100101;
        end
        424: begin
            cosine_reg0 <= 36'sb11001011101110111111011110100110001;
            sine_reg0   <= 36'sb10011011000000101100010110001000001;
        end
        425: begin
            cosine_reg0 <= 36'sb11001011011111110000100010001110111;
            sine_reg0   <= 36'sb10011011010100101011101100101100000;
        end
        426: begin
            cosine_reg0 <= 36'sb11001011010000011111101000010101111;
            sine_reg0   <= 36'sb10011011101000101001100011011100000;
        end
        427: begin
            cosine_reg0 <= 36'sb11001011000001001100110001000100100;
            sine_reg0   <= 36'sb10011011111100100101111010001011110;
        end
        428: begin
            cosine_reg0 <= 36'sb11001010110001110111111100100100011;
            sine_reg0   <= 36'sb10011100010000100000110000101110111;
        end
        429: begin
            cosine_reg0 <= 36'sb11001010100010100001001010111110110;
            sine_reg0   <= 36'sb10011100100100011010000110111001011;
        end
        430: begin
            cosine_reg0 <= 36'sb11001010010011001000011100011101010;
            sine_reg0   <= 36'sb10011100111000010001111100011110101;
        end
        431: begin
            cosine_reg0 <= 36'sb11001010000011101101110001001001011;
            sine_reg0   <= 36'sb10011101001100001000010001010010101;
        end
        432: begin
            cosine_reg0 <= 36'sb11001001110100010001001001001100100;
            sine_reg0   <= 36'sb10011101011111111101000101001000111;
        end
        433: begin
            cosine_reg0 <= 36'sb11001001100100110010100100110000010;
            sine_reg0   <= 36'sb10011101110011110000010111110101100;
        end
        434: begin
            cosine_reg0 <= 36'sb11001001010101010010000011111110001;
            sine_reg0   <= 36'sb10011110000111100010001001001100000;
        end
        435: begin
            cosine_reg0 <= 36'sb11001001000101101111100110111111101;
            sine_reg0   <= 36'sb10011110011011010010011001000000010;
        end
        436: begin
            cosine_reg0 <= 36'sb11001000110110001011001101111110100;
            sine_reg0   <= 36'sb10011110101111000001000111000110001;
        end
        437: begin
            cosine_reg0 <= 36'sb11001000100110100100111001000100011;
            sine_reg0   <= 36'sb10011111000010101110010011010001011;
        end
        438: begin
            cosine_reg0 <= 36'sb11001000010110111100101000011010101;
            sine_reg0   <= 36'sb10011111010110011001111101010101111;
        end
        439: begin
            cosine_reg0 <= 36'sb11001000000111010010011100001011001;
            sine_reg0   <= 36'sb10011111101010000100000101000111100;
        end
        440: begin
            cosine_reg0 <= 36'sb11000111110111100110010100011111011;
            sine_reg0   <= 36'sb10011111111101101100101010011010001;
        end
        441: begin
            cosine_reg0 <= 36'sb11000111100111111000010001100001001;
            sine_reg0   <= 36'sb10100000010001010011101101000001101;
        end
        442: begin
            cosine_reg0 <= 36'sb11000111011000001000010011011010001;
            sine_reg0   <= 36'sb10100000100100111001001100110001111;
        end
        443: begin
            cosine_reg0 <= 36'sb11000111001000010110011010010100001;
            sine_reg0   <= 36'sb10100000111000011101001001011110110;
        end
        444: begin
            cosine_reg0 <= 36'sb11000110111000100010100110011000101;
            sine_reg0   <= 36'sb10100001001011111111100010111100011;
        end
        445: begin
            cosine_reg0 <= 36'sb11000110101000101100110111110001100;
            sine_reg0   <= 36'sb10100001011111100000011000111110100;
        end
        446: begin
            cosine_reg0 <= 36'sb11000110011000110101001110101000101;
            sine_reg0   <= 36'sb10100001110010111111101011011001010;
        end
        447: begin
            cosine_reg0 <= 36'sb11000110001000111011101011000111110;
            sine_reg0   <= 36'sb10100010000110011101011010000000100;
        end
        448: begin
            cosine_reg0 <= 36'sb11000101111001000000001101011000100;
            sine_reg0   <= 36'sb10100010011001111001100100101000010;
        end
        449: begin
            cosine_reg0 <= 36'sb11000101101001000010110101100101000;
            sine_reg0   <= 36'sb10100010101101010100001011000100100;
        end
        450: begin
            cosine_reg0 <= 36'sb11000101011001000011100011110110111;
            sine_reg0   <= 36'sb10100011000000101101001101001001010;
        end
        451: begin
            cosine_reg0 <= 36'sb11000101001001000010011000011000000;
            sine_reg0   <= 36'sb10100011010100000100101010101010101;
        end
        452: begin
            cosine_reg0 <= 36'sb11000100111000111111010011010010011;
            sine_reg0   <= 36'sb10100011100111011010100011011100101;
        end
        453: begin
            cosine_reg0 <= 36'sb11000100101000111010010100101111110;
            sine_reg0   <= 36'sb10100011111010101110110111010011011;
        end
        454: begin
            cosine_reg0 <= 36'sb11000100011000110011011100111010001;
            sine_reg0   <= 36'sb10100100001110000001100110000011000;
        end
        455: begin
            cosine_reg0 <= 36'sb11000100001000101010101011111011100;
            sine_reg0   <= 36'sb10100100100001010010101111011111011;
        end
        456: begin
            cosine_reg0 <= 36'sb11000011111000100000000001111101110;
            sine_reg0   <= 36'sb10100100110100100010010011011100110;
        end
        457: begin
            cosine_reg0 <= 36'sb11000011101000010011011111001010110;
            sine_reg0   <= 36'sb10100101000111110000010001101111011;
        end
        458: begin
            cosine_reg0 <= 36'sb11000011011000000101000011101100110;
            sine_reg0   <= 36'sb10100101011010111100101010001011001;
        end
        459: begin
            cosine_reg0 <= 36'sb11000011000111110100101111101101100;
            sine_reg0   <= 36'sb10100101101110000111011100100100011;
        end
        460: begin
            cosine_reg0 <= 36'sb11000010110111100010100011010111010;
            sine_reg0   <= 36'sb10100110000001010000101000101111010;
        end
        461: begin
            cosine_reg0 <= 36'sb11000010100111001110011110110011110;
            sine_reg0   <= 36'sb10100110010100011000001110100000000;
        end
        462: begin
            cosine_reg0 <= 36'sb11000010010110111000100010001101011;
            sine_reg0   <= 36'sb10100110100111011110001101101010110;
        end
        463: begin
            cosine_reg0 <= 36'sb11000010000110100000101101101110000;
            sine_reg0   <= 36'sb10100110111010100010100110000011101;
        end
        464: begin
            cosine_reg0 <= 36'sb11000001110110000111000001011111111;
            sine_reg0   <= 36'sb10100111001101100101010111011111000;
        end
        465: begin
            cosine_reg0 <= 36'sb11000001100101101011011101101101000;
            sine_reg0   <= 36'sb10100111100000100110100001110001001;
        end
        466: begin
            cosine_reg0 <= 36'sb11000001010101001110000010011111101;
            sine_reg0   <= 36'sb10100111110011100110000100101110011;
        end
        467: begin
            cosine_reg0 <= 36'sb11000001000100101110110000000001110;
            sine_reg0   <= 36'sb10101000000110100100000000001010110;
        end
        468: begin
            cosine_reg0 <= 36'sb11000000110100001101100110011101101;
            sine_reg0   <= 36'sb10101000011001100000010011111010110;
        end
        469: begin
            cosine_reg0 <= 36'sb11000000100011101010100101111101011;
            sine_reg0   <= 36'sb10101000101100011010111111110010101;
        end
        470: begin
            cosine_reg0 <= 36'sb11000000010011000101101110101011011;
            sine_reg0   <= 36'sb10101000111111010100000011100110110;
        end
        471: begin
            cosine_reg0 <= 36'sb11000000000010011111000000110001101;
            sine_reg0   <= 36'sb10101001010010001011011111001011011;
        end
        472: begin
            cosine_reg0 <= 36'sb10111111110001110110011100011010101;
            sine_reg0   <= 36'sb10101001100101000001010010010101000;
        end
        473: begin
            cosine_reg0 <= 36'sb10111111100001001100000001110000100;
            sine_reg0   <= 36'sb10101001110111110101011100111000000;
        end
        474: begin
            cosine_reg0 <= 36'sb10111111010000011111110000111101011;
            sine_reg0   <= 36'sb10101010001010100111111110101000101;
        end
        475: begin
            cosine_reg0 <= 36'sb10111110111111110001101010001011111;
            sine_reg0   <= 36'sb10101010011101011000110111011011011;
        end
        476: begin
            cosine_reg0 <= 36'sb10111110101111000001101101100110000;
            sine_reg0   <= 36'sb10101010110000001000000111000100101;
        end
        477: begin
            cosine_reg0 <= 36'sb10111110011110001111111011010110010;
            sine_reg0   <= 36'sb10101011000010110101101101011000111;
        end
        478: begin
            cosine_reg0 <= 36'sb10111110001101011100010011100111000;
            sine_reg0   <= 36'sb10101011010101100001101010001100101;
        end
        479: begin
            cosine_reg0 <= 36'sb10111101111100100110110110100010100;
            sine_reg0   <= 36'sb10101011101000001011111101010100010;
        end
        480: begin
            cosine_reg0 <= 36'sb10111101101011101111100100010011010;
            sine_reg0   <= 36'sb10101011111010110100100110100100011;
        end
        481: begin
            cosine_reg0 <= 36'sb10111101011010110110011101000011100;
            sine_reg0   <= 36'sb10101100001101011011100101110001010;
        end
        482: begin
            cosine_reg0 <= 36'sb10111101001001111011100000111101111;
            sine_reg0   <= 36'sb10101100100000000000111010101111101;
        end
        483: begin
            cosine_reg0 <= 36'sb10111100111000111110110000001100101;
            sine_reg0   <= 36'sb10101100110010100100100101010100000;
        end
        484: begin
            cosine_reg0 <= 36'sb10111100101000000000001010111010011;
            sine_reg0   <= 36'sb10101101000101000110100101010010111;
        end
        485: begin
            cosine_reg0 <= 36'sb10111100010110111111110001010001100;
            sine_reg0   <= 36'sb10101101010111100110111010100000110;
        end
        486: begin
            cosine_reg0 <= 36'sb10111100000101111101100011011100011;
            sine_reg0   <= 36'sb10101101101010000101100100110010011;
        end
        487: begin
            cosine_reg0 <= 36'sb10111011110100111001100001100101110;
            sine_reg0   <= 36'sb10101101111100100010100011111100010;
        end
        488: begin
            cosine_reg0 <= 36'sb10111011100011110011101011111000000;
            sine_reg0   <= 36'sb10101110001110111101110111110011001;
        end
        489: begin
            cosine_reg0 <= 36'sb10111011010010101100000010011101110;
            sine_reg0   <= 36'sb10101110100001010111100000001011011;
        end
        490: begin
            cosine_reg0 <= 36'sb10111011000001100010100101100001011;
            sine_reg0   <= 36'sb10101110110011101111011100111001111;
        end
        491: begin
            cosine_reg0 <= 36'sb10111010110000010111010101001101110;
            sine_reg0   <= 36'sb10101111000110000101101101110011001;
        end
        492: begin
            cosine_reg0 <= 36'sb10111010011111001010010001101101001;
            sine_reg0   <= 36'sb10101111011000011010010010101100000;
        end
        493: begin
            cosine_reg0 <= 36'sb10111010001101111011011011001010100;
            sine_reg0   <= 36'sb10101111101010101101001011011001001;
        end
        494: begin
            cosine_reg0 <= 36'sb10111001111100101010110001110000001;
            sine_reg0   <= 36'sb10101111111100111110010111101111001;
        end
        495: begin
            cosine_reg0 <= 36'sb10111001101011011000010101101000111;
            sine_reg0   <= 36'sb10110000001111001101110111100010110;
        end
        496: begin
            cosine_reg0 <= 36'sb10111001011010000100000110111111011;
            sine_reg0   <= 36'sb10110000100001011011101010101000111;
        end
        497: begin
            cosine_reg0 <= 36'sb10111001001000101110000101111110011;
            sine_reg0   <= 36'sb10110000110011100111110000110110001;
        end
        498: begin
            cosine_reg0 <= 36'sb10111000110111010110010010110000011;
            sine_reg0   <= 36'sb10110001000101110010001001111111010;
        end
        499: begin
            cosine_reg0 <= 36'sb10111000100101111100101101100000010;
            sine_reg0   <= 36'sb10110001010111111010110101111001010;
        end
        500: begin
            cosine_reg0 <= 36'sb10111000010100100001010110011000101;
            sine_reg0   <= 36'sb10110001101010000001110100011000110;
        end
        501: begin
            cosine_reg0 <= 36'sb10111000000011000100001101100100011;
            sine_reg0   <= 36'sb10110001111100000111000101010010110;
        end
        502: begin
            cosine_reg0 <= 36'sb10110111110001100101010011001110010;
            sine_reg0   <= 36'sb10110010001110001010101000011011111;
        end
        503: begin
            cosine_reg0 <= 36'sb10110111100000000100100111100000111;
            sine_reg0   <= 36'sb10110010100000001100011101101001001;
        end
        504: begin
            cosine_reg0 <= 36'sb10110111001110100010001010100111010;
            sine_reg0   <= 36'sb10110010110010001100100100101111011;
        end
        505: begin
            cosine_reg0 <= 36'sb10110110111100111101111100101100001;
            sine_reg0   <= 36'sb10110011000100001010111101100011101;
        end
        506: begin
            cosine_reg0 <= 36'sb10110110101011010111111101111010010;
            sine_reg0   <= 36'sb10110011010110000111100111111010100;
        end
        507: begin
            cosine_reg0 <= 36'sb10110110011001110000001110011100101;
            sine_reg0   <= 36'sb10110011101000000010100011101001001;
        end
        508: begin
            cosine_reg0 <= 36'sb10110110001000000110101110011110000;
            sine_reg0   <= 36'sb10110011111001111011110000100100100;
        end
        509: begin
            cosine_reg0 <= 36'sb10110101110110011011011110001001010;
            sine_reg0   <= 36'sb10110100001011110011001110100001011;
        end
        510: begin
            cosine_reg0 <= 36'sb10110101100100101110011101101001011;
            sine_reg0   <= 36'sb10110100011101101000111101010101000;
        end
        511: begin
            cosine_reg0 <= 36'sb10110101010010111111101101001001010;
            sine_reg0   <= 36'sb10110100101111011100111100110100001;
        end
        512: begin
            cosine_reg0 <= 36'sb10110101000001001111001100110011111;
            sine_reg0   <= 36'sb10110101000001001111001100110011111;
        end
        513: begin
            cosine_reg0 <= 36'sb10110100101111011100111100110100001;
            sine_reg0   <= 36'sb10110101010010111111101101001001010;
        end
        514: begin
            cosine_reg0 <= 36'sb10110100011101101000111101010101000;
            sine_reg0   <= 36'sb10110101100100101110011101101001011;
        end
        515: begin
            cosine_reg0 <= 36'sb10110100001011110011001110100001011;
            sine_reg0   <= 36'sb10110101110110011011011110001001010;
        end
        516: begin
            cosine_reg0 <= 36'sb10110011111001111011110000100100100;
            sine_reg0   <= 36'sb10110110001000000110101110011110000;
        end
        517: begin
            cosine_reg0 <= 36'sb10110011101000000010100011101001001;
            sine_reg0   <= 36'sb10110110011001110000001110011100101;
        end
        518: begin
            cosine_reg0 <= 36'sb10110011010110000111100111111010100;
            sine_reg0   <= 36'sb10110110101011010111111101111010010;
        end
        519: begin
            cosine_reg0 <= 36'sb10110011000100001010111101100011101;
            sine_reg0   <= 36'sb10110110111100111101111100101100001;
        end
        520: begin
            cosine_reg0 <= 36'sb10110010110010001100100100101111011;
            sine_reg0   <= 36'sb10110111001110100010001010100111010;
        end
        521: begin
            cosine_reg0 <= 36'sb10110010100000001100011101101001001;
            sine_reg0   <= 36'sb10110111100000000100100111100000111;
        end
        522: begin
            cosine_reg0 <= 36'sb10110010001110001010101000011011111;
            sine_reg0   <= 36'sb10110111110001100101010011001110010;
        end
        523: begin
            cosine_reg0 <= 36'sb10110001111100000111000101010010110;
            sine_reg0   <= 36'sb10111000000011000100001101100100011;
        end
        524: begin
            cosine_reg0 <= 36'sb10110001101010000001110100011000110;
            sine_reg0   <= 36'sb10111000010100100001010110011000101;
        end
        525: begin
            cosine_reg0 <= 36'sb10110001010111111010110101111001010;
            sine_reg0   <= 36'sb10111000100101111100101101100000010;
        end
        526: begin
            cosine_reg0 <= 36'sb10110001000101110010001001111111010;
            sine_reg0   <= 36'sb10111000110111010110010010110000011;
        end
        527: begin
            cosine_reg0 <= 36'sb10110000110011100111110000110110001;
            sine_reg0   <= 36'sb10111001001000101110000101111110011;
        end
        528: begin
            cosine_reg0 <= 36'sb10110000100001011011101010101000111;
            sine_reg0   <= 36'sb10111001011010000100000110111111011;
        end
        529: begin
            cosine_reg0 <= 36'sb10110000001111001101110111100010110;
            sine_reg0   <= 36'sb10111001101011011000010101101000111;
        end
        530: begin
            cosine_reg0 <= 36'sb10101111111100111110010111101111001;
            sine_reg0   <= 36'sb10111001111100101010110001110000001;
        end
        531: begin
            cosine_reg0 <= 36'sb10101111101010101101001011011001001;
            sine_reg0   <= 36'sb10111010001101111011011011001010100;
        end
        532: begin
            cosine_reg0 <= 36'sb10101111011000011010010010101100000;
            sine_reg0   <= 36'sb10111010011111001010010001101101001;
        end
        533: begin
            cosine_reg0 <= 36'sb10101111000110000101101101110011001;
            sine_reg0   <= 36'sb10111010110000010111010101001101110;
        end
        534: begin
            cosine_reg0 <= 36'sb10101110110011101111011100111001111;
            sine_reg0   <= 36'sb10111011000001100010100101100001011;
        end
        535: begin
            cosine_reg0 <= 36'sb10101110100001010111100000001011011;
            sine_reg0   <= 36'sb10111011010010101100000010011101110;
        end
        536: begin
            cosine_reg0 <= 36'sb10101110001110111101110111110011001;
            sine_reg0   <= 36'sb10111011100011110011101011111000000;
        end
        537: begin
            cosine_reg0 <= 36'sb10101101111100100010100011111100010;
            sine_reg0   <= 36'sb10111011110100111001100001100101110;
        end
        538: begin
            cosine_reg0 <= 36'sb10101101101010000101100100110010011;
            sine_reg0   <= 36'sb10111100000101111101100011011100011;
        end
        539: begin
            cosine_reg0 <= 36'sb10101101010111100110111010100000110;
            sine_reg0   <= 36'sb10111100010110111111110001010001100;
        end
        540: begin
            cosine_reg0 <= 36'sb10101101000101000110100101010010111;
            sine_reg0   <= 36'sb10111100101000000000001010111010011;
        end
        541: begin
            cosine_reg0 <= 36'sb10101100110010100100100101010100000;
            sine_reg0   <= 36'sb10111100111000111110110000001100101;
        end
        542: begin
            cosine_reg0 <= 36'sb10101100100000000000111010101111101;
            sine_reg0   <= 36'sb10111101001001111011100000111101111;
        end
        543: begin
            cosine_reg0 <= 36'sb10101100001101011011100101110001010;
            sine_reg0   <= 36'sb10111101011010110110011101000011100;
        end
        544: begin
            cosine_reg0 <= 36'sb10101011111010110100100110100100011;
            sine_reg0   <= 36'sb10111101101011101111100100010011010;
        end
        545: begin
            cosine_reg0 <= 36'sb10101011101000001011111101010100010;
            sine_reg0   <= 36'sb10111101111100100110110110100010100;
        end
        546: begin
            cosine_reg0 <= 36'sb10101011010101100001101010001100101;
            sine_reg0   <= 36'sb10111110001101011100010011100111000;
        end
        547: begin
            cosine_reg0 <= 36'sb10101011000010110101101101011000111;
            sine_reg0   <= 36'sb10111110011110001111111011010110010;
        end
        548: begin
            cosine_reg0 <= 36'sb10101010110000001000000111000100101;
            sine_reg0   <= 36'sb10111110101111000001101101100110000;
        end
        549: begin
            cosine_reg0 <= 36'sb10101010011101011000110111011011011;
            sine_reg0   <= 36'sb10111110111111110001101010001011111;
        end
        550: begin
            cosine_reg0 <= 36'sb10101010001010100111111110101000101;
            sine_reg0   <= 36'sb10111111010000011111110000111101011;
        end
        551: begin
            cosine_reg0 <= 36'sb10101001110111110101011100111000000;
            sine_reg0   <= 36'sb10111111100001001100000001110000100;
        end
        552: begin
            cosine_reg0 <= 36'sb10101001100101000001010010010101000;
            sine_reg0   <= 36'sb10111111110001110110011100011010101;
        end
        553: begin
            cosine_reg0 <= 36'sb10101001010010001011011111001011011;
            sine_reg0   <= 36'sb11000000000010011111000000110001101;
        end
        554: begin
            cosine_reg0 <= 36'sb10101000111111010100000011100110110;
            sine_reg0   <= 36'sb11000000010011000101101110101011011;
        end
        555: begin
            cosine_reg0 <= 36'sb10101000101100011010111111110010101;
            sine_reg0   <= 36'sb11000000100011101010100101111101011;
        end
        556: begin
            cosine_reg0 <= 36'sb10101000011001100000010011111010110;
            sine_reg0   <= 36'sb11000000110100001101100110011101101;
        end
        557: begin
            cosine_reg0 <= 36'sb10101000000110100100000000001010110;
            sine_reg0   <= 36'sb11000001000100101110110000000001110;
        end
        558: begin
            cosine_reg0 <= 36'sb10100111110011100110000100101110011;
            sine_reg0   <= 36'sb11000001010101001110000010011111101;
        end
        559: begin
            cosine_reg0 <= 36'sb10100111100000100110100001110001001;
            sine_reg0   <= 36'sb11000001100101101011011101101101000;
        end
        560: begin
            cosine_reg0 <= 36'sb10100111001101100101010111011111000;
            sine_reg0   <= 36'sb11000001110110000111000001011111111;
        end
        561: begin
            cosine_reg0 <= 36'sb10100110111010100010100110000011101;
            sine_reg0   <= 36'sb11000010000110100000101101101110000;
        end
        562: begin
            cosine_reg0 <= 36'sb10100110100111011110001101101010110;
            sine_reg0   <= 36'sb11000010010110111000100010001101011;
        end
        563: begin
            cosine_reg0 <= 36'sb10100110010100011000001110100000000;
            sine_reg0   <= 36'sb11000010100111001110011110110011110;
        end
        564: begin
            cosine_reg0 <= 36'sb10100110000001010000101000101111010;
            sine_reg0   <= 36'sb11000010110111100010100011010111010;
        end
        565: begin
            cosine_reg0 <= 36'sb10100101101110000111011100100100011;
            sine_reg0   <= 36'sb11000011000111110100101111101101100;
        end
        566: begin
            cosine_reg0 <= 36'sb10100101011010111100101010001011001;
            sine_reg0   <= 36'sb11000011011000000101000011101100110;
        end
        567: begin
            cosine_reg0 <= 36'sb10100101000111110000010001101111011;
            sine_reg0   <= 36'sb11000011101000010011011111001010110;
        end
        568: begin
            cosine_reg0 <= 36'sb10100100110100100010010011011100110;
            sine_reg0   <= 36'sb11000011111000100000000001111101110;
        end
        569: begin
            cosine_reg0 <= 36'sb10100100100001010010101111011111011;
            sine_reg0   <= 36'sb11000100001000101010101011111011100;
        end
        570: begin
            cosine_reg0 <= 36'sb10100100001110000001100110000011000;
            sine_reg0   <= 36'sb11000100011000110011011100111010001;
        end
        571: begin
            cosine_reg0 <= 36'sb10100011111010101110110111010011011;
            sine_reg0   <= 36'sb11000100101000111010010100101111110;
        end
        572: begin
            cosine_reg0 <= 36'sb10100011100111011010100011011100101;
            sine_reg0   <= 36'sb11000100111000111111010011010010011;
        end
        573: begin
            cosine_reg0 <= 36'sb10100011010100000100101010101010101;
            sine_reg0   <= 36'sb11000101001001000010011000011000000;
        end
        574: begin
            cosine_reg0 <= 36'sb10100011000000101101001101001001010;
            sine_reg0   <= 36'sb11000101011001000011100011110110111;
        end
        575: begin
            cosine_reg0 <= 36'sb10100010101101010100001011000100100;
            sine_reg0   <= 36'sb11000101101001000010110101100101000;
        end
        576: begin
            cosine_reg0 <= 36'sb10100010011001111001100100101000010;
            sine_reg0   <= 36'sb11000101111001000000001101011000100;
        end
        577: begin
            cosine_reg0 <= 36'sb10100010000110011101011010000000100;
            sine_reg0   <= 36'sb11000110001000111011101011000111110;
        end
        578: begin
            cosine_reg0 <= 36'sb10100001110010111111101011011001010;
            sine_reg0   <= 36'sb11000110011000110101001110101000101;
        end
        579: begin
            cosine_reg0 <= 36'sb10100001011111100000011000111110100;
            sine_reg0   <= 36'sb11000110101000101100110111110001100;
        end
        580: begin
            cosine_reg0 <= 36'sb10100001001011111111100010111100011;
            sine_reg0   <= 36'sb11000110111000100010100110011000101;
        end
        581: begin
            cosine_reg0 <= 36'sb10100000111000011101001001011110110;
            sine_reg0   <= 36'sb11000111001000010110011010010100001;
        end
        582: begin
            cosine_reg0 <= 36'sb10100000100100111001001100110001111;
            sine_reg0   <= 36'sb11000111011000001000010011011010001;
        end
        583: begin
            cosine_reg0 <= 36'sb10100000010001010011101101000001101;
            sine_reg0   <= 36'sb11000111100111111000010001100001001;
        end
        584: begin
            cosine_reg0 <= 36'sb10011111111101101100101010011010001;
            sine_reg0   <= 36'sb11000111110111100110010100011111011;
        end
        585: begin
            cosine_reg0 <= 36'sb10011111101010000100000101000111100;
            sine_reg0   <= 36'sb11001000000111010010011100001011001;
        end
        586: begin
            cosine_reg0 <= 36'sb10011111010110011001111101010101111;
            sine_reg0   <= 36'sb11001000010110111100101000011010101;
        end
        587: begin
            cosine_reg0 <= 36'sb10011111000010101110010011010001011;
            sine_reg0   <= 36'sb11001000100110100100111001000100011;
        end
        588: begin
            cosine_reg0 <= 36'sb10011110101111000001000111000110001;
            sine_reg0   <= 36'sb11001000110110001011001101111110100;
        end
        589: begin
            cosine_reg0 <= 36'sb10011110011011010010011001000000010;
            sine_reg0   <= 36'sb11001001000101101111100110111111101;
        end
        590: begin
            cosine_reg0 <= 36'sb10011110000111100010001001001100000;
            sine_reg0   <= 36'sb11001001010101010010000011111110001;
        end
        591: begin
            cosine_reg0 <= 36'sb10011101110011110000010111110101100;
            sine_reg0   <= 36'sb11001001100100110010100100110000010;
        end
        592: begin
            cosine_reg0 <= 36'sb10011101011111111101000101001000111;
            sine_reg0   <= 36'sb11001001110100010001001001001100100;
        end
        593: begin
            cosine_reg0 <= 36'sb10011101001100001000010001010010101;
            sine_reg0   <= 36'sb11001010000011101101110001001001011;
        end
        594: begin
            cosine_reg0 <= 36'sb10011100111000010001111100011110101;
            sine_reg0   <= 36'sb11001010010011001000011100011101010;
        end
        595: begin
            cosine_reg0 <= 36'sb10011100100100011010000110111001011;
            sine_reg0   <= 36'sb11001010100010100001001010111110110;
        end
        596: begin
            cosine_reg0 <= 36'sb10011100010000100000110000101110111;
            sine_reg0   <= 36'sb11001010110001110111111100100100011;
        end
        597: begin
            cosine_reg0 <= 36'sb10011011111100100101111010001011110;
            sine_reg0   <= 36'sb11001011000001001100110001000100100;
        end
        598: begin
            cosine_reg0 <= 36'sb10011011101000101001100011011100000;
            sine_reg0   <= 36'sb11001011010000011111101000010101111;
        end
        599: begin
            cosine_reg0 <= 36'sb10011011010100101011101100101100000;
            sine_reg0   <= 36'sb11001011011111110000100010001110111;
        end
        600: begin
            cosine_reg0 <= 36'sb10011011000000101100010110001000001;
            sine_reg0   <= 36'sb11001011101110111111011110100110001;
        end
        601: begin
            cosine_reg0 <= 36'sb10011010101100101011011111111100101;
            sine_reg0   <= 36'sb11001011111110001100011101010010011;
        end
        602: begin
            cosine_reg0 <= 36'sb10011010011000101001001010010110000;
            sine_reg0   <= 36'sb11001100001101010111011110001010001;
        end
        603: begin
            cosine_reg0 <= 36'sb10011010000100100101010101100000011;
            sine_reg0   <= 36'sb11001100011100100000100001000100000;
        end
        604: begin
            cosine_reg0 <= 36'sb10011001110000100000000001101000011;
            sine_reg0   <= 36'sb11001100101011100111100101110110101;
        end
        605: begin
            cosine_reg0 <= 36'sb10011001011100011001001110111010001;
            sine_reg0   <= 36'sb11001100111010101100101100011000111;
        end
        606: begin
            cosine_reg0 <= 36'sb10011001001000010000111101100010010;
            sine_reg0   <= 36'sb11001101001001101111110100100001010;
        end
        607: begin
            cosine_reg0 <= 36'sb10011000110100000111001101101101000;
            sine_reg0   <= 36'sb11001101011000110000111110000110100;
        end
        608: begin
            cosine_reg0 <= 36'sb10011000011111111011111111100111000;
            sine_reg0   <= 36'sb11001101100111110000001000111111100;
        end
        609: begin
            cosine_reg0 <= 36'sb10011000001011101111010011011100100;
            sine_reg0   <= 36'sb11001101110110101101010101000010111;
        end
        610: begin
            cosine_reg0 <= 36'sb10010111110111100001001001011010000;
            sine_reg0   <= 36'sb11001110000101101000100010000111011;
        end
        611: begin
            cosine_reg0 <= 36'sb10010111100011010001100001101100001;
            sine_reg0   <= 36'sb11001110010100100001110000000011111;
        end
        612: begin
            cosine_reg0 <= 36'sb10010111001111000000011100011111010;
            sine_reg0   <= 36'sb11001110100011011000111110101111010;
        end
        613: begin
            cosine_reg0 <= 36'sb10010110111010101101111001111111110;
            sine_reg0   <= 36'sb11001110110010001110001110000000001;
        end
        614: begin
            cosine_reg0 <= 36'sb10010110100110011001111010011010011;
            sine_reg0   <= 36'sb11001111000001000001011101101101100;
        end
        615: begin
            cosine_reg0 <= 36'sb10010110010010000100011101111011100;
            sine_reg0   <= 36'sb11001111001111110010101101101110010;
        end
        616: begin
            cosine_reg0 <= 36'sb10010101111101101101100100101111110;
            sine_reg0   <= 36'sb11001111011110100001111101111001010;
        end
        617: begin
            cosine_reg0 <= 36'sb10010101101001010101001111000011101;
            sine_reg0   <= 36'sb11001111101101001111001110000101010;
        end
        618: begin
            cosine_reg0 <= 36'sb10010101010100111011011101000011110;
            sine_reg0   <= 36'sb11001111111011111010011110001001100;
        end
        619: begin
            cosine_reg0 <= 36'sb10010101000000100000001110111100101;
            sine_reg0   <= 36'sb11010000001010100011101101111100101;
        end
        620: begin
            cosine_reg0 <= 36'sb10010100101100000011100100111011000;
            sine_reg0   <= 36'sb11010000011001001010111101010101110;
        end
        621: begin
            cosine_reg0 <= 36'sb10010100010111100101011111001011011;
            sine_reg0   <= 36'sb11010000100111110000001100001011111;
        end
        622: begin
            cosine_reg0 <= 36'sb10010100000011000101111101111010011;
            sine_reg0   <= 36'sb11010000110110010011011010010101111;
        end
        623: begin
            cosine_reg0 <= 36'sb10010011101110100101000001010100101;
            sine_reg0   <= 36'sb11010001000100110100100111101011000;
        end
        624: begin
            cosine_reg0 <= 36'sb10010011011010000010101001100110111;
            sine_reg0   <= 36'sb11010001010011010011110100000010001;
        end
        625: begin
            cosine_reg0 <= 36'sb10010011000101011110110110111101101;
            sine_reg0   <= 36'sb11010001100001110000111111010010010;
        end
        626: begin
            cosine_reg0 <= 36'sb10010010110000111001101001100101110;
            sine_reg0   <= 36'sb11010001110000001100001001010010101;
        end
        627: begin
            cosine_reg0 <= 36'sb10010010011100010011000001101011111;
            sine_reg0   <= 36'sb11010001111110100101010001111010011;
        end
        628: begin
            cosine_reg0 <= 36'sb10010010000111101010111111011100110;
            sine_reg0   <= 36'sb11010010001100111100011001000000100;
        end
        629: begin
            cosine_reg0 <= 36'sb10010001110011000001100011000100111;
            sine_reg0   <= 36'sb11010010011011010001011110011100001;
        end
        630: begin
            cosine_reg0 <= 36'sb10010001011110010110101100110001010;
            sine_reg0   <= 36'sb11010010101001100100100010000100011;
        end
        631: begin
            cosine_reg0 <= 36'sb10010001001001101010011100101110101;
            sine_reg0   <= 36'sb11010010110111110101100011110000101;
        end
        632: begin
            cosine_reg0 <= 36'sb10010000110100111100110011001001100;
            sine_reg0   <= 36'sb11010011000110000100100011011000000;
        end
        633: begin
            cosine_reg0 <= 36'sb10010000100000001101110000001111000;
            sine_reg0   <= 36'sb11010011010100010001100000110001101;
        end
        634: begin
            cosine_reg0 <= 36'sb10010000001011011101010100001011101;
            sine_reg0   <= 36'sb11010011100010011100011011110100111;
        end
        635: begin
            cosine_reg0 <= 36'sb10001111110110101011011111001100010;
            sine_reg0   <= 36'sb11010011110000100101010100011000110;
        end
        636: begin
            cosine_reg0 <= 36'sb10001111100001111000010001011101111;
            sine_reg0   <= 36'sb11010011111110101100001010010100111;
        end
        637: begin
            cosine_reg0 <= 36'sb10001111001101000011101011001101000;
            sine_reg0   <= 36'sb11010100001100110000111101100000011;
        end
        638: begin
            cosine_reg0 <= 36'sb10001110111000001101101100100110111;
            sine_reg0   <= 36'sb11010100011010110011101101110010100;
        end
        639: begin
            cosine_reg0 <= 36'sb10001110100011010110010101111000000;
            sine_reg0   <= 36'sb11010100101000110100011011000010110;
        end
        640: begin
            cosine_reg0 <= 36'sb10001110001110011101100111001101011;
            sine_reg0   <= 36'sb11010100110110110011000101001000011;
        end
        641: begin
            cosine_reg0 <= 36'sb10001101111001100011100000110100000;
            sine_reg0   <= 36'sb11010101000100101111101011111010110;
        end
        642: begin
            cosine_reg0 <= 36'sb10001101100100101000000010111000100;
            sine_reg0   <= 36'sb11010101010010101010001111010001010;
        end
        643: begin
            cosine_reg0 <= 36'sb10001101001111101011001101101000001;
            sine_reg0   <= 36'sb11010101100000100010101111000011100;
        end
        644: begin
            cosine_reg0 <= 36'sb10001100111010101101000001001111100;
            sine_reg0   <= 36'sb11010101101110011001001011001000101;
        end
        645: begin
            cosine_reg0 <= 36'sb10001100100101101101011101111011110;
            sine_reg0   <= 36'sb11010101111100001101100011011000010;
        end
        646: begin
            cosine_reg0 <= 36'sb10001100010000101100100011111001110;
            sine_reg0   <= 36'sb11010110001001111111110111101001111;
        end
        647: begin
            cosine_reg0 <= 36'sb10001011111011101010010011010110100;
            sine_reg0   <= 36'sb11010110010111110000000111110100111;
        end
        648: begin
            cosine_reg0 <= 36'sb10001011100110100110101100011110111;
            sine_reg0   <= 36'sb11010110100101011110010011110001000;
        end
        649: begin
            cosine_reg0 <= 36'sb10001011010001100001101111100000000;
            sine_reg0   <= 36'sb11010110110011001010011011010101100;
        end
        650: begin
            cosine_reg0 <= 36'sb10001010111100011011011100100110110;
            sine_reg0   <= 36'sb11010111000000110100011110011010001;
        end
        651: begin
            cosine_reg0 <= 36'sb10001010100111010011110100000000010;
            sine_reg0   <= 36'sb11010111001110011100011100110110010;
        end
        652: begin
            cosine_reg0 <= 36'sb10001010010010001010110101111001100;
            sine_reg0   <= 36'sb11010111011100000010010110100001110;
        end
        653: begin
            cosine_reg0 <= 36'sb10001001111101000000100010011111100;
            sine_reg0   <= 36'sb11010111101001100110001011010100001;
        end
        654: begin
            cosine_reg0 <= 36'sb10001001100111110100111001111111011;
            sine_reg0   <= 36'sb11010111110111000111111011000100111;
        end
        655: begin
            cosine_reg0 <= 36'sb10001001010010100111111100100110001;
            sine_reg0   <= 36'sb11011000000100100111100101101011110;
        end
        656: begin
            cosine_reg0 <= 36'sb10001000111101011001101010100000110;
            sine_reg0   <= 36'sb11011000010010000101001011000000100;
        end
        657: begin
            cosine_reg0 <= 36'sb10001000101000001010000011111100100;
            sine_reg0   <= 36'sb11011000011111100000101010111010110;
        end
        658: begin
            cosine_reg0 <= 36'sb10001000010010111001001001000110100;
            sine_reg0   <= 36'sb11011000101100111010000101010010010;
        end
        659: begin
            cosine_reg0 <= 36'sb10000111111101100110111010001011101;
            sine_reg0   <= 36'sb11011000111010010001011001111110110;
        end
        660: begin
            cosine_reg0 <= 36'sb10000111101000010011010111011001010;
            sine_reg0   <= 36'sb11011001000111100110101000110111111;
        end
        661: begin
            cosine_reg0 <= 36'sb10000111010010111110100000111100011;
            sine_reg0   <= 36'sb11011001010100111001110001110101100;
        end
        662: begin
            cosine_reg0 <= 36'sb10000110111101101000010111000010010;
            sine_reg0   <= 36'sb11011001100010001010110100101111100;
        end
        663: begin
            cosine_reg0 <= 36'sb10000110101000010000111001111000000;
            sine_reg0   <= 36'sb11011001101111011001110001011101100;
        end
        664: begin
            cosine_reg0 <= 36'sb10000110010010111000001001101010111;
            sine_reg0   <= 36'sb11011001111100100110100111110111100;
        end
        665: begin
            cosine_reg0 <= 36'sb10000101111101011110000110100111111;
            sine_reg0   <= 36'sb11011010001001110001010111110101011;
        end
        666: begin
            cosine_reg0 <= 36'sb10000101101000000010110000111100011;
            sine_reg0   <= 36'sb11011010010110111010000001001110111;
        end
        667: begin
            cosine_reg0 <= 36'sb10000101010010100110001000110101101;
            sine_reg0   <= 36'sb11011010100100000000100011111011111;
        end
        668: begin
            cosine_reg0 <= 36'sb10000100111101001000001110100000101;
            sine_reg0   <= 36'sb11011010110001000100111111110100100;
        end
        669: begin
            cosine_reg0 <= 36'sb10000100100111101001000010001010111;
            sine_reg0   <= 36'sb11011010111110000111010100110000100;
        end
        670: begin
            cosine_reg0 <= 36'sb10000100010010001000100100000001100;
            sine_reg0   <= 36'sb11011011001011000111100010100111111;
        end
        671: begin
            cosine_reg0 <= 36'sb10000011111100100110110100010001110;
            sine_reg0   <= 36'sb11011011011000000101101001010010101;
        end
        672: begin
            cosine_reg0 <= 36'sb10000011100111000011110011001001000;
            sine_reg0   <= 36'sb11011011100101000001101000101000101;
        end
        673: begin
            cosine_reg0 <= 36'sb10000011010001011111100000110100100;
            sine_reg0   <= 36'sb11011011110001111011100000100010010;
        end
        674: begin
            cosine_reg0 <= 36'sb10000010111011111001111101100001100;
            sine_reg0   <= 36'sb11011011111110110011010000110111001;
        end
        675: begin
            cosine_reg0 <= 36'sb10000010100110010011001001011101011;
            sine_reg0   <= 36'sb11011100001011101000111001011111100;
        end
        676: begin
            cosine_reg0 <= 36'sb10000010010000101011000100110101011;
            sine_reg0   <= 36'sb11011100011000011100011010010011100;
        end
        677: begin
            cosine_reg0 <= 36'sb10000001111011000001101111110110111;
            sine_reg0   <= 36'sb11011100100101001101110011001011010;
        end
        678: begin
            cosine_reg0 <= 36'sb10000001100101010111001010101111011;
            sine_reg0   <= 36'sb11011100110001111101000011111110101;
        end
        679: begin
            cosine_reg0 <= 36'sb10000001001111101011010101101100000;
            sine_reg0   <= 36'sb11011100111110101010001100100110001;
        end
        680: begin
            cosine_reg0 <= 36'sb10000000111001111110010000111010011;
            sine_reg0   <= 36'sb11011101001011010101001100111001101;
        end
        681: begin
            cosine_reg0 <= 36'sb10000000100100001111111100100111101;
            sine_reg0   <= 36'sb11011101010111111110000100110001011;
        end
        682: begin
            cosine_reg0 <= 36'sb10000000001110100000011001000001010;
            sine_reg0   <= 36'sb11011101100100100100110100000101101;
        end
        683: begin
            cosine_reg0 <= 36'sb1111111111000101111100110010100110;
            sine_reg0   <= 36'sb11011101110001001001011010101110101;
        end
        684: begin
            cosine_reg0 <= 36'sb1111111100010111101100100101111100;
            sine_reg0   <= 36'sb11011101111101101011111000100100100;
        end
        685: begin
            cosine_reg0 <= 36'sb1111111001101001010010100011111000;
            sine_reg0   <= 36'sb11011110001010001100001101011111101;
        end
        686: begin
            cosine_reg0 <= 36'sb1111110110111010101110101110000100;
            sine_reg0   <= 36'sb11011110010110101010011001011000010;
        end
        687: begin
            cosine_reg0 <= 36'sb1111110100001100000001000110001101;
            sine_reg0   <= 36'sb11011110100011000110011100000110110;
        end
        688: begin
            cosine_reg0 <= 36'sb1111110001011101001001101101111111;
            sine_reg0   <= 36'sb11011110101111100000010101100011011;
        end
        689: begin
            cosine_reg0 <= 36'sb1111101110101110001000100111000100;
            sine_reg0   <= 36'sb11011110111011111000000101100110100;
        end
        690: begin
            cosine_reg0 <= 36'sb1111101011111110111101110011001010;
            sine_reg0   <= 36'sb11011111001000001101101100001000011;
        end
        691: begin
            cosine_reg0 <= 36'sb1111101001001111101001010011111101;
            sine_reg0   <= 36'sb11011111010100100001001001000001101;
        end
        692: begin
            cosine_reg0 <= 36'sb1111100110100000001011001011000111;
            sine_reg0   <= 36'sb11011111100000110010011100001010100;
        end
        693: begin
            cosine_reg0 <= 36'sb1111100011110000100011011010010111;
            sine_reg0   <= 36'sb11011111101101000001100101011011100;
        end
        694: begin
            cosine_reg0 <= 36'sb1111100001000000110010000011011000;
            sine_reg0   <= 36'sb11011111111001001110100100101101000;
        end
        695: begin
            cosine_reg0 <= 36'sb1111011110010000110111000111110101;
            sine_reg0   <= 36'sb11100000000101011001011001110111100;
        end
        696: begin
            cosine_reg0 <= 36'sb1111011011100000110010101001011101;
            sine_reg0   <= 36'sb11100000010001100010000100110011100;
        end
        697: begin
            cosine_reg0 <= 36'sb1111011000110000100100101001111100;
            sine_reg0   <= 36'sb11100000011101101000100101011001100;
        end
        698: begin
            cosine_reg0 <= 36'sb1111010110000000001101001010111110;
            sine_reg0   <= 36'sb11100000101001101100111011100010001;
        end
        699: begin
            cosine_reg0 <= 36'sb1111010011001111101100001110010000;
            sine_reg0   <= 36'sb11100000110101101111000111000101110;
        end
        700: begin
            cosine_reg0 <= 36'sb1111010000011111000001110101011111;
            sine_reg0   <= 36'sb11100001000001101111000111111101001;
        end
        701: begin
            cosine_reg0 <= 36'sb1111001101101110001110000010010111;
            sine_reg0   <= 36'sb11100001001101101100111110000000111;
        end
        702: begin
            cosine_reg0 <= 36'sb1111001010111101010000110110100111;
            sine_reg0   <= 36'sb11100001011001101000101001001001100;
        end
        703: begin
            cosine_reg0 <= 36'sb1111001000001100001010010011111011;
            sine_reg0   <= 36'sb11100001100101100010001001001111101;
        end
        704: begin
            cosine_reg0 <= 36'sb1111000101011010111010011100000000;
            sine_reg0   <= 36'sb11100001110001011001011110001011111;
        end
        705: begin
            cosine_reg0 <= 36'sb1111000010101001100001010000100100;
            sine_reg0   <= 36'sb11100001111101001110100111110111001;
        end
        706: begin
            cosine_reg0 <= 36'sb1110111111110111111110110011010101;
            sine_reg0   <= 36'sb11100010001001000001100110001010000;
        end
        707: begin
            cosine_reg0 <= 36'sb1110111101000110010011000101111111;
            sine_reg0   <= 36'sb11100010010100110010011000111101001;
        end
        708: begin
            cosine_reg0 <= 36'sb1110111010010100011110001010010000;
            sine_reg0   <= 36'sb11100010100000100001000000001001010;
        end
        709: begin
            cosine_reg0 <= 36'sb1110110111100010100000000001110110;
            sine_reg0   <= 36'sb11100010101100001101011011100111010;
        end
        710: begin
            cosine_reg0 <= 36'sb1110110100110000011000101110011111;
            sine_reg0   <= 36'sb11100010110111110111101011001111111;
        end
        711: begin
            cosine_reg0 <= 36'sb1110110001111110001000010001111000;
            sine_reg0   <= 36'sb11100011000011011111101110111011111;
        end
        712: begin
            cosine_reg0 <= 36'sb1110101111001011101110101101110000;
            sine_reg0   <= 36'sb11100011001111000101100110100100001;
        end
        713: begin
            cosine_reg0 <= 36'sb1110101100011001001100000011110101;
            sine_reg0   <= 36'sb11100011011010101001010010000001100;
        end
        714: begin
            cosine_reg0 <= 36'sb1110101001100110100000010101110101;
            sine_reg0   <= 36'sb11100011100110001010110001001100111;
        end
        715: begin
            cosine_reg0 <= 36'sb1110100110110011101011100101011101;
            sine_reg0   <= 36'sb11100011110001101010000011111111000;
        end
        716: begin
            cosine_reg0 <= 36'sb1110100100000000101101110100011101;
            sine_reg0   <= 36'sb11100011111101000111001010010001000;
        end
        717: begin
            cosine_reg0 <= 36'sb1110100001001101100111000100100010;
            sine_reg0   <= 36'sb11100100001000100010000011111011101;
        end
        718: begin
            cosine_reg0 <= 36'sb1110011110011010010111010111011100;
            sine_reg0   <= 36'sb11100100010011111010110000111000000;
        end
        719: begin
            cosine_reg0 <= 36'sb1110011011100110111110101110111000;
            sine_reg0   <= 36'sb11100100011111010001010000111110111;
        end
        720: begin
            cosine_reg0 <= 36'sb1110011000110011011101001100100110;
            sine_reg0   <= 36'sb11100100101010100101100100001001100;
        end
        721: begin
            cosine_reg0 <= 36'sb1110010101111111110010110010010100;
            sine_reg0   <= 36'sb11100100110101110111101010010000110;
        end
        722: begin
            cosine_reg0 <= 36'sb1110010011001011111111100001110000;
            sine_reg0   <= 36'sb11100101000001000111100011001101110;
        end
        723: begin
            cosine_reg0 <= 36'sb1110010000011000000011011100101011;
            sine_reg0   <= 36'sb11100101001100010101001110111001011;
        end
        724: begin
            cosine_reg0 <= 36'sb1110001101100011111110100100110010;
            sine_reg0   <= 36'sb11100101010111100000101101001100111;
        end
        725: begin
            cosine_reg0 <= 36'sb1110001010101111110000111011110110;
            sine_reg0   <= 36'sb11100101100010101001111110000001011;
        end
        726: begin
            cosine_reg0 <= 36'sb1110000111111011011010100011100100;
            sine_reg0   <= 36'sb11100101101101110001000001001111111;
        end
        727: begin
            cosine_reg0 <= 36'sb1110000101000110111011011101101101;
            sine_reg0   <= 36'sb11100101111000110101110110110001101;
        end
        728: begin
            cosine_reg0 <= 36'sb1110000010010010010011101100000000;
            sine_reg0   <= 36'sb11100110000011111000011110011111110;
        end
        729: begin
            cosine_reg0 <= 36'sb1101111111011101100011010000001011;
            sine_reg0   <= 36'sb11100110001110111000111000010011100;
        end
        730: begin
            cosine_reg0 <= 36'sb1101111100101000101010001100000000;
            sine_reg0   <= 36'sb11100110011001110111000100000110000;
        end
        731: begin
            cosine_reg0 <= 36'sb1101111001110011101000100001001100;
            sine_reg0   <= 36'sb11100110100100110011000001110000100;
        end
        732: begin
            cosine_reg0 <= 36'sb1101110110111110011110010001100000;
            sine_reg0   <= 36'sb11100110101111101100110001001100010;
        end
        733: begin
            cosine_reg0 <= 36'sb1101110100001001001011011110101100;
            sine_reg0   <= 36'sb11100110111010100100010010010010100;
        end
        734: begin
            cosine_reg0 <= 36'sb1101110001010011110000001010011111;
            sine_reg0   <= 36'sb11100111000101011001100100111100110;
        end
        735: begin
            cosine_reg0 <= 36'sb1101101110011110001100010110101010;
            sine_reg0   <= 36'sb11100111010000001100101001000100000;
        end
        736: begin
            cosine_reg0 <= 36'sb1101101011101000100000000100111100;
            sine_reg0   <= 36'sb11100111011010111101011110100001110;
        end
        737: begin
            cosine_reg0 <= 36'sb1101101000110010101011010111000101;
            sine_reg0   <= 36'sb11100111100101101100000101001111100;
        end
        738: begin
            cosine_reg0 <= 36'sb1101100101111100101110001110110110;
            sine_reg0   <= 36'sb11100111110000011000011101000110011;
        end
        739: begin
            cosine_reg0 <= 36'sb1101100011000110101000101101111111;
            sine_reg0   <= 36'sb11100111111011000010100101111111111;
        end
        740: begin
            cosine_reg0 <= 36'sb1101100000010000011010110110001111;
            sine_reg0   <= 36'sb11101000000101101010011111110101100;
        end
        741: begin
            cosine_reg0 <= 36'sb1101011101011010000100101001011001;
            sine_reg0   <= 36'sb11101000010000010000001010100000101;
        end
        742: begin
            cosine_reg0 <= 36'sb1101011010100011100110001001001011;
            sine_reg0   <= 36'sb11101000011010110011100101111010110;
        end
        743: begin
            cosine_reg0 <= 36'sb1101010111101100111111010111010111;
            sine_reg0   <= 36'sb11101000100101010100110001111101010;
        end
        744: begin
            cosine_reg0 <= 36'sb1101010100110110010000010101101101;
            sine_reg0   <= 36'sb11101000101111110011101110100001111;
        end
        745: begin
            cosine_reg0 <= 36'sb1101010001111111011001000101111110;
            sine_reg0   <= 36'sb11101000111010010000011011100001111;
        end
        746: begin
            cosine_reg0 <= 36'sb1101001111001000011001101001111011;
            sine_reg0   <= 36'sb11101001000100101010111000110111001;
        end
        747: begin
            cosine_reg0 <= 36'sb1101001100010001010010000011010100;
            sine_reg0   <= 36'sb11101001001111000011000110011010111;
        end
        748: begin
            cosine_reg0 <= 36'sb1101001001011010000010010011111011;
            sine_reg0   <= 36'sb11101001011001011001000100000110111;
        end
        749: begin
            cosine_reg0 <= 36'sb1101000110100010101010011101100001;
            sine_reg0   <= 36'sb11101001100011101100110001110100111;
        end
        750: begin
            cosine_reg0 <= 36'sb1101000011101011001010100001110110;
            sine_reg0   <= 36'sb11101001101101111110001111011110010;
        end
        751: begin
            cosine_reg0 <= 36'sb1101000000110011100010100010101100;
            sine_reg0   <= 36'sb11101001111000001101011100111100111;
        end
        752: begin
            cosine_reg0 <= 36'sb1100111101111011110010100001110101;
            sine_reg0   <= 36'sb11101010000010011010011010001010011;
        end
        753: begin
            cosine_reg0 <= 36'sb1100111011000011111010100001000001;
            sine_reg0   <= 36'sb11101010001100100101000111000000011;
        end
        754: begin
            cosine_reg0 <= 36'sb1100111000001011111010100010000001;
            sine_reg0   <= 36'sb11101010010110101101100011011000101;
        end
        755: begin
            cosine_reg0 <= 36'sb1100110101010011110010100110101001;
            sine_reg0   <= 36'sb11101010100000110011101111001101000;
        end
        756: begin
            cosine_reg0 <= 36'sb1100110010011011100010110000101000;
            sine_reg0   <= 36'sb11101010101010110111101010010111001;
        end
        757: begin
            cosine_reg0 <= 36'sb1100101111100011001011000001110001;
            sine_reg0   <= 36'sb11101010110100111001010100110001000;
        end
        758: begin
            cosine_reg0 <= 36'sb1100101100101010101011011011110101;
            sine_reg0   <= 36'sb11101010111110111000101110010100001;
        end
        759: begin
            cosine_reg0 <= 36'sb1100101001110010000100000000100111;
            sine_reg0   <= 36'sb11101011001000110101110110111010101;
        end
        760: begin
            cosine_reg0 <= 36'sb1100100110111001010100110001110111;
            sine_reg0   <= 36'sb11101011010010110000101110011110010;
        end
        761: begin
            cosine_reg0 <= 36'sb1100100100000000011101110001011001;
            sine_reg0   <= 36'sb11101011011100101001010100111000110;
        end
        762: begin
            cosine_reg0 <= 36'sb1100100001000111011111000000111110;
            sine_reg0   <= 36'sb11101011100110011111101010000100010;
        end
        763: begin
            cosine_reg0 <= 36'sb1100011110001110011000100010010111;
            sine_reg0   <= 36'sb11101011110000010011101101111010101;
        end
        764: begin
            cosine_reg0 <= 36'sb1100011011010101001010010111011001;
            sine_reg0   <= 36'sb11101011111010000101100000010101101;
        end
        765: begin
            cosine_reg0 <= 36'sb1100011000011011110100100001110100;
            sine_reg0   <= 36'sb11101100000011110101000001001111100;
        end
        766: begin
            cosine_reg0 <= 36'sb1100010101100010010111000011011010;
            sine_reg0   <= 36'sb11101100001101100010010000100010000;
        end
        767: begin
            cosine_reg0 <= 36'sb1100010010101000110001111101111111;
            sine_reg0   <= 36'sb11101100010111001101001110000111011;
        end
        768: begin
            cosine_reg0 <= 36'sb1100001111101111000101010011010101;
            sine_reg0   <= 36'sb11101100100000110101111001111001100;
        end
        769: begin
            cosine_reg0 <= 36'sb1100001100110101010001000101001111;
            sine_reg0   <= 36'sb11101100101010011100010011110010011;
        end
        770: begin
            cosine_reg0 <= 36'sb1100001001111011010101010101011110;
            sine_reg0   <= 36'sb11101100110100000000011011101100010;
        end
        771: begin
            cosine_reg0 <= 36'sb1100000111000001010010000101110110;
            sine_reg0   <= 36'sb11101100111101100010010001100001001;
        end
        772: begin
            cosine_reg0 <= 36'sb1100000100000111000111011000001001;
            sine_reg0   <= 36'sb11101101000111000001110101001011001;
        end
        773: begin
            cosine_reg0 <= 36'sb1100000001001100110101001110001011;
            sine_reg0   <= 36'sb11101101010000011111000110100100011;
        end
        774: begin
            cosine_reg0 <= 36'sb1011111110010010011011101001101110;
            sine_reg0   <= 36'sb11101101011001111010000101100111001;
        end
        775: begin
            cosine_reg0 <= 36'sb1011111011010111111010101100100101;
            sine_reg0   <= 36'sb11101101100011010010110010001101100;
        end
        776: begin
            cosine_reg0 <= 36'sb1011111000011101010010011000100011;
            sine_reg0   <= 36'sb11101101101100101001001100010001101;
        end
        777: begin
            cosine_reg0 <= 36'sb1011110101100010100010101111011100;
            sine_reg0   <= 36'sb11101101110101111101010011101110000;
        end
        778: begin
            cosine_reg0 <= 36'sb1011110010100111101011110011000010;
            sine_reg0   <= 36'sb11101101111111001111001000011100100;
        end
        779: begin
            cosine_reg0 <= 36'sb1011101111101100101101100101001001;
            sine_reg0   <= 36'sb11101110001000011110101010010111110;
        end
        780: begin
            cosine_reg0 <= 36'sb1011101100110001101000000111100100;
            sine_reg0   <= 36'sb11101110010001101011111001011001111;
        end
        781: begin
            cosine_reg0 <= 36'sb1011101001110110011011011100000111;
            sine_reg0   <= 36'sb11101110011010110110110101011101010;
        end
        782: begin
            cosine_reg0 <= 36'sb1011100110111011000111100100100100;
            sine_reg0   <= 36'sb11101110100011111111011110011100010;
        end
        783: begin
            cosine_reg0 <= 36'sb1011100011111111101100100010110001;
            sine_reg0   <= 36'sb11101110101101000101110100010001001;
        end
        784: begin
            cosine_reg0 <= 36'sb1011100001000100001010011000011111;
            sine_reg0   <= 36'sb11101110110110001001110110110110010;
        end
        785: begin
            cosine_reg0 <= 36'sb1011011110001000100001000111100011;
            sine_reg0   <= 36'sb11101110111111001011100110000110010;
        end
        786: begin
            cosine_reg0 <= 36'sb1011011011001100110000110001110001;
            sine_reg0   <= 36'sb11101111001000001011000001111011010;
        end
        787: begin
            cosine_reg0 <= 36'sb1011011000010000111001011000111100;
            sine_reg0   <= 36'sb11101111010001001000001010010000000;
        end
        788: begin
            cosine_reg0 <= 36'sb1011010101010100111010111110111001;
            sine_reg0   <= 36'sb11101111011010000010111110111110111;
        end
        789: begin
            cosine_reg0 <= 36'sb1011010010011000110101100101011010;
            sine_reg0   <= 36'sb11101111100010111011100000000010010;
        end
        790: begin
            cosine_reg0 <= 36'sb1011001111011100101001001110010101;
            sine_reg0   <= 36'sb11101111101011110001101101010100110;
        end
        791: begin
            cosine_reg0 <= 36'sb1011001100100000010101111011011110;
            sine_reg0   <= 36'sb11101111110100100101100110110000111;
        end
        792: begin
            cosine_reg0 <= 36'sb1011001001100011111011101110101000;
            sine_reg0   <= 36'sb11101111111101010111001100010001010;
        end
        793: begin
            cosine_reg0 <= 36'sb1011000110100111011010101001100111;
            sine_reg0   <= 36'sb11110000000110000110011101110000100;
        end
        794: begin
            cosine_reg0 <= 36'sb1011000011101010110010101110010001;
            sine_reg0   <= 36'sb11110000001110110011011011001001001;
        end
        795: begin
            cosine_reg0 <= 36'sb1011000000101110000011111110011001;
            sine_reg0   <= 36'sb11110000010111011110000100010101110;
        end
        796: begin
            cosine_reg0 <= 36'sb1010111101110001001110011011110011;
            sine_reg0   <= 36'sb11110000100000000110011001010001001;
        end
        797: begin
            cosine_reg0 <= 36'sb1010111010110100010010001000010110;
            sine_reg0   <= 36'sb11110000101000101100011001110101111;
        end
        798: begin
            cosine_reg0 <= 36'sb1010110111110111001111000101110011;
            sine_reg0   <= 36'sb11110000110001010000000101111110110;
        end
        799: begin
            cosine_reg0 <= 36'sb1010110100111010000101010110000010;
            sine_reg0   <= 36'sb11110000111001110001011101100110011;
        end
        800: begin
            cosine_reg0 <= 36'sb1010110001111100110100111010110101;
            sine_reg0   <= 36'sb11110001000010010000100000100111101;
        end
        801: begin
            cosine_reg0 <= 36'sb1010101110111111011101110110000010;
            sine_reg0   <= 36'sb11110001001010101101001110111101001;
        end
        802: begin
            cosine_reg0 <= 36'sb1010101100000010000000001001011110;
            sine_reg0   <= 36'sb11110001010011000111101000100001101;
        end
        803: begin
            cosine_reg0 <= 36'sb1010101001000100011011110110111110;
            sine_reg0   <= 36'sb11110001011011011111101101010000001;
        end
        804: begin
            cosine_reg0 <= 36'sb1010100110000110110001000000010110;
            sine_reg0   <= 36'sb11110001100011110101011101000011011;
        end
        805: begin
            cosine_reg0 <= 36'sb1010100011001000111111100111011011;
            sine_reg0   <= 36'sb11110001101100001000110111110110010;
        end
        806: begin
            cosine_reg0 <= 36'sb1010100000001011000111101110000011;
            sine_reg0   <= 36'sb11110001110100011001111101100011101;
        end
        807: begin
            cosine_reg0 <= 36'sb1010011101001101001001010110000010;
            sine_reg0   <= 36'sb11110001111100101000101110000110010;
        end
        808: begin
            cosine_reg0 <= 36'sb1010011010001111000100100001001111;
            sine_reg0   <= 36'sb11110010000100110101001001011001010;
        end
        809: begin
            cosine_reg0 <= 36'sb1010010111010000111001010001011101;
            sine_reg0   <= 36'sb11110010001100111111001111010111100;
        end
        810: begin
            cosine_reg0 <= 36'sb1010010100010010100111101000100011;
            sine_reg0   <= 36'sb11110010010101000110111111111100000;
        end
        811: begin
            cosine_reg0 <= 36'sb1010010001010100001111101000010110;
            sine_reg0   <= 36'sb11110010011101001100011011000001101;
        end
        812: begin
            cosine_reg0 <= 36'sb1010001110010101110001010010101011;
            sine_reg0   <= 36'sb11110010100101001111100000100011100;
        end
        813: begin
            cosine_reg0 <= 36'sb1010001011010111001100101001010111;
            sine_reg0   <= 36'sb11110010101101010000010000011100101;
        end
        814: begin
            cosine_reg0 <= 36'sb1010001000011000100001101110010001;
            sine_reg0   <= 36'sb11110010110101001110101010101000000;
        end
        815: begin
            cosine_reg0 <= 36'sb1010000101011001110000100011001101;
            sine_reg0   <= 36'sb11110010111101001010101111000000111;
        end
        816: begin
            cosine_reg0 <= 36'sb1010000010011010111001001010000011;
            sine_reg0   <= 36'sb11110011000101000100011101100010001;
        end
        817: begin
            cosine_reg0 <= 36'sb1001111111011011111011100100100110;
            sine_reg0   <= 36'sb11110011001100111011110110000111001;
        end
        818: begin
            cosine_reg0 <= 36'sb1001111100011100110111110100101110;
            sine_reg0   <= 36'sb11110011010100110000111000101010110;
        end
        819: begin
            cosine_reg0 <= 36'sb1001111001011101101101111100001111;
            sine_reg0   <= 36'sb11110011011100100011100101001000100;
        end
        820: begin
            cosine_reg0 <= 36'sb1001110110011110011101111101000000;
            sine_reg0   <= 36'sb11110011100100010011111011011011010;
        end
        821: begin
            cosine_reg0 <= 36'sb1001110011011111000111111000110111;
            sine_reg0   <= 36'sb11110011101100000001111011011110011;
        end
        822: begin
            cosine_reg0 <= 36'sb1001110000011111101011110001101010;
            sine_reg0   <= 36'sb11110011110011101101100101001101000;
        end
        823: begin
            cosine_reg0 <= 36'sb1001101101100000001001101001001111;
            sine_reg0   <= 36'sb11110011111011010110111000100010101;
        end
        824: begin
            cosine_reg0 <= 36'sb1001101010100000100001100001011100;
            sine_reg0   <= 36'sb11110100000010111101110101011010010;
        end
        825: begin
            cosine_reg0 <= 36'sb1001100111100000110011011100000111;
            sine_reg0   <= 36'sb11110100001010100010011011101111011;
        end
        826: begin
            cosine_reg0 <= 36'sb1001100100100000111111011011000111;
            sine_reg0   <= 36'sb11110100010010000100101011011101010;
        end
        827: begin
            cosine_reg0 <= 36'sb1001100001100001000101100000010001;
            sine_reg0   <= 36'sb11110100011001100100100100011111010;
        end
        828: begin
            cosine_reg0 <= 36'sb1001011110100001000101101101011101;
            sine_reg0   <= 36'sb11110100100001000010000110110000111;
        end
        829: begin
            cosine_reg0 <= 36'sb1001011011100001000000000100100001;
            sine_reg0   <= 36'sb11110100101000011101010010001101010;
        end
        830: begin
            cosine_reg0 <= 36'sb1001011000100000110100100111010010;
            sine_reg0   <= 36'sb11110100101111110110000110101111111;
        end
        831: begin
            cosine_reg0 <= 36'sb1001010101100000100011010111101001;
            sine_reg0   <= 36'sb11110100110111001100100100010100011;
        end
        832: begin
            cosine_reg0 <= 36'sb1001010010100000001100010111011010;
            sine_reg0   <= 36'sb11110100111110100000101010110110001;
        end
        833: begin
            cosine_reg0 <= 36'sb1001001111011111101111101000011110;
            sine_reg0   <= 36'sb11110101000101110010011010010000100;
        end
        834: begin
            cosine_reg0 <= 36'sb1001001100011111001101001100101010;
            sine_reg0   <= 36'sb11110101001101000001110010011111001;
        end
        835: begin
            cosine_reg0 <= 36'sb1001001001011110100101000101110110;
            sine_reg0   <= 36'sb11110101010100001110110011011101100;
        end
        836: begin
            cosine_reg0 <= 36'sb1001000110011101110111010101111000;
            sine_reg0   <= 36'sb11110101011011011001011101000111001;
        end
        837: begin
            cosine_reg0 <= 36'sb1001000011011101000011111110100111;
            sine_reg0   <= 36'sb11110101100010100001101111010111101;
        end
        838: begin
            cosine_reg0 <= 36'sb1001000000011100001011000001111011;
            sine_reg0   <= 36'sb11110101101001100111101010001010110;
        end
        839: begin
            cosine_reg0 <= 36'sb1000111101011011001100100001101001;
            sine_reg0   <= 36'sb11110101110000101011001101011011111;
        end
        840: begin
            cosine_reg0 <= 36'sb1000111010011010001000011111101001;
            sine_reg0   <= 36'sb11110101110111101100011001000110111;
        end
        841: begin
            cosine_reg0 <= 36'sb1000110111011000111110111101110011;
            sine_reg0   <= 36'sb11110101111110101011001101000111010;
        end
        842: begin
            cosine_reg0 <= 36'sb1000110100010111101111111101111101;
            sine_reg0   <= 36'sb11110110000101100111101001011000110;
        end
        843: begin
            cosine_reg0 <= 36'sb1000110001010110011011100001111110;
            sine_reg0   <= 36'sb11110110001100100001101101110111001;
        end
        844: begin
            cosine_reg0 <= 36'sb1000101110010101000001101011101111;
            sine_reg0   <= 36'sb11110110010011011001011010011110000;
        end
        845: begin
            cosine_reg0 <= 36'sb1000101011010011100010011101000101;
            sine_reg0   <= 36'sb11110110011010001110101111001001010;
        end
        846: begin
            cosine_reg0 <= 36'sb1000101000010001111101110111111001;
            sine_reg0   <= 36'sb11110110100001000001101011110100101;
        end
        847: begin
            cosine_reg0 <= 36'sb1000100101010000010011111110000001;
            sine_reg0   <= 36'sb11110110100111110010010000011100000;
        end
        848: begin
            cosine_reg0 <= 36'sb1000100010001110100100110001010110;
            sine_reg0   <= 36'sb11110110101110100000011100111011001;
        end
        849: begin
            cosine_reg0 <= 36'sb1000011111001100110000010011101111;
            sine_reg0   <= 36'sb11110110110101001100010001001101111;
        end
        850: begin
            cosine_reg0 <= 36'sb1000011100001010110110100111000011;
            sine_reg0   <= 36'sb11110110111011110101101101010000001;
        end
        851: begin
            cosine_reg0 <= 36'sb1000011001001000110111101101001010;
            sine_reg0   <= 36'sb11110111000010011100110000111101110;
        end
        852: begin
            cosine_reg0 <= 36'sb1000010110000110110011100111111011;
            sine_reg0   <= 36'sb11110111001001000001011100010010110;
        end
        853: begin
            cosine_reg0 <= 36'sb1000010011000100101010011001001111;
            sine_reg0   <= 36'sb11110111001111100011101111001010111;
        end
        854: begin
            cosine_reg0 <= 36'sb1000010000000010011100000010111101;
            sine_reg0   <= 36'sb11110111010110000011101001100010011;
        end
        855: begin
            cosine_reg0 <= 36'sb1000001101000000001000100110111101;
            sine_reg0   <= 36'sb11110111011100100001001011010101001;
        end
        856: begin
            cosine_reg0 <= 36'sb1000001001111101110000000111000111;
            sine_reg0   <= 36'sb11110111100010111100010100011111000;
        end
        857: begin
            cosine_reg0 <= 36'sb1000000110111011010010100101010010;
            sine_reg0   <= 36'sb11110111101001010101000100111100010;
        end
        858: begin
            cosine_reg0 <= 36'sb1000000011111000110000000011010111;
            sine_reg0   <= 36'sb11110111101111101011011100101000110;
        end
        859: begin
            cosine_reg0 <= 36'sb1000000000110110001000100011001110;
            sine_reg0   <= 36'sb11110111110101111111011011100000110;
        end
        860: begin
            cosine_reg0 <= 36'sb111111101110011011100000110101110;
            sine_reg0   <= 36'sb11110111111100010001000001100000010;
        end
        861: begin
            cosine_reg0 <= 36'sb111111010110000101010101111110000;
            sine_reg0   <= 36'sb11111000000010100000001110100011011;
        end
        862: begin
            cosine_reg0 <= 36'sb111110111101101110100100000001100;
            sine_reg0   <= 36'sb11111000001000101101000010100110011;
        end
        863: begin
            cosine_reg0 <= 36'sb111110100101010111001011001111010;
            sine_reg0   <= 36'sb11111000001110110111011101100101011;
        end
        864: begin
            cosine_reg0 <= 36'sb111110001100111111001011110110010;
            sine_reg0   <= 36'sb11111000010100111111011111011100100;
        end
        865: begin
            cosine_reg0 <= 36'sb111101110100100110100110000101101;
            sine_reg0   <= 36'sb11111000011011000101001000001000000;
        end
        866: begin
            cosine_reg0 <= 36'sb111101011100001101011010001100011;
            sine_reg0   <= 36'sb11111000100001001000010111100100001;
        end
        867: begin
            cosine_reg0 <= 36'sb111101000011110011101000011001100;
            sine_reg0   <= 36'sb11111000100111001001001101101101010;
        end
        868: begin
            cosine_reg0 <= 36'sb111100101011011001010000111100001;
            sine_reg0   <= 36'sb11111000101101000111101010011111101;
        end
        869: begin
            cosine_reg0 <= 36'sb111100010010111110010100000011010;
            sine_reg0   <= 36'sb11111000110011000011101101110111100;
        end
        870: begin
            cosine_reg0 <= 36'sb111011111010100010110001111110000;
            sine_reg0   <= 36'sb11111000111000111101010111110001001;
        end
        871: begin
            cosine_reg0 <= 36'sb111011100010000110101010111011011;
            sine_reg0   <= 36'sb11111000111110110100101000001001000;
        end
        872: begin
            cosine_reg0 <= 36'sb111011001001101001111111001010100;
            sine_reg0   <= 36'sb11111001000100101001011110111011101;
        end
        873: begin
            cosine_reg0 <= 36'sb111010110001001100101110111010100;
            sine_reg0   <= 36'sb11111001001010011011111100000101001;
        end
        874: begin
            cosine_reg0 <= 36'sb111010011000101110111010011010011;
            sine_reg0   <= 36'sb11111001010000001011111111100010001;
        end
        875: begin
            cosine_reg0 <= 36'sb111010000000010000100001111001001;
            sine_reg0   <= 36'sb11111001010101111001101001001110111;
        end
        876: begin
            cosine_reg0 <= 36'sb111001100111110001100101100110001;
            sine_reg0   <= 36'sb11111001011011100100111001001000001;
        end
        877: begin
            cosine_reg0 <= 36'sb111001001111010010000101110000010;
            sine_reg0   <= 36'sb11111001100001001101101111001010010;
        end
        878: begin
            cosine_reg0 <= 36'sb111000110110110010000010100110110;
            sine_reg0   <= 36'sb11111001100110110100001011010001110;
        end
        879: begin
            cosine_reg0 <= 36'sb111000011110010001011100011000101;
            sine_reg0   <= 36'sb11111001101100011000001101011011001;
        end
        880: begin
            cosine_reg0 <= 36'sb111000000101110000010011010101000;
            sine_reg0   <= 36'sb11111001110001111001110101100011000;
        end
        881: begin
            cosine_reg0 <= 36'sb110111101101001110100111101011000;
            sine_reg0   <= 36'sb11111001110111011001000011100110000;
        end
        882: begin
            cosine_reg0 <= 36'sb110111010100101100011001101001111;
            sine_reg0   <= 36'sb11111001111100110101110111100000110;
        end
        883: begin
            cosine_reg0 <= 36'sb110110111100001001101001100000101;
            sine_reg0   <= 36'sb11111010000010010000010001001111110;
        end
        884: begin
            cosine_reg0 <= 36'sb110110100011100110010111011110100;
            sine_reg0   <= 36'sb11111010000111101000010000101111111;
        end
        885: begin
            cosine_reg0 <= 36'sb110110001011000010100011110010100;
            sine_reg0   <= 36'sb11111010001100111101110101111101101;
        end
        886: begin
            cosine_reg0 <= 36'sb110101110010011110001110101011111;
            sine_reg0   <= 36'sb11111010010010010001000000110101110;
        end
        887: begin
            cosine_reg0 <= 36'sb110101011001111001011000011001110;
            sine_reg0   <= 36'sb11111010010111100001110001010101000;
        end
        888: begin
            cosine_reg0 <= 36'sb110101000001010100000001001011011;
            sine_reg0   <= 36'sb11111010011100110000000111011000010;
        end
        889: begin
            cosine_reg0 <= 36'sb110100101000101110001001001111110;
            sine_reg0   <= 36'sb11111010100001111100000010111100000;
        end
        890: begin
            cosine_reg0 <= 36'sb110100010000000111110000110110001;
            sine_reg0   <= 36'sb11111010100111000101100011111101011;
        end
        891: begin
            cosine_reg0 <= 36'sb110011110111100000111000001101110;
            sine_reg0   <= 36'sb11111010101100001100101010011000111;
        end
        892: begin
            cosine_reg0 <= 36'sb110011011110111001011111100101110;
            sine_reg0   <= 36'sb11111010110001010001010110001011101;
        end
        893: begin
            cosine_reg0 <= 36'sb110011000110010001100111001101001;
            sine_reg0   <= 36'sb11111010110110010011100111010010011;
        end
        894: begin
            cosine_reg0 <= 36'sb110010101101101001001111010011011;
            sine_reg0   <= 36'sb11111010111011010011011101101010000;
        end
        895: begin
            cosine_reg0 <= 36'sb110010010101000000011000000111100;
            sine_reg0   <= 36'sb11111011000000010000111001001111011;
        end
        896: begin
            cosine_reg0 <= 36'sb110001111100010111000001111000110;
            sine_reg0   <= 36'sb11111011000101001011111001111111101;
        end
        897: begin
            cosine_reg0 <= 36'sb110001100011101101001100110110011;
            sine_reg0   <= 36'sb11111011001010000100011111110111100;
        end
        898: begin
            cosine_reg0 <= 36'sb110001001011000010111001001111100;
            sine_reg0   <= 36'sb11111011001110111010101010110100001;
        end
        899: begin
            cosine_reg0 <= 36'sb110000110010011000000111010011011;
            sine_reg0   <= 36'sb11111011010011101110011010110010100;
        end
        900: begin
            cosine_reg0 <= 36'sb110000011001101100110111010001010;
            sine_reg0   <= 36'sb11111011011000011111101111101111100;
        end
        901: begin
            cosine_reg0 <= 36'sb110000000001000001001001011000010;
            sine_reg0   <= 36'sb11111011011101001110101001101000100;
        end
        902: begin
            cosine_reg0 <= 36'sb101111101000010100111101110111101;
            sine_reg0   <= 36'sb11111011100001111011001000011010010;
        end
        903: begin
            cosine_reg0 <= 36'sb101111001111101000010100111110101;
            sine_reg0   <= 36'sb11111011100110100101001100000010000;
        end
        904: begin
            cosine_reg0 <= 36'sb101110110110111011001110111100101;
            sine_reg0   <= 36'sb11111011101011001100110100011100111;
        end
        905: begin
            cosine_reg0 <= 36'sb101110011110001101101100000000101;
            sine_reg0   <= 36'sb11111011101111110010000001101000001;
        end
        906: begin
            cosine_reg0 <= 36'sb101110000101011111101100011010000;
            sine_reg0   <= 36'sb11111011110100010100110011100000110;
        end
        907: begin
            cosine_reg0 <= 36'sb101101101100110001010000011000000;
            sine_reg0   <= 36'sb11111011111000110101001010000100000;
        end
        908: begin
            cosine_reg0 <= 36'sb101101010100000010011000001001111;
            sine_reg0   <= 36'sb11111011111101010011000101001111001;
        end
        909: begin
            cosine_reg0 <= 36'sb101100111011010011000011111110111;
            sine_reg0   <= 36'sb11111100000001101110100100111111010;
        end
        910: begin
            cosine_reg0 <= 36'sb101100100010100011010100000110010;
            sine_reg0   <= 36'sb11111100000110000111101001010001111;
        end
        911: begin
            cosine_reg0 <= 36'sb101100001001110011001000101111001;
            sine_reg0   <= 36'sb11111100001010011110010010000100001;
        end
        912: begin
            cosine_reg0 <= 36'sb101011110001000010100010001001001;
            sine_reg0   <= 36'sb11111100001110110010011111010011011;
        end
        913: begin
            cosine_reg0 <= 36'sb101011011000010001100000100011001;
            sine_reg0   <= 36'sb11111100010011000100010000111101000;
        end
        914: begin
            cosine_reg0 <= 36'sb101010111111100000000100001100101;
            sine_reg0   <= 36'sb11111100010111010011100110111110010;
        end
        915: begin
            cosine_reg0 <= 36'sb101010100110101110001101010100111;
            sine_reg0   <= 36'sb11111100011011100000100001010100100;
        end
        916: begin
            cosine_reg0 <= 36'sb101010001101111011111100001011001;
            sine_reg0   <= 36'sb11111100011111101010111111111101011;
        end
        917: begin
            cosine_reg0 <= 36'sb101001110101001001010000111110110;
            sine_reg0   <= 36'sb11111100100011110011000010110110000;
        end
        918: begin
            cosine_reg0 <= 36'sb101001011100010110001011111110111;
            sine_reg0   <= 36'sb11111100100111111000101001111100000;
        end
        919: begin
            cosine_reg0 <= 36'sb101001000011100010101101011011000;
            sine_reg0   <= 36'sb11111100101011111011110101001100111;
        end
        920: begin
            cosine_reg0 <= 36'sb101000101010101110110101100010010;
            sine_reg0   <= 36'sb11111100101111111100100100100110001;
        end
        921: begin
            cosine_reg0 <= 36'sb101000010001111010100100100100001;
            sine_reg0   <= 36'sb11111100110011111010111000000101010;
        end
        922: begin
            cosine_reg0 <= 36'sb100111111001000101111010101111110;
            sine_reg0   <= 36'sb11111100110111110110101111100111110;
        end
        923: begin
            cosine_reg0 <= 36'sb100111100000010000111000010100011;
            sine_reg0   <= 36'sb11111100111011110000001011001011010;
        end
        924: begin
            cosine_reg0 <= 36'sb100111000111011011011101100001101;
            sine_reg0   <= 36'sb11111100111111100111001010101101010;
        end
        925: begin
            cosine_reg0 <= 36'sb100110101110100101101010100110100;
            sine_reg0   <= 36'sb11111101000011011011101110001011101;
        end
        926: begin
            cosine_reg0 <= 36'sb100110010101101111011111110010100;
            sine_reg0   <= 36'sb11111101000111001101110101100011110;
        end
        927: begin
            cosine_reg0 <= 36'sb100101111100111000111101010101000;
            sine_reg0   <= 36'sb11111101001010111101100000110011011;
        end
        928: begin
            cosine_reg0 <= 36'sb100101100100000010000011011101001;
            sine_reg0   <= 36'sb11111101001110101010101111111000001;
        end
        929: begin
            cosine_reg0 <= 36'sb100101001011001010110010011010011;
            sine_reg0   <= 36'sb11111101010010010101100010101111111;
        end
        930: begin
            cosine_reg0 <= 36'sb100100110010010011001010011100000;
            sine_reg0   <= 36'sb11111101010101111101111001011000010;
        end
        931: begin
            cosine_reg0 <= 36'sb100100011001011011001011110001011;
            sine_reg0   <= 36'sb11111101011001100011110011101111001;
        end
        932: begin
            cosine_reg0 <= 36'sb100100000000100010110110101001111;
            sine_reg0   <= 36'sb11111101011101000111010001110010001;
        end
        933: begin
            cosine_reg0 <= 36'sb100011100111101010001011010100110;
            sine_reg0   <= 36'sb11111101100000101000010011011111001;
        end
        934: begin
            cosine_reg0 <= 36'sb100011001110110001001010000001100;
            sine_reg0   <= 36'sb11111101100100000110111000110011111;
        end
        935: begin
            cosine_reg0 <= 36'sb100010110101110111110010111111011;
            sine_reg0   <= 36'sb11111101100111100011000001101110100;
        end
        936: begin
            cosine_reg0 <= 36'sb100010011100111110000110011101110;
            sine_reg0   <= 36'sb11111101101010111100101110001100100;
        end
        937: begin
            cosine_reg0 <= 36'sb100010000100000100000100101011111;
            sine_reg0   <= 36'sb11111101101110010011111110001100001;
        end
        938: begin
            cosine_reg0 <= 36'sb100001101011001001101101111001011;
            sine_reg0   <= 36'sb11111101110001101000110001101011001;
        end
        939: begin
            cosine_reg0 <= 36'sb100001010010001111000010010101011;
            sine_reg0   <= 36'sb11111101110100111011001000100111011;
        end
        940: begin
            cosine_reg0 <= 36'sb100000111001010100000010001111100;
            sine_reg0   <= 36'sb11111101111000001011000010111111000;
        end
        941: begin
            cosine_reg0 <= 36'sb100000100000011000101101110110110;
            sine_reg0   <= 36'sb11111101111011011000100000110000000;
        end
        942: begin
            cosine_reg0 <= 36'sb100000000111011101000101011010111;
            sine_reg0   <= 36'sb11111101111110100011100001111000010;
        end
        943: begin
            cosine_reg0 <= 36'sb11111101110100001001001001011000;
            sine_reg0   <= 36'sb11111110000001101100000110010101111;
        end
        944: begin
            cosine_reg0 <= 36'sb11111010101100100111001010110101;
            sine_reg0   <= 36'sb11111110000100110010001110000110111;
        end
        945: begin
            cosine_reg0 <= 36'sb11110111100101000010110001101001;
            sine_reg0   <= 36'sb11111110000111110101111001001001100;
        end
        946: begin
            cosine_reg0 <= 36'sb11110100011101011011111111101111;
            sine_reg0   <= 36'sb11111110001010110111000111011011110;
        end
        947: begin
            cosine_reg0 <= 36'sb11110001010101110010110111000010;
            sine_reg0   <= 36'sb11111110001101110101111000111011111;
        end
        948: begin
            cosine_reg0 <= 36'sb11101110001110000111011001011101;
            sine_reg0   <= 36'sb11111110010000110010001101100111111;
        end
        949: begin
            cosine_reg0 <= 36'sb11101011000110011001101000111100;
            sine_reg0   <= 36'sb11111110010011101100000101011110000;
        end
        950: begin
            cosine_reg0 <= 36'sb11100111111110101001100111011001;
            sine_reg0   <= 36'sb11111110010110100011100000011100011;
        end
        951: begin
            cosine_reg0 <= 36'sb11100100110110110111010110110001;
            sine_reg0   <= 36'sb11111110011001011000011110100001100;
        end
        952: begin
            cosine_reg0 <= 36'sb11100001101111000010111000111101;
            sine_reg0   <= 36'sb11111110011100001010111111101011010;
        end
        953: begin
            cosine_reg0 <= 36'sb11011110100111001100001111111001;
            sine_reg0   <= 36'sb11111110011110111011000011111000010;
        end
        954: begin
            cosine_reg0 <= 36'sb11011011011111010011011101100010;
            sine_reg0   <= 36'sb11111110100001101000101011000110101;
        end
        955: begin
            cosine_reg0 <= 36'sb11011000010111011000100011110001;
            sine_reg0   <= 36'sb11111110100100010011110101010100110;
        end
        956: begin
            cosine_reg0 <= 36'sb11010101001111011011100100100010;
            sine_reg0   <= 36'sb11111110100110111100100010100001000;
        end
        957: begin
            cosine_reg0 <= 36'sb11010010000111011100100001110001;
            sine_reg0   <= 36'sb11111110101001100010110010101001101;
        end
        958: begin
            cosine_reg0 <= 36'sb11001110111111011011011101011001;
            sine_reg0   <= 36'sb11111110101100000110100101101101001;
        end
        959: begin
            cosine_reg0 <= 36'sb11001011110111011000011001010101;
            sine_reg0   <= 36'sb11111110101110100111111011101001111;
        end
        960: begin
            cosine_reg0 <= 36'sb11001000101111010011010111100001;
            sine_reg0   <= 36'sb11111110110001000110110100011110011;
        end
        961: begin
            cosine_reg0 <= 36'sb11000101100111001100011001111000;
            sine_reg0   <= 36'sb11111110110011100011010000001001001;
        end
        962: begin
            cosine_reg0 <= 36'sb11000010011111000011100010010110;
            sine_reg0   <= 36'sb11111110110101111101001110101000100;
        end
        963: begin
            cosine_reg0 <= 36'sb10111111010110111000110010110110;
            sine_reg0   <= 36'sb11111110111000010100101111111011001;
        end
        964: begin
            cosine_reg0 <= 36'sb10111100001110101100001101010011;
            sine_reg0   <= 36'sb11111110111010101001110011111111011;
        end
        965: begin
            cosine_reg0 <= 36'sb10111001000110011101110011101001;
            sine_reg0   <= 36'sb11111110111100111100011010110100001;
        end
        966: begin
            cosine_reg0 <= 36'sb10110101111110001101100111110100;
            sine_reg0   <= 36'sb11111110111111001100100100010111101;
        end
        967: begin
            cosine_reg0 <= 36'sb10110010110101111011101011101110;
            sine_reg0   <= 36'sb11111111000001011010010000101000101;
        end
        968: begin
            cosine_reg0 <= 36'sb10101111101101101000000001010101;
            sine_reg0   <= 36'sb11111111000011100101011111100101110;
        end
        969: begin
            cosine_reg0 <= 36'sb10101100100101010010101010100010;
            sine_reg0   <= 36'sb11111111000101101110010001001101110;
        end
        970: begin
            cosine_reg0 <= 36'sb10101001011100111011101001010010;
            sine_reg0   <= 36'sb11111111000111110100100101011111001;
        end
        971: begin
            cosine_reg0 <= 36'sb10100110010100100010111111100001;
            sine_reg0   <= 36'sb11111111001001111000011100011000110;
        end
        972: begin
            cosine_reg0 <= 36'sb10100011001100001000101111001001;
            sine_reg0   <= 36'sb11111111001011111001110101111001011;
        end
        973: begin
            cosine_reg0 <= 36'sb10100000000011101100111010000111;
            sine_reg0   <= 36'sb11111111001101111000110001111111100;
        end
        974: begin
            cosine_reg0 <= 36'sb10011100111011001111100010010110;
            sine_reg0   <= 36'sb11111111001111110101010000101010001;
        end
        975: begin
            cosine_reg0 <= 36'sb10011001110010110000101001110010;
            sine_reg0   <= 36'sb11111111010001101111010001111000000;
        end
        976: begin
            cosine_reg0 <= 36'sb10010110101010010000010010010110;
            sine_reg0   <= 36'sb11111111010011100110110101100111111;
        end
        977: begin
            cosine_reg0 <= 36'sb10010011100001101110011101111111;
            sine_reg0   <= 36'sb11111111010101011011111011111000110;
        end
        978: begin
            cosine_reg0 <= 36'sb10010000011001001011001110100111;
            sine_reg0   <= 36'sb11111111010111001110100100101001011;
        end
        979: begin
            cosine_reg0 <= 36'sb10001101010000100110100110001011;
            sine_reg0   <= 36'sb11111111011000111110101111111000101;
        end
        980: begin
            cosine_reg0 <= 36'sb10001010001000000000100110100111;
            sine_reg0   <= 36'sb11111111011010101100011101100101101;
        end
        981: begin
            cosine_reg0 <= 36'sb10000110111111011001010001110101;
            sine_reg0   <= 36'sb11111111011100010111101101101111000;
        end
        982: begin
            cosine_reg0 <= 36'sb10000011110110110000101001110010;
            sine_reg0   <= 36'sb11111111011110000000100000010100000;
        end
        983: begin
            cosine_reg0 <= 36'sb10000000101110000110110000011010;
            sine_reg0   <= 36'sb11111111011111100110110101010011011;
        end
        984: begin
            cosine_reg0 <= 36'sb1111101100101011011100111101000;
            sine_reg0   <= 36'sb11111111100001001010101100101100011;
        end
        985: begin
            cosine_reg0 <= 36'sb1111010011100101111010001011000;
            sine_reg0   <= 36'sb11111111100010101100000110011101111;
        end
        986: begin
            cosine_reg0 <= 36'sb1110111010100000001101111100110;
            sine_reg0   <= 36'sb11111111100100001011000010100110111;
        end
        987: begin
            cosine_reg0 <= 36'sb1110100001011010011000100001110;
            sine_reg0   <= 36'sb11111111100101100111100001000110110;
        end
        988: begin
            cosine_reg0 <= 36'sb1110001000010100011010001001011;
            sine_reg0   <= 36'sb11111111100111000001100001111100010;
        end
        989: begin
            cosine_reg0 <= 36'sb1101101111001110010011000011010;
            sine_reg0   <= 36'sb11111111101000011001000101000110111;
        end
        990: begin
            cosine_reg0 <= 36'sb1101010110001000000011011110101;
            sine_reg0   <= 36'sb11111111101001101110001010100101011;
        end
        991: begin
            cosine_reg0 <= 36'sb1100111101000001101011101011010;
            sine_reg0   <= 36'sb11111111101011000000110010010111011;
        end
        992: begin
            cosine_reg0 <= 36'sb1100100011111011001011111000100;
            sine_reg0   <= 36'sb11111111101100010000111100011011101;
        end
        993: begin
            cosine_reg0 <= 36'sb1100001010110100100100010101111;
            sine_reg0   <= 36'sb11111111101101011110101000110001110;
        end
        994: begin
            cosine_reg0 <= 36'sb1011110001101101110101010010110;
            sine_reg0   <= 36'sb11111111101110101001110111011000110;
        end
        995: begin
            cosine_reg0 <= 36'sb1011011000100110111110111110110;
            sine_reg0   <= 36'sb11111111101111110010101000010000000;
        end
        996: begin
            cosine_reg0 <= 36'sb1010111111100000000001101001010;
            sine_reg0   <= 36'sb11111111110000111000111011010110110;
        end
        997: begin
            cosine_reg0 <= 36'sb1010100110011000111101100001111;
            sine_reg0   <= 36'sb11111111110001111100110000101100011;
        end
        998: begin
            cosine_reg0 <= 36'sb1010001101010001110010111000000;
            sine_reg0   <= 36'sb11111111110010111110001000010000001;
        end
        999: begin
            cosine_reg0 <= 36'sb1001110100001010100001111011001;
            sine_reg0   <= 36'sb11111111110011111101000010000001100;
        end
        1000: begin
            cosine_reg0 <= 36'sb1001011011000011001010111010110;
            sine_reg0   <= 36'sb11111111110100111001011101111111111;
        end
        1001: begin
            cosine_reg0 <= 36'sb1001000001111011101110000110100;
            sine_reg0   <= 36'sb11111111110101110011011100001010100;
        end
        1002: begin
            cosine_reg0 <= 36'sb1000101000110100001011101101101;
            sine_reg0   <= 36'sb11111111110110101010111100100001000;
        end
        1003: begin
            cosine_reg0 <= 36'sb1000001111101100100011111111110;
            sine_reg0   <= 36'sb11111111110111011111111111000010111;
        end
        1004: begin
            cosine_reg0 <= 36'sb111110110100100110111001100100;
            sine_reg0   <= 36'sb11111111111000010010100011101111011;
        end
        1005: begin
            cosine_reg0 <= 36'sb111011101011101000101100011001;
            sine_reg0   <= 36'sb11111111111001000010101010100110010;
        end
        1006: begin
            cosine_reg0 <= 36'sb111000100010101001111010011010;
            sine_reg0   <= 36'sb11111111111001110000010011100111000;
        end
        1007: begin
            cosine_reg0 <= 36'sb110101011001101010100101100011;
            sine_reg0   <= 36'sb11111111111010011011011110110001000;
        end
        1008: begin
            cosine_reg0 <= 36'sb110010010000101010101111101111;
            sine_reg0   <= 36'sb11111111111011000100001100000100000;
        end
        1009: begin
            cosine_reg0 <= 36'sb101111000111101010011010111100;
            sine_reg0   <= 36'sb11111111111011101010011011011111101;
        end
        1010: begin
            cosine_reg0 <= 36'sb101011111110101001101001000100;
            sine_reg0   <= 36'sb11111111111100001110001101000011011;
        end
        1011: begin
            cosine_reg0 <= 36'sb101000110101101000011100000100;
            sine_reg0   <= 36'sb11111111111100101111100000101111000;
        end
        1012: begin
            cosine_reg0 <= 36'sb100101101100100110110101111000;
            sine_reg0   <= 36'sb11111111111101001110010110100010010;
        end
        1013: begin
            cosine_reg0 <= 36'sb100010100011100100111000011011;
            sine_reg0   <= 36'sb11111111111101101010101110011100101;
        end
        1014: begin
            cosine_reg0 <= 36'sb11111011010100010100101101011;
            sine_reg0   <= 36'sb11111111111110000100101000011110000;
        end
        1015: begin
            cosine_reg0 <= 36'sb11100010001011111111111100010;
            sine_reg0   <= 36'sb11111111111110011100000100100110001;
        end
        1016: begin
            cosine_reg0 <= 36'sb11001001000011101000111111101;
            sine_reg0   <= 36'sb11111111111110110001000010110100110;
        end
        1017: begin
            cosine_reg0 <= 36'sb10101111111011010000000111000;
            sine_reg0   <= 36'sb11111111111111000011100011001001101;
        end
        1018: begin
            cosine_reg0 <= 36'sb10010110110010110101100001110;
            sine_reg0   <= 36'sb11111111111111010011100101100100101;
        end
        1019: begin
            cosine_reg0 <= 36'sb1111101101010011001011111101;
            sine_reg0   <= 36'sb11111111111111100001001010000101100;
        end
        1020: begin
            cosine_reg0 <= 36'sb1100100100001111100001111111;
            sine_reg0   <= 36'sb11111111111111101100010000101100011;
        end
        1021: begin
            cosine_reg0 <= 36'sb1001011011001011110000010001;
            sine_reg0   <= 36'sb11111111111111110100111001011000111;
        end
        1022: begin
            cosine_reg0 <= 36'sb110010010000111111000110000;
            sine_reg0   <= 36'sb11111111111111111011000100001011000;
        end
        1023: begin
            cosine_reg0 <= 36'sb11001001000011111101010110;
            sine_reg0   <= 36'sb11111111111111111110110001000010101;
        end
        1024: begin
            cosine_reg0 <= 36'sb0;
            sine_reg0   <= 36'sb11111111111111111111111111111111111;
        end
        1025: begin
            cosine_reg0 <= 36'sb111111111100110110111100000010101010;
            sine_reg0   <= 36'sb11111111111111111110110001000010101;
        end
        1026: begin
            cosine_reg0 <= 36'sb111111111001101101111000000111010000;
            sine_reg0   <= 36'sb11111111111111111011000100001011000;
        end
        1027: begin
            cosine_reg0 <= 36'sb111111110110100100110100001111101111;
            sine_reg0   <= 36'sb11111111111111110100111001011000111;
        end
        1028: begin
            cosine_reg0 <= 36'sb111111110011011011110000011110000001;
            sine_reg0   <= 36'sb11111111111111101100010000101100011;
        end
        1029: begin
            cosine_reg0 <= 36'sb111111110000010010101100110100000011;
            sine_reg0   <= 36'sb11111111111111100001001010000101100;
        end
        1030: begin
            cosine_reg0 <= 36'sb111111101101001001101001010011110010;
            sine_reg0   <= 36'sb11111111111111010011100101100100101;
        end
        1031: begin
            cosine_reg0 <= 36'sb111111101010000000100101111111001000;
            sine_reg0   <= 36'sb11111111111111000011100011001001101;
        end
        1032: begin
            cosine_reg0 <= 36'sb111111100110110111100010111000000011;
            sine_reg0   <= 36'sb11111111111110110001000010110100110;
        end
        1033: begin
            cosine_reg0 <= 36'sb111111100011101110100000000000011110;
            sine_reg0   <= 36'sb11111111111110011100000100100110001;
        end
        1034: begin
            cosine_reg0 <= 36'sb111111100000100101011101011010010101;
            sine_reg0   <= 36'sb11111111111110000100101000011110000;
        end
        1035: begin
            cosine_reg0 <= 36'sb111111011101011100011011000111100101;
            sine_reg0   <= 36'sb11111111111101101010101110011100101;
        end
        1036: begin
            cosine_reg0 <= 36'sb111111011010010011011001001010001000;
            sine_reg0   <= 36'sb11111111111101001110010110100010010;
        end
        1037: begin
            cosine_reg0 <= 36'sb111111010111001010010111100011111100;
            sine_reg0   <= 36'sb11111111111100101111100000101111000;
        end
        1038: begin
            cosine_reg0 <= 36'sb111111010100000001010110010110111100;
            sine_reg0   <= 36'sb11111111111100001110001101000011011;
        end
        1039: begin
            cosine_reg0 <= 36'sb111111010000111000010101100101000100;
            sine_reg0   <= 36'sb11111111111011101010011011011111101;
        end
        1040: begin
            cosine_reg0 <= 36'sb111111001101101111010101010000010001;
            sine_reg0   <= 36'sb11111111111011000100001100000100000;
        end
        1041: begin
            cosine_reg0 <= 36'sb111111001010100110010101011010011101;
            sine_reg0   <= 36'sb11111111111010011011011110110001000;
        end
        1042: begin
            cosine_reg0 <= 36'sb111111000111011101010110000101100110;
            sine_reg0   <= 36'sb11111111111001110000010011100111000;
        end
        1043: begin
            cosine_reg0 <= 36'sb111111000100010100010111010011100111;
            sine_reg0   <= 36'sb11111111111001000010101010100110010;
        end
        1044: begin
            cosine_reg0 <= 36'sb111111000001001011011001000110011100;
            sine_reg0   <= 36'sb11111111111000010010100011101111011;
        end
        1045: begin
            cosine_reg0 <= 36'sb111110111110000010011011100000000010;
            sine_reg0   <= 36'sb11111111110111011111111111000010111;
        end
        1046: begin
            cosine_reg0 <= 36'sb111110111010111001011110100010010011;
            sine_reg0   <= 36'sb11111111110110101010111100100001000;
        end
        1047: begin
            cosine_reg0 <= 36'sb111110110111110000100010001111001100;
            sine_reg0   <= 36'sb11111111110101110011011100001010100;
        end
        1048: begin
            cosine_reg0 <= 36'sb111110110100100111100110101000101010;
            sine_reg0   <= 36'sb11111111110100111001011101111111111;
        end
        1049: begin
            cosine_reg0 <= 36'sb111110110001011110101011110000100111;
            sine_reg0   <= 36'sb11111111110011111101000010000001100;
        end
        1050: begin
            cosine_reg0 <= 36'sb111110101110010101110001101001000000;
            sine_reg0   <= 36'sb11111111110010111110001000010000001;
        end
        1051: begin
            cosine_reg0 <= 36'sb111110101011001100111000010011110001;
            sine_reg0   <= 36'sb11111111110001111100110000101100011;
        end
        1052: begin
            cosine_reg0 <= 36'sb111110101000000011111111110010110110;
            sine_reg0   <= 36'sb11111111110000111000111011010110110;
        end
        1053: begin
            cosine_reg0 <= 36'sb111110100100111011001000001000001010;
            sine_reg0   <= 36'sb11111111101111110010101000010000000;
        end
        1054: begin
            cosine_reg0 <= 36'sb111110100001110010010001010101101010;
            sine_reg0   <= 36'sb11111111101110101001110111011000110;
        end
        1055: begin
            cosine_reg0 <= 36'sb111110011110101001011011011101010001;
            sine_reg0   <= 36'sb11111111101101011110101000110001110;
        end
        1056: begin
            cosine_reg0 <= 36'sb111110011011100000100110100000111100;
            sine_reg0   <= 36'sb11111111101100010000111100011011101;
        end
        1057: begin
            cosine_reg0 <= 36'sb111110011000010111110010100010100110;
            sine_reg0   <= 36'sb11111111101011000000110010010111011;
        end
        1058: begin
            cosine_reg0 <= 36'sb111110010101001110111111100100001011;
            sine_reg0   <= 36'sb11111111101001101110001010100101011;
        end
        1059: begin
            cosine_reg0 <= 36'sb111110010010000110001101100111100110;
            sine_reg0   <= 36'sb11111111101000011001000101000110111;
        end
        1060: begin
            cosine_reg0 <= 36'sb111110001110111101011100101110110101;
            sine_reg0   <= 36'sb11111111100111000001100001111100010;
        end
        1061: begin
            cosine_reg0 <= 36'sb111110001011110100101100111011110010;
            sine_reg0   <= 36'sb11111111100101100111100001000110110;
        end
        1062: begin
            cosine_reg0 <= 36'sb111110001000101011111110010000011010;
            sine_reg0   <= 36'sb11111111100100001011000010100110111;
        end
        1063: begin
            cosine_reg0 <= 36'sb111110000101100011010000101110101000;
            sine_reg0   <= 36'sb11111111100010101100000110011101111;
        end
        1064: begin
            cosine_reg0 <= 36'sb111110000010011010100100011000011000;
            sine_reg0   <= 36'sb11111111100001001010101100101100011;
        end
        1065: begin
            cosine_reg0 <= 36'sb111101111111010001111001001111100110;
            sine_reg0   <= 36'sb11111111011111100110110101010011011;
        end
        1066: begin
            cosine_reg0 <= 36'sb111101111100001001001111010110001110;
            sine_reg0   <= 36'sb11111111011110000000100000010100000;
        end
        1067: begin
            cosine_reg0 <= 36'sb111101111001000000100110101110001011;
            sine_reg0   <= 36'sb11111111011100010111101101101111000;
        end
        1068: begin
            cosine_reg0 <= 36'sb111101110101110111111111011001011001;
            sine_reg0   <= 36'sb11111111011010101100011101100101101;
        end
        1069: begin
            cosine_reg0 <= 36'sb111101110010101111011001011001110101;
            sine_reg0   <= 36'sb11111111011000111110101111111000101;
        end
        1070: begin
            cosine_reg0 <= 36'sb111101101111100110110100110001011001;
            sine_reg0   <= 36'sb11111111010111001110100100101001011;
        end
        1071: begin
            cosine_reg0 <= 36'sb111101101100011110010001100010000001;
            sine_reg0   <= 36'sb11111111010101011011111011111000110;
        end
        1072: begin
            cosine_reg0 <= 36'sb111101101001010101101111101101101010;
            sine_reg0   <= 36'sb11111111010011100110110101100111111;
        end
        1073: begin
            cosine_reg0 <= 36'sb111101100110001101001111010110001110;
            sine_reg0   <= 36'sb11111111010001101111010001111000000;
        end
        1074: begin
            cosine_reg0 <= 36'sb111101100011000100110000011101101010;
            sine_reg0   <= 36'sb11111111001111110101010000101010001;
        end
        1075: begin
            cosine_reg0 <= 36'sb111101011111111100010011000101111001;
            sine_reg0   <= 36'sb11111111001101111000110001111111100;
        end
        1076: begin
            cosine_reg0 <= 36'sb111101011100110011110111010000110111;
            sine_reg0   <= 36'sb11111111001011111001110101111001011;
        end
        1077: begin
            cosine_reg0 <= 36'sb111101011001101011011101000000011111;
            sine_reg0   <= 36'sb11111111001001111000011100011000110;
        end
        1078: begin
            cosine_reg0 <= 36'sb111101010110100011000100010110101110;
            sine_reg0   <= 36'sb11111111000111110100100101011111001;
        end
        1079: begin
            cosine_reg0 <= 36'sb111101010011011010101101010101011110;
            sine_reg0   <= 36'sb11111111000101101110010001001101110;
        end
        1080: begin
            cosine_reg0 <= 36'sb111101010000010010010111111110101011;
            sine_reg0   <= 36'sb11111111000011100101011111100101110;
        end
        1081: begin
            cosine_reg0 <= 36'sb111101001101001010000100010100010010;
            sine_reg0   <= 36'sb11111111000001011010010000101000101;
        end
        1082: begin
            cosine_reg0 <= 36'sb111101001010000001110010011000001100;
            sine_reg0   <= 36'sb11111110111111001100100100010111101;
        end
        1083: begin
            cosine_reg0 <= 36'sb111101000110111001100010001100010111;
            sine_reg0   <= 36'sb11111110111100111100011010110100001;
        end
        1084: begin
            cosine_reg0 <= 36'sb111101000011110001010011110010101101;
            sine_reg0   <= 36'sb11111110111010101001110011111111011;
        end
        1085: begin
            cosine_reg0 <= 36'sb111101000000101001000111001101001010;
            sine_reg0   <= 36'sb11111110111000010100101111111011001;
        end
        1086: begin
            cosine_reg0 <= 36'sb111100111101100000111100011101101010;
            sine_reg0   <= 36'sb11111110110101111101001110101000100;
        end
        1087: begin
            cosine_reg0 <= 36'sb111100111010011000110011100110001000;
            sine_reg0   <= 36'sb11111110110011100011010000001001001;
        end
        1088: begin
            cosine_reg0 <= 36'sb111100110111010000101100101000011111;
            sine_reg0   <= 36'sb11111110110001000110110100011110011;
        end
        1089: begin
            cosine_reg0 <= 36'sb111100110100001000100111100110101011;
            sine_reg0   <= 36'sb11111110101110100111111011101001111;
        end
        1090: begin
            cosine_reg0 <= 36'sb111100110001000000100100100010100111;
            sine_reg0   <= 36'sb11111110101100000110100101101101001;
        end
        1091: begin
            cosine_reg0 <= 36'sb111100101101111000100011011110001111;
            sine_reg0   <= 36'sb11111110101001100010110010101001101;
        end
        1092: begin
            cosine_reg0 <= 36'sb111100101010110000100100011011011110;
            sine_reg0   <= 36'sb11111110100110111100100010100001000;
        end
        1093: begin
            cosine_reg0 <= 36'sb111100100111101000100111011100001111;
            sine_reg0   <= 36'sb11111110100100010011110101010100110;
        end
        1094: begin
            cosine_reg0 <= 36'sb111100100100100000101100100010011110;
            sine_reg0   <= 36'sb11111110100001101000101011000110101;
        end
        1095: begin
            cosine_reg0 <= 36'sb111100100001011000110011110000000111;
            sine_reg0   <= 36'sb11111110011110111011000011111000010;
        end
        1096: begin
            cosine_reg0 <= 36'sb111100011110010000111101000111000011;
            sine_reg0   <= 36'sb11111110011100001010111111101011010;
        end
        1097: begin
            cosine_reg0 <= 36'sb111100011011001001001000101001001111;
            sine_reg0   <= 36'sb11111110011001011000011110100001100;
        end
        1098: begin
            cosine_reg0 <= 36'sb111100011000000001010110011000100111;
            sine_reg0   <= 36'sb11111110010110100011100000011100011;
        end
        1099: begin
            cosine_reg0 <= 36'sb111100010100111001100110010111000100;
            sine_reg0   <= 36'sb11111110010011101100000101011110000;
        end
        1100: begin
            cosine_reg0 <= 36'sb111100010001110001111000100110100011;
            sine_reg0   <= 36'sb11111110010000110010001101100111111;
        end
        1101: begin
            cosine_reg0 <= 36'sb111100001110101010001101001000111110;
            sine_reg0   <= 36'sb11111110001101110101111000111011111;
        end
        1102: begin
            cosine_reg0 <= 36'sb111100001011100010100100000000010001;
            sine_reg0   <= 36'sb11111110001010110111000111011011110;
        end
        1103: begin
            cosine_reg0 <= 36'sb111100001000011010111101001110010111;
            sine_reg0   <= 36'sb11111110000111110101111001001001100;
        end
        1104: begin
            cosine_reg0 <= 36'sb111100000101010011011000110101001011;
            sine_reg0   <= 36'sb11111110000100110010001110000110111;
        end
        1105: begin
            cosine_reg0 <= 36'sb111100000010001011110110110110101000;
            sine_reg0   <= 36'sb11111110000001101100000110010101111;
        end
        1106: begin
            cosine_reg0 <= 36'sb111011111111000100010111010100101001;
            sine_reg0   <= 36'sb11111101111110100011100001111000010;
        end
        1107: begin
            cosine_reg0 <= 36'sb111011111011111100111010010001001010;
            sine_reg0   <= 36'sb11111101111011011000100000110000000;
        end
        1108: begin
            cosine_reg0 <= 36'sb111011111000110101011111101110000100;
            sine_reg0   <= 36'sb11111101111000001011000010111111000;
        end
        1109: begin
            cosine_reg0 <= 36'sb111011110101101110000111101101010101;
            sine_reg0   <= 36'sb11111101110100111011001000100111011;
        end
        1110: begin
            cosine_reg0 <= 36'sb111011110010100110110010010000110101;
            sine_reg0   <= 36'sb11111101110001101000110001101011001;
        end
        1111: begin
            cosine_reg0 <= 36'sb111011101111011111011111011010100001;
            sine_reg0   <= 36'sb11111101101110010011111110001100001;
        end
        1112: begin
            cosine_reg0 <= 36'sb111011101100011000001111001100010010;
            sine_reg0   <= 36'sb11111101101010111100101110001100100;
        end
        1113: begin
            cosine_reg0 <= 36'sb111011101001010001000001101000000101;
            sine_reg0   <= 36'sb11111101100111100011000001101110100;
        end
        1114: begin
            cosine_reg0 <= 36'sb111011100110001001110110101111110100;
            sine_reg0   <= 36'sb11111101100100000110111000110011111;
        end
        1115: begin
            cosine_reg0 <= 36'sb111011100011000010101110100101011010;
            sine_reg0   <= 36'sb11111101100000101000010011011111001;
        end
        1116: begin
            cosine_reg0 <= 36'sb111011011111111011101001001010110001;
            sine_reg0   <= 36'sb11111101011101000111010001110010001;
        end
        1117: begin
            cosine_reg0 <= 36'sb111011011100110100100110100001110101;
            sine_reg0   <= 36'sb11111101011001100011110011101111001;
        end
        1118: begin
            cosine_reg0 <= 36'sb111011011001101101100110101100100000;
            sine_reg0   <= 36'sb11111101010101111101111001011000010;
        end
        1119: begin
            cosine_reg0 <= 36'sb111011010110100110101001101100101101;
            sine_reg0   <= 36'sb11111101010010010101100010101111111;
        end
        1120: begin
            cosine_reg0 <= 36'sb111011010011011111101111100100010111;
            sine_reg0   <= 36'sb11111101001110101010101111111000001;
        end
        1121: begin
            cosine_reg0 <= 36'sb111011010000011000111000010101011000;
            sine_reg0   <= 36'sb11111101001010111101100000110011011;
        end
        1122: begin
            cosine_reg0 <= 36'sb111011001101010010000100000001101100;
            sine_reg0   <= 36'sb11111101000111001101110101100011110;
        end
        1123: begin
            cosine_reg0 <= 36'sb111011001010001011010010101011001100;
            sine_reg0   <= 36'sb11111101000011011011101110001011101;
        end
        1124: begin
            cosine_reg0 <= 36'sb111011000111000100100100010011110011;
            sine_reg0   <= 36'sb11111100111111100111001010101101010;
        end
        1125: begin
            cosine_reg0 <= 36'sb111011000011111101111000111101011101;
            sine_reg0   <= 36'sb11111100111011110000001011001011010;
        end
        1126: begin
            cosine_reg0 <= 36'sb111011000000110111010000101010000010;
            sine_reg0   <= 36'sb11111100110111110110101111100111110;
        end
        1127: begin
            cosine_reg0 <= 36'sb111010111101110000101011011011011111;
            sine_reg0   <= 36'sb11111100110011111010111000000101010;
        end
        1128: begin
            cosine_reg0 <= 36'sb111010111010101010001001010011101110;
            sine_reg0   <= 36'sb11111100101111111100100100100110001;
        end
        1129: begin
            cosine_reg0 <= 36'sb111010110111100011101010010100101000;
            sine_reg0   <= 36'sb11111100101011111011110101001100111;
        end
        1130: begin
            cosine_reg0 <= 36'sb111010110100011101001110100000001001;
            sine_reg0   <= 36'sb11111100100111111000101001111100000;
        end
        1131: begin
            cosine_reg0 <= 36'sb111010110001010110110101111000001010;
            sine_reg0   <= 36'sb11111100100011110011000010110110000;
        end
        1132: begin
            cosine_reg0 <= 36'sb111010101110010000100000011110100111;
            sine_reg0   <= 36'sb11111100011111101010111111111101011;
        end
        1133: begin
            cosine_reg0 <= 36'sb111010101011001010001110010101011001;
            sine_reg0   <= 36'sb11111100011011100000100001010100100;
        end
        1134: begin
            cosine_reg0 <= 36'sb111010101000000011111111011110011011;
            sine_reg0   <= 36'sb11111100010111010011100110111110010;
        end
        1135: begin
            cosine_reg0 <= 36'sb111010100100111101110011111011100111;
            sine_reg0   <= 36'sb11111100010011000100010000111101000;
        end
        1136: begin
            cosine_reg0 <= 36'sb111010100001110111101011101110110111;
            sine_reg0   <= 36'sb11111100001110110010011111010011011;
        end
        1137: begin
            cosine_reg0 <= 36'sb111010011110110001100110111010000111;
            sine_reg0   <= 36'sb11111100001010011110010010000100001;
        end
        1138: begin
            cosine_reg0 <= 36'sb111010011011101011100101011111001110;
            sine_reg0   <= 36'sb11111100000110000111101001010001111;
        end
        1139: begin
            cosine_reg0 <= 36'sb111010011000100101100111100000001001;
            sine_reg0   <= 36'sb11111100000001101110100100111111010;
        end
        1140: begin
            cosine_reg0 <= 36'sb111010010101011111101100111110110001;
            sine_reg0   <= 36'sb11111011111101010011000101001111001;
        end
        1141: begin
            cosine_reg0 <= 36'sb111010010010011001110101111101000000;
            sine_reg0   <= 36'sb11111011111000110101001010000100000;
        end
        1142: begin
            cosine_reg0 <= 36'sb111010001111010100000010011100110000;
            sine_reg0   <= 36'sb11111011110100010100110011100000110;
        end
        1143: begin
            cosine_reg0 <= 36'sb111010001100001110010010011111111011;
            sine_reg0   <= 36'sb11111011101111110010000001101000001;
        end
        1144: begin
            cosine_reg0 <= 36'sb111010001001001000100110001000011011;
            sine_reg0   <= 36'sb11111011101011001100110100011100111;
        end
        1145: begin
            cosine_reg0 <= 36'sb111010000110000010111101011000001011;
            sine_reg0   <= 36'sb11111011100110100101001100000010000;
        end
        1146: begin
            cosine_reg0 <= 36'sb111010000010111101011000010001000011;
            sine_reg0   <= 36'sb11111011100001111011001000011010010;
        end
        1147: begin
            cosine_reg0 <= 36'sb111001111111110111110110110100111110;
            sine_reg0   <= 36'sb11111011011101001110101001101000100;
        end
        1148: begin
            cosine_reg0 <= 36'sb111001111100110010011001000101110110;
            sine_reg0   <= 36'sb11111011011000011111101111101111100;
        end
        1149: begin
            cosine_reg0 <= 36'sb111001111001101100111111000101100101;
            sine_reg0   <= 36'sb11111011010011101110011010110010100;
        end
        1150: begin
            cosine_reg0 <= 36'sb111001110110100111101000110110000100;
            sine_reg0   <= 36'sb11111011001110111010101010110100001;
        end
        1151: begin
            cosine_reg0 <= 36'sb111001110011100010010110011001001101;
            sine_reg0   <= 36'sb11111011001010000100011111110111100;
        end
        1152: begin
            cosine_reg0 <= 36'sb111001110000011101000111110000111010;
            sine_reg0   <= 36'sb11111011000101001011111001111111101;
        end
        1153: begin
            cosine_reg0 <= 36'sb111001101101010111111100111111000100;
            sine_reg0   <= 36'sb11111011000000010000111001001111011;
        end
        1154: begin
            cosine_reg0 <= 36'sb111001101010010010110110000101100101;
            sine_reg0   <= 36'sb11111010111011010011011101101010000;
        end
        1155: begin
            cosine_reg0 <= 36'sb111001100111001101110011000110010111;
            sine_reg0   <= 36'sb11111010110110010011100111010010011;
        end
        1156: begin
            cosine_reg0 <= 36'sb111001100100001000110100000011010010;
            sine_reg0   <= 36'sb11111010110001010001010110001011101;
        end
        1157: begin
            cosine_reg0 <= 36'sb111001100001000011111000111110010010;
            sine_reg0   <= 36'sb11111010101100001100101010011000111;
        end
        1158: begin
            cosine_reg0 <= 36'sb111001011101111111000001111001001111;
            sine_reg0   <= 36'sb11111010100111000101100011111101011;
        end
        1159: begin
            cosine_reg0 <= 36'sb111001011010111010001110110110000010;
            sine_reg0   <= 36'sb11111010100001111100000010111100000;
        end
        1160: begin
            cosine_reg0 <= 36'sb111001010111110101011111110110100101;
            sine_reg0   <= 36'sb11111010011100110000000111011000010;
        end
        1161: begin
            cosine_reg0 <= 36'sb111001010100110000110100111100110010;
            sine_reg0   <= 36'sb11111010010111100001110001010101000;
        end
        1162: begin
            cosine_reg0 <= 36'sb111001010001101100001110001010100001;
            sine_reg0   <= 36'sb11111010010010010001000000110101110;
        end
        1163: begin
            cosine_reg0 <= 36'sb111001001110100111101011100001101100;
            sine_reg0   <= 36'sb11111010001100111101110101111101101;
        end
        1164: begin
            cosine_reg0 <= 36'sb111001001011100011001101000100001100;
            sine_reg0   <= 36'sb11111010000111101000010000101111111;
        end
        1165: begin
            cosine_reg0 <= 36'sb111001001000011110110010110011111011;
            sine_reg0   <= 36'sb11111010000010010000010001001111110;
        end
        1166: begin
            cosine_reg0 <= 36'sb111001000101011010011100110010110001;
            sine_reg0   <= 36'sb11111001111100110101110111100000110;
        end
        1167: begin
            cosine_reg0 <= 36'sb111001000010010110001011000010101000;
            sine_reg0   <= 36'sb11111001110111011001000011100110000;
        end
        1168: begin
            cosine_reg0 <= 36'sb111000111111010001111101100101011000;
            sine_reg0   <= 36'sb11111001110001111001110101100011000;
        end
        1169: begin
            cosine_reg0 <= 36'sb111000111100001101110100011100111011;
            sine_reg0   <= 36'sb11111001101100011000001101011011001;
        end
        1170: begin
            cosine_reg0 <= 36'sb111000111001001001101111101011001010;
            sine_reg0   <= 36'sb11111001100110110100001011010001110;
        end
        1171: begin
            cosine_reg0 <= 36'sb111000110110000101101111010001111110;
            sine_reg0   <= 36'sb11111001100001001101101111001010010;
        end
        1172: begin
            cosine_reg0 <= 36'sb111000110011000001110011010011001111;
            sine_reg0   <= 36'sb11111001011011100100111001001000001;
        end
        1173: begin
            cosine_reg0 <= 36'sb111000101111111101111011110000110111;
            sine_reg0   <= 36'sb11111001010101111001101001001110111;
        end
        1174: begin
            cosine_reg0 <= 36'sb111000101100111010001000101100101101;
            sine_reg0   <= 36'sb11111001010000001011111111100010001;
        end
        1175: begin
            cosine_reg0 <= 36'sb111000101001110110011010001000101100;
            sine_reg0   <= 36'sb11111001001010011011111100000101001;
        end
        1176: begin
            cosine_reg0 <= 36'sb111000100110110010110000000110101100;
            sine_reg0   <= 36'sb11111001000100101001011110111011101;
        end
        1177: begin
            cosine_reg0 <= 36'sb111000100011101111001010101000100101;
            sine_reg0   <= 36'sb11111000111110110100101000001001000;
        end
        1178: begin
            cosine_reg0 <= 36'sb111000100000101011101001110000010000;
            sine_reg0   <= 36'sb11111000111000111101010111110001001;
        end
        1179: begin
            cosine_reg0 <= 36'sb111000011101101000001101011111100110;
            sine_reg0   <= 36'sb11111000110011000011101101110111100;
        end
        1180: begin
            cosine_reg0 <= 36'sb111000011010100100110101111000011111;
            sine_reg0   <= 36'sb11111000101101000111101010011111101;
        end
        1181: begin
            cosine_reg0 <= 36'sb111000010111100001100010111100110100;
            sine_reg0   <= 36'sb11111000100111001001001101101101010;
        end
        1182: begin
            cosine_reg0 <= 36'sb111000010100011110010100101110011101;
            sine_reg0   <= 36'sb11111000100001001000010111100100001;
        end
        1183: begin
            cosine_reg0 <= 36'sb111000010001011011001011001111010011;
            sine_reg0   <= 36'sb11111000011011000101001000001000000;
        end
        1184: begin
            cosine_reg0 <= 36'sb111000001110011000000110100001001110;
            sine_reg0   <= 36'sb11111000010100111111011111011100100;
        end
        1185: begin
            cosine_reg0 <= 36'sb111000001011010101000110100110000110;
            sine_reg0   <= 36'sb11111000001110110111011101100101011;
        end
        1186: begin
            cosine_reg0 <= 36'sb111000001000010010001011011111110100;
            sine_reg0   <= 36'sb11111000001000101101000010100110011;
        end
        1187: begin
            cosine_reg0 <= 36'sb111000000101001111010101010000010000;
            sine_reg0   <= 36'sb11111000000010100000001110100011011;
        end
        1188: begin
            cosine_reg0 <= 36'sb111000000010001100100011111001010010;
            sine_reg0   <= 36'sb11110111111100010001000001100000010;
        end
        1189: begin
            cosine_reg0 <= 36'sb110111111111001001110111011100110010;
            sine_reg0   <= 36'sb11110111110101111111011011100000110;
        end
        1190: begin
            cosine_reg0 <= 36'sb110111111100000111001111111100101001;
            sine_reg0   <= 36'sb11110111101111101011011100101000110;
        end
        1191: begin
            cosine_reg0 <= 36'sb110111111001000100101101011010101110;
            sine_reg0   <= 36'sb11110111101001010101000100111100010;
        end
        1192: begin
            cosine_reg0 <= 36'sb110111110110000010001111111000111001;
            sine_reg0   <= 36'sb11110111100010111100010100011111000;
        end
        1193: begin
            cosine_reg0 <= 36'sb110111110010111111110111011001000011;
            sine_reg0   <= 36'sb11110111011100100001001011010101001;
        end
        1194: begin
            cosine_reg0 <= 36'sb110111101111111101100011111101000011;
            sine_reg0   <= 36'sb11110111010110000011101001100010011;
        end
        1195: begin
            cosine_reg0 <= 36'sb110111101100111011010101100110110001;
            sine_reg0   <= 36'sb11110111001111100011101111001010111;
        end
        1196: begin
            cosine_reg0 <= 36'sb110111101001111001001100011000000101;
            sine_reg0   <= 36'sb11110111001001000001011100010010110;
        end
        1197: begin
            cosine_reg0 <= 36'sb110111100110110111001000010010110110;
            sine_reg0   <= 36'sb11110111000010011100110000111101110;
        end
        1198: begin
            cosine_reg0 <= 36'sb110111100011110101001001011000111101;
            sine_reg0   <= 36'sb11110110111011110101101101010000001;
        end
        1199: begin
            cosine_reg0 <= 36'sb110111100000110011001111101100010001;
            sine_reg0   <= 36'sb11110110110101001100010001001101111;
        end
        1200: begin
            cosine_reg0 <= 36'sb110111011101110001011011001110101010;
            sine_reg0   <= 36'sb11110110101110100000011100111011001;
        end
        1201: begin
            cosine_reg0 <= 36'sb110111011010101111101100000001111111;
            sine_reg0   <= 36'sb11110110100111110010010000011100000;
        end
        1202: begin
            cosine_reg0 <= 36'sb110111010111101110000010001000000111;
            sine_reg0   <= 36'sb11110110100001000001101011110100101;
        end
        1203: begin
            cosine_reg0 <= 36'sb110111010100101100011101100010111011;
            sine_reg0   <= 36'sb11110110011010001110101111001001010;
        end
        1204: begin
            cosine_reg0 <= 36'sb110111010001101010111110010100010001;
            sine_reg0   <= 36'sb11110110010011011001011010011110000;
        end
        1205: begin
            cosine_reg0 <= 36'sb110111001110101001100100011110000010;
            sine_reg0   <= 36'sb11110110001100100001101101110111001;
        end
        1206: begin
            cosine_reg0 <= 36'sb110111001011101000010000000010000011;
            sine_reg0   <= 36'sb11110110000101100111101001011000110;
        end
        1207: begin
            cosine_reg0 <= 36'sb110111001000100111000001000010001101;
            sine_reg0   <= 36'sb11110101111110101011001101000111010;
        end
        1208: begin
            cosine_reg0 <= 36'sb110111000101100101110111100000010111;
            sine_reg0   <= 36'sb11110101110111101100011001000110111;
        end
        1209: begin
            cosine_reg0 <= 36'sb110111000010100100110011011110010111;
            sine_reg0   <= 36'sb11110101110000101011001101011011111;
        end
        1210: begin
            cosine_reg0 <= 36'sb110110111111100011110100111110000101;
            sine_reg0   <= 36'sb11110101101001100111101010001010110;
        end
        1211: begin
            cosine_reg0 <= 36'sb110110111100100010111100000001011001;
            sine_reg0   <= 36'sb11110101100010100001101111010111101;
        end
        1212: begin
            cosine_reg0 <= 36'sb110110111001100010001000101010001000;
            sine_reg0   <= 36'sb11110101011011011001011101000111001;
        end
        1213: begin
            cosine_reg0 <= 36'sb110110110110100001011010111010001010;
            sine_reg0   <= 36'sb11110101010100001110110011011101100;
        end
        1214: begin
            cosine_reg0 <= 36'sb110110110011100000110010110011010110;
            sine_reg0   <= 36'sb11110101001101000001110010011111001;
        end
        1215: begin
            cosine_reg0 <= 36'sb110110110000100000010000010111100010;
            sine_reg0   <= 36'sb11110101000101110010011010010000100;
        end
        1216: begin
            cosine_reg0 <= 36'sb110110101101011111110011101000100110;
            sine_reg0   <= 36'sb11110100111110100000101010110110001;
        end
        1217: begin
            cosine_reg0 <= 36'sb110110101010011111011100101000010111;
            sine_reg0   <= 36'sb11110100110111001100100100010100011;
        end
        1218: begin
            cosine_reg0 <= 36'sb110110100111011111001011011000101110;
            sine_reg0   <= 36'sb11110100101111110110000110101111111;
        end
        1219: begin
            cosine_reg0 <= 36'sb110110100100011110111111111011011111;
            sine_reg0   <= 36'sb11110100101000011101010010001101010;
        end
        1220: begin
            cosine_reg0 <= 36'sb110110100001011110111010010010100011;
            sine_reg0   <= 36'sb11110100100001000010000110110000111;
        end
        1221: begin
            cosine_reg0 <= 36'sb110110011110011110111010011111101111;
            sine_reg0   <= 36'sb11110100011001100100100100011111010;
        end
        1222: begin
            cosine_reg0 <= 36'sb110110011011011111000000100100111001;
            sine_reg0   <= 36'sb11110100010010000100101011011101010;
        end
        1223: begin
            cosine_reg0 <= 36'sb110110011000011111001100100011111001;
            sine_reg0   <= 36'sb11110100001010100010011011101111011;
        end
        1224: begin
            cosine_reg0 <= 36'sb110110010101011111011110011110100100;
            sine_reg0   <= 36'sb11110100000010111101110101011010010;
        end
        1225: begin
            cosine_reg0 <= 36'sb110110010010011111110110010110110001;
            sine_reg0   <= 36'sb11110011111011010110111000100010101;
        end
        1226: begin
            cosine_reg0 <= 36'sb110110001111100000010100001110010110;
            sine_reg0   <= 36'sb11110011110011101101100101001101000;
        end
        1227: begin
            cosine_reg0 <= 36'sb110110001100100000111000000111001001;
            sine_reg0   <= 36'sb11110011101100000001111011011110011;
        end
        1228: begin
            cosine_reg0 <= 36'sb110110001001100001100010000011000000;
            sine_reg0   <= 36'sb11110011100100010011111011011011010;
        end
        1229: begin
            cosine_reg0 <= 36'sb110110000110100010010010000011110001;
            sine_reg0   <= 36'sb11110011011100100011100101001000100;
        end
        1230: begin
            cosine_reg0 <= 36'sb110110000011100011001000001011010010;
            sine_reg0   <= 36'sb11110011010100110000111000101010110;
        end
        1231: begin
            cosine_reg0 <= 36'sb110110000000100100000100011011011010;
            sine_reg0   <= 36'sb11110011001100111011110110000111001;
        end
        1232: begin
            cosine_reg0 <= 36'sb110101111101100101000110110101111101;
            sine_reg0   <= 36'sb11110011000101000100011101100010001;
        end
        1233: begin
            cosine_reg0 <= 36'sb110101111010100110001111011100110011;
            sine_reg0   <= 36'sb11110010111101001010101111000000111;
        end
        1234: begin
            cosine_reg0 <= 36'sb110101110111100111011110010001101111;
            sine_reg0   <= 36'sb11110010110101001110101010101000000;
        end
        1235: begin
            cosine_reg0 <= 36'sb110101110100101000110011010110101001;
            sine_reg0   <= 36'sb11110010101101010000010000011100101;
        end
        1236: begin
            cosine_reg0 <= 36'sb110101110001101010001110101101010101;
            sine_reg0   <= 36'sb11110010100101001111100000100011100;
        end
        1237: begin
            cosine_reg0 <= 36'sb110101101110101011110000010111101010;
            sine_reg0   <= 36'sb11110010011101001100011011000001101;
        end
        1238: begin
            cosine_reg0 <= 36'sb110101101011101101011000010111011101;
            sine_reg0   <= 36'sb11110010010101000110111111111100000;
        end
        1239: begin
            cosine_reg0 <= 36'sb110101101000101111000110101110100011;
            sine_reg0   <= 36'sb11110010001100111111001111010111100;
        end
        1240: begin
            cosine_reg0 <= 36'sb110101100101110000111011011110110001;
            sine_reg0   <= 36'sb11110010000100110101001001011001010;
        end
        1241: begin
            cosine_reg0 <= 36'sb110101100010110010110110101001111110;
            sine_reg0   <= 36'sb11110001111100101000101110000110010;
        end
        1242: begin
            cosine_reg0 <= 36'sb110101011111110100111000010001111101;
            sine_reg0   <= 36'sb11110001110100011001111101100011101;
        end
        1243: begin
            cosine_reg0 <= 36'sb110101011100110111000000011000100101;
            sine_reg0   <= 36'sb11110001101100001000110111110110010;
        end
        1244: begin
            cosine_reg0 <= 36'sb110101011001111001001110111111101010;
            sine_reg0   <= 36'sb11110001100011110101011101000011011;
        end
        1245: begin
            cosine_reg0 <= 36'sb110101010110111011100100001001000010;
            sine_reg0   <= 36'sb11110001011011011111101101010000001;
        end
        1246: begin
            cosine_reg0 <= 36'sb110101010011111101111111110110100010;
            sine_reg0   <= 36'sb11110001010011000111101000100001101;
        end
        1247: begin
            cosine_reg0 <= 36'sb110101010001000000100010001001111110;
            sine_reg0   <= 36'sb11110001001010101101001110111101001;
        end
        1248: begin
            cosine_reg0 <= 36'sb110101001110000011001011000101001011;
            sine_reg0   <= 36'sb11110001000010010000100000100111101;
        end
        1249: begin
            cosine_reg0 <= 36'sb110101001011000101111010101001111110;
            sine_reg0   <= 36'sb11110000111001110001011101100110011;
        end
        1250: begin
            cosine_reg0 <= 36'sb110101001000001000110000111010001101;
            sine_reg0   <= 36'sb11110000110001010000000101111110110;
        end
        1251: begin
            cosine_reg0 <= 36'sb110101000101001011101101110111101010;
            sine_reg0   <= 36'sb11110000101000101100011001110101111;
        end
        1252: begin
            cosine_reg0 <= 36'sb110101000010001110110001100100001101;
            sine_reg0   <= 36'sb11110000100000000110011001010001001;
        end
        1253: begin
            cosine_reg0 <= 36'sb110100111111010001111100000001100111;
            sine_reg0   <= 36'sb11110000010111011110000100010101110;
        end
        1254: begin
            cosine_reg0 <= 36'sb110100111100010101001101010001101111;
            sine_reg0   <= 36'sb11110000001110110011011011001001001;
        end
        1255: begin
            cosine_reg0 <= 36'sb110100111001011000100101010110011001;
            sine_reg0   <= 36'sb11110000000110000110011101110000100;
        end
        1256: begin
            cosine_reg0 <= 36'sb110100110110011100000100010001011000;
            sine_reg0   <= 36'sb11101111111101010111001100010001010;
        end
        1257: begin
            cosine_reg0 <= 36'sb110100110011011111101010000100100010;
            sine_reg0   <= 36'sb11101111110100100101100110110000111;
        end
        1258: begin
            cosine_reg0 <= 36'sb110100110000100011010110110001101011;
            sine_reg0   <= 36'sb11101111101011110001101101010100110;
        end
        1259: begin
            cosine_reg0 <= 36'sb110100101101100111001010011010100110;
            sine_reg0   <= 36'sb11101111100010111011100000000010010;
        end
        1260: begin
            cosine_reg0 <= 36'sb110100101010101011000101000001000111;
            sine_reg0   <= 36'sb11101111011010000010111110111110111;
        end
        1261: begin
            cosine_reg0 <= 36'sb110100100111101111000110100111000100;
            sine_reg0   <= 36'sb11101111010001001000001010010000000;
        end
        1262: begin
            cosine_reg0 <= 36'sb110100100100110011001111001110001111;
            sine_reg0   <= 36'sb11101111001000001011000001111011010;
        end
        1263: begin
            cosine_reg0 <= 36'sb110100100001110111011110111000011101;
            sine_reg0   <= 36'sb11101110111111001011100110000110010;
        end
        1264: begin
            cosine_reg0 <= 36'sb110100011110111011110101100111100001;
            sine_reg0   <= 36'sb11101110110110001001110110110110010;
        end
        1265: begin
            cosine_reg0 <= 36'sb110100011100000000010011011101001111;
            sine_reg0   <= 36'sb11101110101101000101110100010001001;
        end
        1266: begin
            cosine_reg0 <= 36'sb110100011001000100111000011011011100;
            sine_reg0   <= 36'sb11101110100011111111011110011100010;
        end
        1267: begin
            cosine_reg0 <= 36'sb110100010110001001100100100011111001;
            sine_reg0   <= 36'sb11101110011010110110110101011101010;
        end
        1268: begin
            cosine_reg0 <= 36'sb110100010011001110010111111000011100;
            sine_reg0   <= 36'sb11101110010001101011111001011001111;
        end
        1269: begin
            cosine_reg0 <= 36'sb110100010000010011010010011010110111;
            sine_reg0   <= 36'sb11101110001000011110101010010111110;
        end
        1270: begin
            cosine_reg0 <= 36'sb110100001101011000010100001100111110;
            sine_reg0   <= 36'sb11101101111111001111001000011100100;
        end
        1271: begin
            cosine_reg0 <= 36'sb110100001010011101011101010000100100;
            sine_reg0   <= 36'sb11101101110101111101010011101110000;
        end
        1272: begin
            cosine_reg0 <= 36'sb110100000111100010101101100111011101;
            sine_reg0   <= 36'sb11101101101100101001001100010001101;
        end
        1273: begin
            cosine_reg0 <= 36'sb110100000100101000000101010011011011;
            sine_reg0   <= 36'sb11101101100011010010110010001101100;
        end
        1274: begin
            cosine_reg0 <= 36'sb110100000001101101100100010110010010;
            sine_reg0   <= 36'sb11101101011001111010000101100111001;
        end
        1275: begin
            cosine_reg0 <= 36'sb110011111110110011001010110001110101;
            sine_reg0   <= 36'sb11101101010000011111000110100100011;
        end
        1276: begin
            cosine_reg0 <= 36'sb110011111011111000111000100111110111;
            sine_reg0   <= 36'sb11101101000111000001110101001011001;
        end
        1277: begin
            cosine_reg0 <= 36'sb110011111000111110101101111010001010;
            sine_reg0   <= 36'sb11101100111101100010010001100001001;
        end
        1278: begin
            cosine_reg0 <= 36'sb110011110110000100101010101010100010;
            sine_reg0   <= 36'sb11101100110100000000011011101100010;
        end
        1279: begin
            cosine_reg0 <= 36'sb110011110011001010101110111010110001;
            sine_reg0   <= 36'sb11101100101010011100010011110010011;
        end
        1280: begin
            cosine_reg0 <= 36'sb110011110000010000111010101100101011;
            sine_reg0   <= 36'sb11101100100000110101111001111001100;
        end
        1281: begin
            cosine_reg0 <= 36'sb110011101101010111001110000010000001;
            sine_reg0   <= 36'sb11101100010111001101001110000111011;
        end
        1282: begin
            cosine_reg0 <= 36'sb110011101010011101101000111100100110;
            sine_reg0   <= 36'sb11101100001101100010010000100010000;
        end
        1283: begin
            cosine_reg0 <= 36'sb110011100111100100001011011110001100;
            sine_reg0   <= 36'sb11101100000011110101000001001111100;
        end
        1284: begin
            cosine_reg0 <= 36'sb110011100100101010110101101000100111;
            sine_reg0   <= 36'sb11101011111010000101100000010101101;
        end
        1285: begin
            cosine_reg0 <= 36'sb110011100001110001100111011101101001;
            sine_reg0   <= 36'sb11101011110000010011101101111010101;
        end
        1286: begin
            cosine_reg0 <= 36'sb110011011110111000100000111111000010;
            sine_reg0   <= 36'sb11101011100110011111101010000100010;
        end
        1287: begin
            cosine_reg0 <= 36'sb110011011011111111100010001110100111;
            sine_reg0   <= 36'sb11101011011100101001010100111000110;
        end
        1288: begin
            cosine_reg0 <= 36'sb110011011001000110101011001110001001;
            sine_reg0   <= 36'sb11101011010010110000101110011110010;
        end
        1289: begin
            cosine_reg0 <= 36'sb110011010110001101111011111111011001;
            sine_reg0   <= 36'sb11101011001000110101110110111010101;
        end
        1290: begin
            cosine_reg0 <= 36'sb110011010011010101010100100100001011;
            sine_reg0   <= 36'sb11101010111110111000101110010100001;
        end
        1291: begin
            cosine_reg0 <= 36'sb110011010000011100110100111110001111;
            sine_reg0   <= 36'sb11101010110100111001010100110001000;
        end
        1292: begin
            cosine_reg0 <= 36'sb110011001101100100011101001111011000;
            sine_reg0   <= 36'sb11101010101010110111101010010111001;
        end
        1293: begin
            cosine_reg0 <= 36'sb110011001010101100001101011001010111;
            sine_reg0   <= 36'sb11101010100000110011101111001101000;
        end
        1294: begin
            cosine_reg0 <= 36'sb110011000111110100000101011101111111;
            sine_reg0   <= 36'sb11101010010110101101100011011000101;
        end
        1295: begin
            cosine_reg0 <= 36'sb110011000100111100000101011110111111;
            sine_reg0   <= 36'sb11101010001100100101000111000000011;
        end
        1296: begin
            cosine_reg0 <= 36'sb110011000010000100001101011110001011;
            sine_reg0   <= 36'sb11101010000010011010011010001010011;
        end
        1297: begin
            cosine_reg0 <= 36'sb110010111111001100011101011101010100;
            sine_reg0   <= 36'sb11101001111000001101011100111100111;
        end
        1298: begin
            cosine_reg0 <= 36'sb110010111100010100110101011110001010;
            sine_reg0   <= 36'sb11101001101101111110001111011110010;
        end
        1299: begin
            cosine_reg0 <= 36'sb110010111001011101010101100010011111;
            sine_reg0   <= 36'sb11101001100011101100110001110100111;
        end
        1300: begin
            cosine_reg0 <= 36'sb110010110110100101111101101100000101;
            sine_reg0   <= 36'sb11101001011001011001000100000110111;
        end
        1301: begin
            cosine_reg0 <= 36'sb110010110011101110101101111100101100;
            sine_reg0   <= 36'sb11101001001111000011000110011010111;
        end
        1302: begin
            cosine_reg0 <= 36'sb110010110000110111100110010110000101;
            sine_reg0   <= 36'sb11101001000100101010111000110111001;
        end
        1303: begin
            cosine_reg0 <= 36'sb110010101110000000100110111010000010;
            sine_reg0   <= 36'sb11101000111010010000011011100001111;
        end
        1304: begin
            cosine_reg0 <= 36'sb110010101011001001101111101010010011;
            sine_reg0   <= 36'sb11101000101111110011101110100001111;
        end
        1305: begin
            cosine_reg0 <= 36'sb110010101000010011000000101000101001;
            sine_reg0   <= 36'sb11101000100101010100110001111101010;
        end
        1306: begin
            cosine_reg0 <= 36'sb110010100101011100011001110110110101;
            sine_reg0   <= 36'sb11101000011010110011100101111010110;
        end
        1307: begin
            cosine_reg0 <= 36'sb110010100010100101111011010110100111;
            sine_reg0   <= 36'sb11101000010000010000001010100000101;
        end
        1308: begin
            cosine_reg0 <= 36'sb110010011111101111100101001001110001;
            sine_reg0   <= 36'sb11101000000101101010011111110101100;
        end
        1309: begin
            cosine_reg0 <= 36'sb110010011100111001010111010010000001;
            sine_reg0   <= 36'sb11100111111011000010100101111111111;
        end
        1310: begin
            cosine_reg0 <= 36'sb110010011010000011010001110001001010;
            sine_reg0   <= 36'sb11100111110000011000011101000110011;
        end
        1311: begin
            cosine_reg0 <= 36'sb110010010111001101010100101000111011;
            sine_reg0   <= 36'sb11100111100101101100000101001111100;
        end
        1312: begin
            cosine_reg0 <= 36'sb110010010100010111011111111011000100;
            sine_reg0   <= 36'sb11100111011010111101011110100001110;
        end
        1313: begin
            cosine_reg0 <= 36'sb110010010001100001110011101001010110;
            sine_reg0   <= 36'sb11100111010000001100101001000100000;
        end
        1314: begin
            cosine_reg0 <= 36'sb110010001110101100001111110101100001;
            sine_reg0   <= 36'sb11100111000101011001100100111100110;
        end
        1315: begin
            cosine_reg0 <= 36'sb110010001011110110110100100001010100;
            sine_reg0   <= 36'sb11100110111010100100010010010010100;
        end
        1316: begin
            cosine_reg0 <= 36'sb110010001001000001100001101110100000;
            sine_reg0   <= 36'sb11100110101111101100110001001100010;
        end
        1317: begin
            cosine_reg0 <= 36'sb110010000110001100010111011110110100;
            sine_reg0   <= 36'sb11100110100100110011000001110000100;
        end
        1318: begin
            cosine_reg0 <= 36'sb110010000011010111010101110100000000;
            sine_reg0   <= 36'sb11100110011001110111000100000110000;
        end
        1319: begin
            cosine_reg0 <= 36'sb110010000000100010011100101111110101;
            sine_reg0   <= 36'sb11100110001110111000111000010011100;
        end
        1320: begin
            cosine_reg0 <= 36'sb110001111101101101101100010100000000;
            sine_reg0   <= 36'sb11100110000011111000011110011111110;
        end
        1321: begin
            cosine_reg0 <= 36'sb110001111010111001000100100010010011;
            sine_reg0   <= 36'sb11100101111000110101110110110001101;
        end
        1322: begin
            cosine_reg0 <= 36'sb110001111000000100100101011100011100;
            sine_reg0   <= 36'sb11100101101101110001000001001111111;
        end
        1323: begin
            cosine_reg0 <= 36'sb110001110101010000001111000100001010;
            sine_reg0   <= 36'sb11100101100010101001111110000001011;
        end
        1324: begin
            cosine_reg0 <= 36'sb110001110010011100000001011011001110;
            sine_reg0   <= 36'sb11100101010111100000101101001100111;
        end
        1325: begin
            cosine_reg0 <= 36'sb110001101111100111111100100011010101;
            sine_reg0   <= 36'sb11100101001100010101001110111001011;
        end
        1326: begin
            cosine_reg0 <= 36'sb110001101100110100000000011110010000;
            sine_reg0   <= 36'sb11100101000001000111100011001101110;
        end
        1327: begin
            cosine_reg0 <= 36'sb110001101010000000001101001101101100;
            sine_reg0   <= 36'sb11100100110101110111101010010000110;
        end
        1328: begin
            cosine_reg0 <= 36'sb110001100111001100100010110011011010;
            sine_reg0   <= 36'sb11100100101010100101100100001001100;
        end
        1329: begin
            cosine_reg0 <= 36'sb110001100100011001000001010001001000;
            sine_reg0   <= 36'sb11100100011111010001010000111110111;
        end
        1330: begin
            cosine_reg0 <= 36'sb110001100001100101101000101000100100;
            sine_reg0   <= 36'sb11100100010011111010110000111000000;
        end
        1331: begin
            cosine_reg0 <= 36'sb110001011110110010011000111011011110;
            sine_reg0   <= 36'sb11100100001000100010000011111011101;
        end
        1332: begin
            cosine_reg0 <= 36'sb110001011011111111010010001011100011;
            sine_reg0   <= 36'sb11100011111101000111001010010001000;
        end
        1333: begin
            cosine_reg0 <= 36'sb110001011001001100010100011010100011;
            sine_reg0   <= 36'sb11100011110001101010000011111111000;
        end
        1334: begin
            cosine_reg0 <= 36'sb110001010110011001011111101010001011;
            sine_reg0   <= 36'sb11100011100110001010110001001100111;
        end
        1335: begin
            cosine_reg0 <= 36'sb110001010011100110110011111100001011;
            sine_reg0   <= 36'sb11100011011010101001010010000001100;
        end
        1336: begin
            cosine_reg0 <= 36'sb110001010000110100010001010010010000;
            sine_reg0   <= 36'sb11100011001111000101100110100100001;
        end
        1337: begin
            cosine_reg0 <= 36'sb110001001110000001110111101110001000;
            sine_reg0   <= 36'sb11100011000011011111101110111011111;
        end
        1338: begin
            cosine_reg0 <= 36'sb110001001011001111100111010001100001;
            sine_reg0   <= 36'sb11100010110111110111101011001111111;
        end
        1339: begin
            cosine_reg0 <= 36'sb110001001000011101011111111110001010;
            sine_reg0   <= 36'sb11100010101100001101011011100111010;
        end
        1340: begin
            cosine_reg0 <= 36'sb110001000101101011100001110101110000;
            sine_reg0   <= 36'sb11100010100000100001000000001001010;
        end
        1341: begin
            cosine_reg0 <= 36'sb110001000010111001101100111010000001;
            sine_reg0   <= 36'sb11100010010100110010011000111101001;
        end
        1342: begin
            cosine_reg0 <= 36'sb110001000000001000000001001100101011;
            sine_reg0   <= 36'sb11100010001001000001100110001010000;
        end
        1343: begin
            cosine_reg0 <= 36'sb110000111101010110011110101111011100;
            sine_reg0   <= 36'sb11100001111101001110100111110111001;
        end
        1344: begin
            cosine_reg0 <= 36'sb110000111010100101000101100100000000;
            sine_reg0   <= 36'sb11100001110001011001011110001011111;
        end
        1345: begin
            cosine_reg0 <= 36'sb110000110111110011110101101100000101;
            sine_reg0   <= 36'sb11100001100101100010001001001111101;
        end
        1346: begin
            cosine_reg0 <= 36'sb110000110101000010101111001001011001;
            sine_reg0   <= 36'sb11100001011001101000101001001001100;
        end
        1347: begin
            cosine_reg0 <= 36'sb110000110010010001110001111101101001;
            sine_reg0   <= 36'sb11100001001101101100111110000000111;
        end
        1348: begin
            cosine_reg0 <= 36'sb110000101111100000111110001010100001;
            sine_reg0   <= 36'sb11100001000001101111000111111101001;
        end
        1349: begin
            cosine_reg0 <= 36'sb110000101100110000010011110001110000;
            sine_reg0   <= 36'sb11100000110101101111000111000101110;
        end
        1350: begin
            cosine_reg0 <= 36'sb110000101001111111110010110101000010;
            sine_reg0   <= 36'sb11100000101001101100111011100010001;
        end
        1351: begin
            cosine_reg0 <= 36'sb110000100111001111011011010110000100;
            sine_reg0   <= 36'sb11100000011101101000100101011001100;
        end
        1352: begin
            cosine_reg0 <= 36'sb110000100100011111001101010110100011;
            sine_reg0   <= 36'sb11100000010001100010000100110011100;
        end
        1353: begin
            cosine_reg0 <= 36'sb110000100001101111001000111000001011;
            sine_reg0   <= 36'sb11100000000101011001011001110111100;
        end
        1354: begin
            cosine_reg0 <= 36'sb110000011110111111001101111100101000;
            sine_reg0   <= 36'sb11011111111001001110100100101101000;
        end
        1355: begin
            cosine_reg0 <= 36'sb110000011100001111011100100101101001;
            sine_reg0   <= 36'sb11011111101101000001100101011011100;
        end
        1356: begin
            cosine_reg0 <= 36'sb110000011001011111110100110100111001;
            sine_reg0   <= 36'sb11011111100000110010011100001010100;
        end
        1357: begin
            cosine_reg0 <= 36'sb110000010110110000010110101100000011;
            sine_reg0   <= 36'sb11011111010100100001001001000001101;
        end
        1358: begin
            cosine_reg0 <= 36'sb110000010100000001000010001100110110;
            sine_reg0   <= 36'sb11011111001000001101101100001000011;
        end
        1359: begin
            cosine_reg0 <= 36'sb110000010001010001110111011000111100;
            sine_reg0   <= 36'sb11011110111011111000000101100110100;
        end
        1360: begin
            cosine_reg0 <= 36'sb110000001110100010110110010010000001;
            sine_reg0   <= 36'sb11011110101111100000010101100011011;
        end
        1361: begin
            cosine_reg0 <= 36'sb110000001011110011111110111001110011;
            sine_reg0   <= 36'sb11011110100011000110011100000110110;
        end
        1362: begin
            cosine_reg0 <= 36'sb110000001001000101010001010001111100;
            sine_reg0   <= 36'sb11011110010110101010011001011000010;
        end
        1363: begin
            cosine_reg0 <= 36'sb110000000110010110101101011100001000;
            sine_reg0   <= 36'sb11011110001010001100001101011111101;
        end
        1364: begin
            cosine_reg0 <= 36'sb110000000011101000010011011010000100;
            sine_reg0   <= 36'sb11011101111101101011111000100100100;
        end
        1365: begin
            cosine_reg0 <= 36'sb110000000000111010000011001101011010;
            sine_reg0   <= 36'sb11011101110001001001011010101110101;
        end
        1366: begin
            cosine_reg0 <= 36'sb101111111110001011111100110111110110;
            sine_reg0   <= 36'sb11011101100100100100110100000101101;
        end
        1367: begin
            cosine_reg0 <= 36'sb101111111011011110000000011011000011;
            sine_reg0   <= 36'sb11011101010111111110000100110001011;
        end
        1368: begin
            cosine_reg0 <= 36'sb101111111000110000001101111000101101;
            sine_reg0   <= 36'sb11011101001011010101001100111001101;
        end
        1369: begin
            cosine_reg0 <= 36'sb101111110110000010100101010010100000;
            sine_reg0   <= 36'sb11011100111110101010001100100110001;
        end
        1370: begin
            cosine_reg0 <= 36'sb101111110011010101000110101010000101;
            sine_reg0   <= 36'sb11011100110001111101000011111110101;
        end
        1371: begin
            cosine_reg0 <= 36'sb101111110000100111110010000001001001;
            sine_reg0   <= 36'sb11011100100101001101110011001011010;
        end
        1372: begin
            cosine_reg0 <= 36'sb101111101101111010100111011001010101;
            sine_reg0   <= 36'sb11011100011000011100011010010011100;
        end
        1373: begin
            cosine_reg0 <= 36'sb101111101011001101100110110100010101;
            sine_reg0   <= 36'sb11011100001011101000111001011111100;
        end
        1374: begin
            cosine_reg0 <= 36'sb101111101000100000110000010011110100;
            sine_reg0   <= 36'sb11011011111110110011010000110111001;
        end
        1375: begin
            cosine_reg0 <= 36'sb101111100101110100000011111001011100;
            sine_reg0   <= 36'sb11011011110001111011100000100010010;
        end
        1376: begin
            cosine_reg0 <= 36'sb101111100011000111100001100110111000;
            sine_reg0   <= 36'sb11011011100101000001101000101000101;
        end
        1377: begin
            cosine_reg0 <= 36'sb101111100000011011001001011101110010;
            sine_reg0   <= 36'sb11011011011000000101101001010010101;
        end
        1378: begin
            cosine_reg0 <= 36'sb101111011101101110111011011111110100;
            sine_reg0   <= 36'sb11011011001011000111100010100111111;
        end
        1379: begin
            cosine_reg0 <= 36'sb101111011011000010110111101110101001;
            sine_reg0   <= 36'sb11011010111110000111010100110000100;
        end
        1380: begin
            cosine_reg0 <= 36'sb101111011000010110111110001011111011;
            sine_reg0   <= 36'sb11011010110001000100111111110100100;
        end
        1381: begin
            cosine_reg0 <= 36'sb101111010101101011001110111001010011;
            sine_reg0   <= 36'sb11011010100100000000100011111011111;
        end
        1382: begin
            cosine_reg0 <= 36'sb101111010010111111101001111000011101;
            sine_reg0   <= 36'sb11011010010110111010000001001110111;
        end
        1383: begin
            cosine_reg0 <= 36'sb101111010000010100001111001011000001;
            sine_reg0   <= 36'sb11011010001001110001010111110101011;
        end
        1384: begin
            cosine_reg0 <= 36'sb101111001101101000111110110010101001;
            sine_reg0   <= 36'sb11011001111100100110100111110111100;
        end
        1385: begin
            cosine_reg0 <= 36'sb101111001010111101111000110001000000;
            sine_reg0   <= 36'sb11011001101111011001110001011101100;
        end
        1386: begin
            cosine_reg0 <= 36'sb101111001000010010111101000111101110;
            sine_reg0   <= 36'sb11011001100010001010110100101111100;
        end
        1387: begin
            cosine_reg0 <= 36'sb101111000101101000001011111000011101;
            sine_reg0   <= 36'sb11011001010100111001110001110101100;
        end
        1388: begin
            cosine_reg0 <= 36'sb101111000010111101100101000100110110;
            sine_reg0   <= 36'sb11011001000111100110101000110111111;
        end
        1389: begin
            cosine_reg0 <= 36'sb101111000000010011001000101110100011;
            sine_reg0   <= 36'sb11011000111010010001011001111110110;
        end
        1390: begin
            cosine_reg0 <= 36'sb101110111101101000110110110111001100;
            sine_reg0   <= 36'sb11011000101100111010000101010010010;
        end
        1391: begin
            cosine_reg0 <= 36'sb101110111010111110101111100000011100;
            sine_reg0   <= 36'sb11011000011111100000101010111010110;
        end
        1392: begin
            cosine_reg0 <= 36'sb101110111000010100110010101011111010;
            sine_reg0   <= 36'sb11011000010010000101001011000000100;
        end
        1393: begin
            cosine_reg0 <= 36'sb101110110101101011000000011011001111;
            sine_reg0   <= 36'sb11011000000100100111100101101011110;
        end
        1394: begin
            cosine_reg0 <= 36'sb101110110011000001011000110000000101;
            sine_reg0   <= 36'sb11010111110111000111111011000100111;
        end
        1395: begin
            cosine_reg0 <= 36'sb101110110000010111111011101100000100;
            sine_reg0   <= 36'sb11010111101001100110001011010100001;
        end
        1396: begin
            cosine_reg0 <= 36'sb101110101101101110101001010000110100;
            sine_reg0   <= 36'sb11010111011100000010010110100001110;
        end
        1397: begin
            cosine_reg0 <= 36'sb101110101011000101100001011111111110;
            sine_reg0   <= 36'sb11010111001110011100011100110110010;
        end
        1398: begin
            cosine_reg0 <= 36'sb101110101000011100100100011011001010;
            sine_reg0   <= 36'sb11010111000000110100011110011010001;
        end
        1399: begin
            cosine_reg0 <= 36'sb101110100101110011110010000100000000;
            sine_reg0   <= 36'sb11010110110011001010011011010101100;
        end
        1400: begin
            cosine_reg0 <= 36'sb101110100011001011001010011100001001;
            sine_reg0   <= 36'sb11010110100101011110010011110001000;
        end
        1401: begin
            cosine_reg0 <= 36'sb101110100000100010101101100101001100;
            sine_reg0   <= 36'sb11010110010111110000000111110100111;
        end
        1402: begin
            cosine_reg0 <= 36'sb101110011101111010011011100000110010;
            sine_reg0   <= 36'sb11010110001001111111110111101001111;
        end
        1403: begin
            cosine_reg0 <= 36'sb101110011011010010010100010000100010;
            sine_reg0   <= 36'sb11010101111100001101100011011000010;
        end
        1404: begin
            cosine_reg0 <= 36'sb101110011000101010010111110110000100;
            sine_reg0   <= 36'sb11010101101110011001001011001000101;
        end
        1405: begin
            cosine_reg0 <= 36'sb101110010110000010100110010010111111;
            sine_reg0   <= 36'sb11010101100000100010101111000011100;
        end
        1406: begin
            cosine_reg0 <= 36'sb101110010011011010111111101000111100;
            sine_reg0   <= 36'sb11010101010010101010001111010001010;
        end
        1407: begin
            cosine_reg0 <= 36'sb101110010000110011100011111001100000;
            sine_reg0   <= 36'sb11010101000100101111101011111010110;
        end
        1408: begin
            cosine_reg0 <= 36'sb101110001110001100010011000110010101;
            sine_reg0   <= 36'sb11010100110110110011000101001000011;
        end
        1409: begin
            cosine_reg0 <= 36'sb101110001011100101001101010001000000;
            sine_reg0   <= 36'sb11010100101000110100011011000010110;
        end
        1410: begin
            cosine_reg0 <= 36'sb101110001000111110010010011011001001;
            sine_reg0   <= 36'sb11010100011010110011101101110010100;
        end
        1411: begin
            cosine_reg0 <= 36'sb101110000110010111100010100110011000;
            sine_reg0   <= 36'sb11010100001100110000111101100000011;
        end
        1412: begin
            cosine_reg0 <= 36'sb101110000011110000111101110100010001;
            sine_reg0   <= 36'sb11010011111110101100001010010100111;
        end
        1413: begin
            cosine_reg0 <= 36'sb101110000001001010100100000110011110;
            sine_reg0   <= 36'sb11010011110000100101010100011000110;
        end
        1414: begin
            cosine_reg0 <= 36'sb101101111110100100010101011110100011;
            sine_reg0   <= 36'sb11010011100010011100011011110100111;
        end
        1415: begin
            cosine_reg0 <= 36'sb101101111011111110010001111110001000;
            sine_reg0   <= 36'sb11010011010100010001100000110001101;
        end
        1416: begin
            cosine_reg0 <= 36'sb101101111001011000011001100110110100;
            sine_reg0   <= 36'sb11010011000110000100100011011000000;
        end
        1417: begin
            cosine_reg0 <= 36'sb101101110110110010101100011010001011;
            sine_reg0   <= 36'sb11010010110111110101100011110000101;
        end
        1418: begin
            cosine_reg0 <= 36'sb101101110100001101001010011001110110;
            sine_reg0   <= 36'sb11010010101001100100100010000100011;
        end
        1419: begin
            cosine_reg0 <= 36'sb101101110001100111110011100111011001;
            sine_reg0   <= 36'sb11010010011011010001011110011100001;
        end
        1420: begin
            cosine_reg0 <= 36'sb101101101111000010101000000100011010;
            sine_reg0   <= 36'sb11010010001100111100011001000000100;
        end
        1421: begin
            cosine_reg0 <= 36'sb101101101100011101100111110010100001;
            sine_reg0   <= 36'sb11010001111110100101010001111010011;
        end
        1422: begin
            cosine_reg0 <= 36'sb101101101001111000110010110011010010;
            sine_reg0   <= 36'sb11010001110000001100001001010010101;
        end
        1423: begin
            cosine_reg0 <= 36'sb101101100111010100001001001000010011;
            sine_reg0   <= 36'sb11010001100001110000111111010010010;
        end
        1424: begin
            cosine_reg0 <= 36'sb101101100100101111101010110011001001;
            sine_reg0   <= 36'sb11010001010011010011110100000010001;
        end
        1425: begin
            cosine_reg0 <= 36'sb101101100010001011010111110101011011;
            sine_reg0   <= 36'sb11010001000100110100100111101011000;
        end
        1426: begin
            cosine_reg0 <= 36'sb101101011111100111010000010000101101;
            sine_reg0   <= 36'sb11010000110110010011011010010101111;
        end
        1427: begin
            cosine_reg0 <= 36'sb101101011101000011010100000110100101;
            sine_reg0   <= 36'sb11010000100111110000001100001011111;
        end
        1428: begin
            cosine_reg0 <= 36'sb101101011010011111100011011000101000;
            sine_reg0   <= 36'sb11010000011001001010111101010101110;
        end
        1429: begin
            cosine_reg0 <= 36'sb101101010111111011111110001000011011;
            sine_reg0   <= 36'sb11010000001010100011101101111100101;
        end
        1430: begin
            cosine_reg0 <= 36'sb101101010101011000100100010111100010;
            sine_reg0   <= 36'sb11001111111011111010011110001001100;
        end
        1431: begin
            cosine_reg0 <= 36'sb101101010010110101010110000111100011;
            sine_reg0   <= 36'sb11001111101101001111001110000101010;
        end
        1432: begin
            cosine_reg0 <= 36'sb101101010000010010010011011010000010;
            sine_reg0   <= 36'sb11001111011110100001111101111001010;
        end
        1433: begin
            cosine_reg0 <= 36'sb101101001101101111011100010000100100;
            sine_reg0   <= 36'sb11001111001111110010101101101110010;
        end
        1434: begin
            cosine_reg0 <= 36'sb101101001011001100110000101100101101;
            sine_reg0   <= 36'sb11001111000001000001011101101101100;
        end
        1435: begin
            cosine_reg0 <= 36'sb101101001000101010010000110000000010;
            sine_reg0   <= 36'sb11001110110010001110001110000000001;
        end
        1436: begin
            cosine_reg0 <= 36'sb101101000110000111111100011100000110;
            sine_reg0   <= 36'sb11001110100011011000111110101111010;
        end
        1437: begin
            cosine_reg0 <= 36'sb101101000011100101110011110010011111;
            sine_reg0   <= 36'sb11001110010100100001110000000011111;
        end
        1438: begin
            cosine_reg0 <= 36'sb101101000001000011110110110100110000;
            sine_reg0   <= 36'sb11001110000101101000100010000111011;
        end
        1439: begin
            cosine_reg0 <= 36'sb101100111110100010000101100100011100;
            sine_reg0   <= 36'sb11001101110110101101010101000010111;
        end
        1440: begin
            cosine_reg0 <= 36'sb101100111100000000100000000011001000;
            sine_reg0   <= 36'sb11001101100111110000001000111111100;
        end
        1441: begin
            cosine_reg0 <= 36'sb101100111001011111000110010010011000;
            sine_reg0   <= 36'sb11001101011000110000111110000110100;
        end
        1442: begin
            cosine_reg0 <= 36'sb101100110110111101111000010011101110;
            sine_reg0   <= 36'sb11001101001001101111110100100001010;
        end
        1443: begin
            cosine_reg0 <= 36'sb101100110100011100110110001000101111;
            sine_reg0   <= 36'sb11001100111010101100101100011000111;
        end
        1444: begin
            cosine_reg0 <= 36'sb101100110001111011111111110010111101;
            sine_reg0   <= 36'sb11001100101011100111100101110110101;
        end
        1445: begin
            cosine_reg0 <= 36'sb101100101111011011010101010011111101;
            sine_reg0   <= 36'sb11001100011100100000100001000100000;
        end
        1446: begin
            cosine_reg0 <= 36'sb101100101100111010110110101101010000;
            sine_reg0   <= 36'sb11001100001101010111011110001010001;
        end
        1447: begin
            cosine_reg0 <= 36'sb101100101010011010100100000000011011;
            sine_reg0   <= 36'sb11001011111110001100011101010010011;
        end
        1448: begin
            cosine_reg0 <= 36'sb101100100111111010011101001110111111;
            sine_reg0   <= 36'sb11001011101110111111011110100110001;
        end
        1449: begin
            cosine_reg0 <= 36'sb101100100101011010100010011010100000;
            sine_reg0   <= 36'sb11001011011111110000100010001110111;
        end
        1450: begin
            cosine_reg0 <= 36'sb101100100010111010110011100100100000;
            sine_reg0   <= 36'sb11001011010000011111101000010101111;
        end
        1451: begin
            cosine_reg0 <= 36'sb101100100000011011010000101110100010;
            sine_reg0   <= 36'sb11001011000001001100110001000100100;
        end
        1452: begin
            cosine_reg0 <= 36'sb101100011101111011111001111010001001;
            sine_reg0   <= 36'sb11001010110001110111111100100100011;
        end
        1453: begin
            cosine_reg0 <= 36'sb101100011011011100101111001000110101;
            sine_reg0   <= 36'sb11001010100010100001001010111110110;
        end
        1454: begin
            cosine_reg0 <= 36'sb101100011000111101110000011100001011;
            sine_reg0   <= 36'sb11001010010011001000011100011101010;
        end
        1455: begin
            cosine_reg0 <= 36'sb101100010110011110111101110101101011;
            sine_reg0   <= 36'sb11001010000011101101110001001001011;
        end
        1456: begin
            cosine_reg0 <= 36'sb101100010100000000010111010110111001;
            sine_reg0   <= 36'sb11001001110100010001001001001100100;
        end
        1457: begin
            cosine_reg0 <= 36'sb101100010001100001111101000001010100;
            sine_reg0   <= 36'sb11001001100100110010100100110000010;
        end
        1458: begin
            cosine_reg0 <= 36'sb101100001111000011101110110110100000;
            sine_reg0   <= 36'sb11001001010101010010000011111110001;
        end
        1459: begin
            cosine_reg0 <= 36'sb101100001100100101101100110111111110;
            sine_reg0   <= 36'sb11001001000101101111100110111111101;
        end
        1460: begin
            cosine_reg0 <= 36'sb101100001010000111110111000111001111;
            sine_reg0   <= 36'sb11001000110110001011001101111110100;
        end
        1461: begin
            cosine_reg0 <= 36'sb101100000111101010001101100101110101;
            sine_reg0   <= 36'sb11001000100110100100111001000100011;
        end
        1462: begin
            cosine_reg0 <= 36'sb101100000101001100110000010101010001;
            sine_reg0   <= 36'sb11001000010110111100101000011010101;
        end
        1463: begin
            cosine_reg0 <= 36'sb101100000010101111011111010111000100;
            sine_reg0   <= 36'sb11001000000111010010011100001011001;
        end
        1464: begin
            cosine_reg0 <= 36'sb101100000000010010011010101100101111;
            sine_reg0   <= 36'sb11000111110111100110010100011111011;
        end
        1465: begin
            cosine_reg0 <= 36'sb101011111101110101100010010111110011;
            sine_reg0   <= 36'sb11000111100111111000010001100001001;
        end
        1466: begin
            cosine_reg0 <= 36'sb101011111011011000110110011001110001;
            sine_reg0   <= 36'sb11000111011000001000010011011010001;
        end
        1467: begin
            cosine_reg0 <= 36'sb101011111000111100010110110100001010;
            sine_reg0   <= 36'sb11000111001000010110011010010100001;
        end
        1468: begin
            cosine_reg0 <= 36'sb101011110110100000000011101000011101;
            sine_reg0   <= 36'sb11000110111000100010100110011000101;
        end
        1469: begin
            cosine_reg0 <= 36'sb101011110100000011111100111000001100;
            sine_reg0   <= 36'sb11000110101000101100110111110001100;
        end
        1470: begin
            cosine_reg0 <= 36'sb101011110001101000000010100100110110;
            sine_reg0   <= 36'sb11000110011000110101001110101000101;
        end
        1471: begin
            cosine_reg0 <= 36'sb101011101111001100010100101111111100;
            sine_reg0   <= 36'sb11000110001000111011101011000111110;
        end
        1472: begin
            cosine_reg0 <= 36'sb101011101100110000110011011010111110;
            sine_reg0   <= 36'sb11000101111001000000001101011000100;
        end
        1473: begin
            cosine_reg0 <= 36'sb101011101010010101011110100111011100;
            sine_reg0   <= 36'sb11000101101001000010110101100101000;
        end
        1474: begin
            cosine_reg0 <= 36'sb101011100111111010010110010110110110;
            sine_reg0   <= 36'sb11000101011001000011100011110110111;
        end
        1475: begin
            cosine_reg0 <= 36'sb101011100101011111011010101010101011;
            sine_reg0   <= 36'sb11000101001001000010011000011000000;
        end
        1476: begin
            cosine_reg0 <= 36'sb101011100011000100101011100100011011;
            sine_reg0   <= 36'sb11000100111000111111010011010010011;
        end
        1477: begin
            cosine_reg0 <= 36'sb101011100000101010001001000101100101;
            sine_reg0   <= 36'sb11000100101000111010010100101111110;
        end
        1478: begin
            cosine_reg0 <= 36'sb101011011110001111110011001111101000;
            sine_reg0   <= 36'sb11000100011000110011011100111010001;
        end
        1479: begin
            cosine_reg0 <= 36'sb101011011011110101101010000100000101;
            sine_reg0   <= 36'sb11000100001000101010101011111011100;
        end
        1480: begin
            cosine_reg0 <= 36'sb101011011001011011101101100100011010;
            sine_reg0   <= 36'sb11000011111000100000000001111101110;
        end
        1481: begin
            cosine_reg0 <= 36'sb101011010111000001111101110010000101;
            sine_reg0   <= 36'sb11000011101000010011011111001010110;
        end
        1482: begin
            cosine_reg0 <= 36'sb101011010100101000011010101110100111;
            sine_reg0   <= 36'sb11000011011000000101000011101100110;
        end
        1483: begin
            cosine_reg0 <= 36'sb101011010010001111000100011011011101;
            sine_reg0   <= 36'sb11000011000111110100101111101101100;
        end
        1484: begin
            cosine_reg0 <= 36'sb101011001111110101111010111010000110;
            sine_reg0   <= 36'sb11000010110111100010100011010111010;
        end
        1485: begin
            cosine_reg0 <= 36'sb101011001101011100111110001100000000;
            sine_reg0   <= 36'sb11000010100111001110011110110011110;
        end
        1486: begin
            cosine_reg0 <= 36'sb101011001011000100001110010010101010;
            sine_reg0   <= 36'sb11000010010110111000100010001101011;
        end
        1487: begin
            cosine_reg0 <= 36'sb101011001000101011101011001111100011;
            sine_reg0   <= 36'sb11000010000110100000101101101110000;
        end
        1488: begin
            cosine_reg0 <= 36'sb101011000110010011010101000100001000;
            sine_reg0   <= 36'sb11000001110110000111000001011111111;
        end
        1489: begin
            cosine_reg0 <= 36'sb101011000011111011001011110001110111;
            sine_reg0   <= 36'sb11000001100101101011011101101101000;
        end
        1490: begin
            cosine_reg0 <= 36'sb101011000001100011001111011010001101;
            sine_reg0   <= 36'sb11000001010101001110000010011111101;
        end
        1491: begin
            cosine_reg0 <= 36'sb101010111111001011011111111110101010;
            sine_reg0   <= 36'sb11000001000100101110110000000001110;
        end
        1492: begin
            cosine_reg0 <= 36'sb101010111100110011111101100000101010;
            sine_reg0   <= 36'sb11000000110100001101100110011101101;
        end
        1493: begin
            cosine_reg0 <= 36'sb101010111010011100101000000001101011;
            sine_reg0   <= 36'sb11000000100011101010100101111101011;
        end
        1494: begin
            cosine_reg0 <= 36'sb101010111000000101011111100011001010;
            sine_reg0   <= 36'sb11000000010011000101101110101011011;
        end
        1495: begin
            cosine_reg0 <= 36'sb101010110101101110100100000110100101;
            sine_reg0   <= 36'sb11000000000010011111000000110001101;
        end
        1496: begin
            cosine_reg0 <= 36'sb101010110011010111110101101101011000;
            sine_reg0   <= 36'sb10111111110001110110011100011010101;
        end
        1497: begin
            cosine_reg0 <= 36'sb101010110001000001010100011001000000;
            sine_reg0   <= 36'sb10111111100001001100000001110000100;
        end
        1498: begin
            cosine_reg0 <= 36'sb101010101110101011000000001010111011;
            sine_reg0   <= 36'sb10111111010000011111110000111101011;
        end
        1499: begin
            cosine_reg0 <= 36'sb101010101100010100111001000100100101;
            sine_reg0   <= 36'sb10111110111111110001101010001011111;
        end
        1500: begin
            cosine_reg0 <= 36'sb101010101001111110111111000111011011;
            sine_reg0   <= 36'sb10111110101111000001101101100110000;
        end
        1501: begin
            cosine_reg0 <= 36'sb101010100111101001010010010100111001;
            sine_reg0   <= 36'sb10111110011110001111111011010110010;
        end
        1502: begin
            cosine_reg0 <= 36'sb101010100101010011110010101110011011;
            sine_reg0   <= 36'sb10111110001101011100010011100111000;
        end
        1503: begin
            cosine_reg0 <= 36'sb101010100010111110100000010101011110;
            sine_reg0   <= 36'sb10111101111100100110110110100010100;
        end
        1504: begin
            cosine_reg0 <= 36'sb101010100000101001011011001011011101;
            sine_reg0   <= 36'sb10111101101011101111100100010011010;
        end
        1505: begin
            cosine_reg0 <= 36'sb101010011110010100100011010001110110;
            sine_reg0   <= 36'sb10111101011010110110011101000011100;
        end
        1506: begin
            cosine_reg0 <= 36'sb101010011011111111111000101010000011;
            sine_reg0   <= 36'sb10111101001001111011100000111101111;
        end
        1507: begin
            cosine_reg0 <= 36'sb101010011001101011011011010101100000;
            sine_reg0   <= 36'sb10111100111000111110110000001100101;
        end
        1508: begin
            cosine_reg0 <= 36'sb101010010111010111001011010101101001;
            sine_reg0   <= 36'sb10111100101000000000001010111010011;
        end
        1509: begin
            cosine_reg0 <= 36'sb101010010101000011001000101011111010;
            sine_reg0   <= 36'sb10111100010110111111110001010001100;
        end
        1510: begin
            cosine_reg0 <= 36'sb101010010010101111010011011001101101;
            sine_reg0   <= 36'sb10111100000101111101100011011100011;
        end
        1511: begin
            cosine_reg0 <= 36'sb101010010000011011101011100000011110;
            sine_reg0   <= 36'sb10111011110100111001100001100101110;
        end
        1512: begin
            cosine_reg0 <= 36'sb101010001110001000010001000001100111;
            sine_reg0   <= 36'sb10111011100011110011101011111000000;
        end
        1513: begin
            cosine_reg0 <= 36'sb101010001011110101000011111110100101;
            sine_reg0   <= 36'sb10111011010010101100000010011101110;
        end
        1514: begin
            cosine_reg0 <= 36'sb101010001001100010000100011000110001;
            sine_reg0   <= 36'sb10111011000001100010100101100001011;
        end
        1515: begin
            cosine_reg0 <= 36'sb101010000111001111010010010001100111;
            sine_reg0   <= 36'sb10111010110000010111010101001101110;
        end
        1516: begin
            cosine_reg0 <= 36'sb101010000100111100101101101010100000;
            sine_reg0   <= 36'sb10111010011111001010010001101101001;
        end
        1517: begin
            cosine_reg0 <= 36'sb101010000010101010010110100100110111;
            sine_reg0   <= 36'sb10111010001101111011011011001010100;
        end
        1518: begin
            cosine_reg0 <= 36'sb101010000000011000001101000010000111;
            sine_reg0   <= 36'sb10111001111100101010110001110000001;
        end
        1519: begin
            cosine_reg0 <= 36'sb101001111110000110010001000011101010;
            sine_reg0   <= 36'sb10111001101011011000010101101000111;
        end
        1520: begin
            cosine_reg0 <= 36'sb101001111011110100100010101010111001;
            sine_reg0   <= 36'sb10111001011010000100000110111111011;
        end
        1521: begin
            cosine_reg0 <= 36'sb101001111001100011000001111001001111;
            sine_reg0   <= 36'sb10111001001000101110000101111110011;
        end
        1522: begin
            cosine_reg0 <= 36'sb101001110111010001101110110000000110;
            sine_reg0   <= 36'sb10111000110111010110010010110000011;
        end
        1523: begin
            cosine_reg0 <= 36'sb101001110101000000101001010000110110;
            sine_reg0   <= 36'sb10111000100101111100101101100000010;
        end
        1524: begin
            cosine_reg0 <= 36'sb101001110010101111110001011100111010;
            sine_reg0   <= 36'sb10111000010100100001010110011000101;
        end
        1525: begin
            cosine_reg0 <= 36'sb101001110000011111000111010101101010;
            sine_reg0   <= 36'sb10111000000011000100001101100100011;
        end
        1526: begin
            cosine_reg0 <= 36'sb101001101110001110101010111100100001;
            sine_reg0   <= 36'sb10110111110001100101010011001110010;
        end
        1527: begin
            cosine_reg0 <= 36'sb101001101011111110011100010010110111;
            sine_reg0   <= 36'sb10110111100000000100100111100000111;
        end
        1528: begin
            cosine_reg0 <= 36'sb101001101001101110011011011010000101;
            sine_reg0   <= 36'sb10110111001110100010001010100111010;
        end
        1529: begin
            cosine_reg0 <= 36'sb101001100111011110101000010011100011;
            sine_reg0   <= 36'sb10110110111100111101111100101100001;
        end
        1530: begin
            cosine_reg0 <= 36'sb101001100101001111000011000000101100;
            sine_reg0   <= 36'sb10110110101011010111111101111010010;
        end
        1531: begin
            cosine_reg0 <= 36'sb101001100010111111101011100010110111;
            sine_reg0   <= 36'sb10110110011001110000001110011100101;
        end
        1532: begin
            cosine_reg0 <= 36'sb101001100000110000100001111011011100;
            sine_reg0   <= 36'sb10110110001000000110101110011110000;
        end
        1533: begin
            cosine_reg0 <= 36'sb101001011110100001100110001011110101;
            sine_reg0   <= 36'sb10110101110110011011011110001001010;
        end
        1534: begin
            cosine_reg0 <= 36'sb101001011100010010111000010101011000;
            sine_reg0   <= 36'sb10110101100100101110011101101001011;
        end
        1535: begin
            cosine_reg0 <= 36'sb101001011010000100011000011001011111;
            sine_reg0   <= 36'sb10110101010010111111101101001001010;
        end
        1536: begin
            cosine_reg0 <= 36'sb101001010111110110000110011001100001;
            sine_reg0   <= 36'sb10110101000001001111001100110011111;
        end
        1537: begin
            cosine_reg0 <= 36'sb101001010101101000000010010110110110;
            sine_reg0   <= 36'sb10110100101111011100111100110100001;
        end
        1538: begin
            cosine_reg0 <= 36'sb101001010011011010001100010010110101;
            sine_reg0   <= 36'sb10110100011101101000111101010101000;
        end
        1539: begin
            cosine_reg0 <= 36'sb101001010001001100100100001110110110;
            sine_reg0   <= 36'sb10110100001011110011001110100001011;
        end
        1540: begin
            cosine_reg0 <= 36'sb101001001110111111001010001100010000;
            sine_reg0   <= 36'sb10110011111001111011110000100100100;
        end
        1541: begin
            cosine_reg0 <= 36'sb101001001100110001111110001100011011;
            sine_reg0   <= 36'sb10110011101000000010100011101001001;
        end
        1542: begin
            cosine_reg0 <= 36'sb101001001010100101000000010000101110;
            sine_reg0   <= 36'sb10110011010110000111100111111010100;
        end
        1543: begin
            cosine_reg0 <= 36'sb101001001000011000010000011010011111;
            sine_reg0   <= 36'sb10110011000100001010111101100011101;
        end
        1544: begin
            cosine_reg0 <= 36'sb101001000110001011101110101011000110;
            sine_reg0   <= 36'sb10110010110010001100100100101111011;
        end
        1545: begin
            cosine_reg0 <= 36'sb101001000011111111011011000011111001;
            sine_reg0   <= 36'sb10110010100000001100011101101001001;
        end
        1546: begin
            cosine_reg0 <= 36'sb101001000001110011010101100110001110;
            sine_reg0   <= 36'sb10110010001110001010101000011011111;
        end
        1547: begin
            cosine_reg0 <= 36'sb101000111111100111011110010011011101;
            sine_reg0   <= 36'sb10110001111100000111000101010010110;
        end
        1548: begin
            cosine_reg0 <= 36'sb101000111101011011110101001100111011;
            sine_reg0   <= 36'sb10110001101010000001110100011000110;
        end
        1549: begin
            cosine_reg0 <= 36'sb101000111011010000011010010011111110;
            sine_reg0   <= 36'sb10110001010111111010110101111001010;
        end
        1550: begin
            cosine_reg0 <= 36'sb101000111001000101001101101001111101;
            sine_reg0   <= 36'sb10110001000101110010001001111111010;
        end
        1551: begin
            cosine_reg0 <= 36'sb101000110110111010001111010000001101;
            sine_reg0   <= 36'sb10110000110011100111110000110110001;
        end
        1552: begin
            cosine_reg0 <= 36'sb101000110100101111011111001000000101;
            sine_reg0   <= 36'sb10110000100001011011101010101000111;
        end
        1553: begin
            cosine_reg0 <= 36'sb101000110010100100111101010010111001;
            sine_reg0   <= 36'sb10110000001111001101110111100010110;
        end
        1554: begin
            cosine_reg0 <= 36'sb101000110000011010101001110001111111;
            sine_reg0   <= 36'sb10101111111100111110010111101111001;
        end
        1555: begin
            cosine_reg0 <= 36'sb101000101110010000100100100110101100;
            sine_reg0   <= 36'sb10101111101010101101001011011001001;
        end
        1556: begin
            cosine_reg0 <= 36'sb101000101100000110101101110010010111;
            sine_reg0   <= 36'sb10101111011000011010010010101100000;
        end
        1557: begin
            cosine_reg0 <= 36'sb101000101001111101000101010110010010;
            sine_reg0   <= 36'sb10101111000110000101101101110011001;
        end
        1558: begin
            cosine_reg0 <= 36'sb101000100111110011101011010011110101;
            sine_reg0   <= 36'sb10101110110011101111011100111001111;
        end
        1559: begin
            cosine_reg0 <= 36'sb101000100101101010011111101100010010;
            sine_reg0   <= 36'sb10101110100001010111100000001011011;
        end
        1560: begin
            cosine_reg0 <= 36'sb101000100011100001100010100001000000;
            sine_reg0   <= 36'sb10101110001110111101110111110011001;
        end
        1561: begin
            cosine_reg0 <= 36'sb101000100001011000110011110011010010;
            sine_reg0   <= 36'sb10101101111100100010100011111100010;
        end
        1562: begin
            cosine_reg0 <= 36'sb101000011111010000010011100100011101;
            sine_reg0   <= 36'sb10101101101010000101100100110010011;
        end
        1563: begin
            cosine_reg0 <= 36'sb101000011101001000000001110101110100;
            sine_reg0   <= 36'sb10101101010111100110111010100000110;
        end
        1564: begin
            cosine_reg0 <= 36'sb101000011010111111111110101000101101;
            sine_reg0   <= 36'sb10101101000101000110100101010010111;
        end
        1565: begin
            cosine_reg0 <= 36'sb101000011000111000001001111110011011;
            sine_reg0   <= 36'sb10101100110010100100100101010100000;
        end
        1566: begin
            cosine_reg0 <= 36'sb101000010110110000100011111000010001;
            sine_reg0   <= 36'sb10101100100000000000111010101111101;
        end
        1567: begin
            cosine_reg0 <= 36'sb101000010100101001001100010111100100;
            sine_reg0   <= 36'sb10101100001101011011100101110001010;
        end
        1568: begin
            cosine_reg0 <= 36'sb101000010010100010000011011101100110;
            sine_reg0   <= 36'sb10101011111010110100100110100100011;
        end
        1569: begin
            cosine_reg0 <= 36'sb101000010000011011001001001011101100;
            sine_reg0   <= 36'sb10101011101000001011111101010100010;
        end
        1570: begin
            cosine_reg0 <= 36'sb101000001110010100011101100011001000;
            sine_reg0   <= 36'sb10101011010101100001101010001100101;
        end
        1571: begin
            cosine_reg0 <= 36'sb101000001100001110000000100101001110;
            sine_reg0   <= 36'sb10101011000010110101101101011000111;
        end
        1572: begin
            cosine_reg0 <= 36'sb101000001010000111110010010011010000;
            sine_reg0   <= 36'sb10101010110000001000000111000100101;
        end
        1573: begin
            cosine_reg0 <= 36'sb101000001000000001110010101110100001;
            sine_reg0   <= 36'sb10101010011101011000110111011011011;
        end
        1574: begin
            cosine_reg0 <= 36'sb101000000101111100000001111000010101;
            sine_reg0   <= 36'sb10101010001010100111111110101000101;
        end
        1575: begin
            cosine_reg0 <= 36'sb101000000011110110011111110001111100;
            sine_reg0   <= 36'sb10101001110111110101011100111000000;
        end
        1576: begin
            cosine_reg0 <= 36'sb101000000001110001001100011100101011;
            sine_reg0   <= 36'sb10101001100101000001010010010101000;
        end
        1577: begin
            cosine_reg0 <= 36'sb100111111111101100000111111001110011;
            sine_reg0   <= 36'sb10101001010010001011011111001011011;
        end
        1578: begin
            cosine_reg0 <= 36'sb100111111101100111010010001010100101;
            sine_reg0   <= 36'sb10101000111111010100000011100110110;
        end
        1579: begin
            cosine_reg0 <= 36'sb100111111011100010101011010000010101;
            sine_reg0   <= 36'sb10101000101100011010111111110010101;
        end
        1580: begin
            cosine_reg0 <= 36'sb100111111001011110010011001100010011;
            sine_reg0   <= 36'sb10101000011001100000010011111010110;
        end
        1581: begin
            cosine_reg0 <= 36'sb100111110111011010001001111111110010;
            sine_reg0   <= 36'sb10101000000110100100000000001010110;
        end
        1582: begin
            cosine_reg0 <= 36'sb100111110101010110001111101100000011;
            sine_reg0   <= 36'sb10100111110011100110000100101110011;
        end
        1583: begin
            cosine_reg0 <= 36'sb100111110011010010100100010010011000;
            sine_reg0   <= 36'sb10100111100000100110100001110001001;
        end
        1584: begin
            cosine_reg0 <= 36'sb100111110001001111000111110100000001;
            sine_reg0   <= 36'sb10100111001101100101010111011111000;
        end
        1585: begin
            cosine_reg0 <= 36'sb100111101111001011111010010010010000;
            sine_reg0   <= 36'sb10100110111010100010100110000011101;
        end
        1586: begin
            cosine_reg0 <= 36'sb100111101101001000111011101110010101;
            sine_reg0   <= 36'sb10100110100111011110001101101010110;
        end
        1587: begin
            cosine_reg0 <= 36'sb100111101011000110001100001001100010;
            sine_reg0   <= 36'sb10100110010100011000001110100000000;
        end
        1588: begin
            cosine_reg0 <= 36'sb100111101001000011101011100101000110;
            sine_reg0   <= 36'sb10100110000001010000101000101111010;
        end
        1589: begin
            cosine_reg0 <= 36'sb100111100111000001011010000010010100;
            sine_reg0   <= 36'sb10100101101110000111011100100100011;
        end
        1590: begin
            cosine_reg0 <= 36'sb100111100100111111010111100010011010;
            sine_reg0   <= 36'sb10100101011010111100101010001011001;
        end
        1591: begin
            cosine_reg0 <= 36'sb100111100010111101100100000110101010;
            sine_reg0   <= 36'sb10100101000111110000010001101111011;
        end
        1592: begin
            cosine_reg0 <= 36'sb100111100000111011111111110000010010;
            sine_reg0   <= 36'sb10100100110100100010010011011100110;
        end
        1593: begin
            cosine_reg0 <= 36'sb100111011110111010101010100000100100;
            sine_reg0   <= 36'sb10100100100001010010101111011111011;
        end
        1594: begin
            cosine_reg0 <= 36'sb100111011100111001100100011000101111;
            sine_reg0   <= 36'sb10100100001110000001100110000011000;
        end
        1595: begin
            cosine_reg0 <= 36'sb100111011010111000101101011010000010;
            sine_reg0   <= 36'sb10100011111010101110110111010011011;
        end
        1596: begin
            cosine_reg0 <= 36'sb100111011000111000000101100101101101;
            sine_reg0   <= 36'sb10100011100111011010100011011100101;
        end
        1597: begin
            cosine_reg0 <= 36'sb100111010110110111101100111101000000;
            sine_reg0   <= 36'sb10100011010100000100101010101010101;
        end
        1598: begin
            cosine_reg0 <= 36'sb100111010100110111100011100001001001;
            sine_reg0   <= 36'sb10100011000000101101001101001001010;
        end
        1599: begin
            cosine_reg0 <= 36'sb100111010010110111101001010011011000;
            sine_reg0   <= 36'sb10100010101101010100001011000100100;
        end
        1600: begin
            cosine_reg0 <= 36'sb100111010000110111111110010100111100;
            sine_reg0   <= 36'sb10100010011001111001100100101000010;
        end
        1601: begin
            cosine_reg0 <= 36'sb100111001110111000100010100111000010;
            sine_reg0   <= 36'sb10100010000110011101011010000000100;
        end
        1602: begin
            cosine_reg0 <= 36'sb100111001100111001010110001010111011;
            sine_reg0   <= 36'sb10100001110010111111101011011001010;
        end
        1603: begin
            cosine_reg0 <= 36'sb100111001010111010011001000001110100;
            sine_reg0   <= 36'sb10100001011111100000011000111110100;
        end
        1604: begin
            cosine_reg0 <= 36'sb100111001000111011101011001100111011;
            sine_reg0   <= 36'sb10100001001011111111100010111100011;
        end
        1605: begin
            cosine_reg0 <= 36'sb100111000110111101001100101101011111;
            sine_reg0   <= 36'sb10100000111000011101001001011110110;
        end
        1606: begin
            cosine_reg0 <= 36'sb100111000100111110111101100100101111;
            sine_reg0   <= 36'sb10100000100100111001001100110001111;
        end
        1607: begin
            cosine_reg0 <= 36'sb100111000011000000111101110011110111;
            sine_reg0   <= 36'sb10100000010001010011101101000001101;
        end
        1608: begin
            cosine_reg0 <= 36'sb100111000001000011001101011100000101;
            sine_reg0   <= 36'sb10011111111101101100101010011010001;
        end
        1609: begin
            cosine_reg0 <= 36'sb100110111111000101101100011110100111;
            sine_reg0   <= 36'sb10011111101010000100000101000111100;
        end
        1610: begin
            cosine_reg0 <= 36'sb100110111101001000011010111100101011;
            sine_reg0   <= 36'sb10011111010110011001111101010101111;
        end
        1611: begin
            cosine_reg0 <= 36'sb100110111011001011011000110111011101;
            sine_reg0   <= 36'sb10011111000010101110010011010001011;
        end
        1612: begin
            cosine_reg0 <= 36'sb100110111001001110100110010000001100;
            sine_reg0   <= 36'sb10011110101111000001000111000110001;
        end
        1613: begin
            cosine_reg0 <= 36'sb100110110111010010000011001000000011;
            sine_reg0   <= 36'sb10011110011011010010011001000000010;
        end
        1614: begin
            cosine_reg0 <= 36'sb100110110101010101101111100000001111;
            sine_reg0   <= 36'sb10011110000111100010001001001100000;
        end
        1615: begin
            cosine_reg0 <= 36'sb100110110011011001101011011001111110;
            sine_reg0   <= 36'sb10011101110011110000010111110101100;
        end
        1616: begin
            cosine_reg0 <= 36'sb100110110001011101110110110110011100;
            sine_reg0   <= 36'sb10011101011111111101000101001000111;
        end
        1617: begin
            cosine_reg0 <= 36'sb100110101111100010010001110110110101;
            sine_reg0   <= 36'sb10011101001100001000010001010010101;
        end
        1618: begin
            cosine_reg0 <= 36'sb100110101101100110111100011100010110;
            sine_reg0   <= 36'sb10011100111000010001111100011110101;
        end
        1619: begin
            cosine_reg0 <= 36'sb100110101011101011110110101000001010;
            sine_reg0   <= 36'sb10011100100100011010000110111001011;
        end
        1620: begin
            cosine_reg0 <= 36'sb100110101001110001000000011011011101;
            sine_reg0   <= 36'sb10011100010000100000110000101110111;
        end
        1621: begin
            cosine_reg0 <= 36'sb100110100111110110011001110111011100;
            sine_reg0   <= 36'sb10011011111100100101111010001011110;
        end
        1622: begin
            cosine_reg0 <= 36'sb100110100101111100000010111101010001;
            sine_reg0   <= 36'sb10011011101000101001100011011100000;
        end
        1623: begin
            cosine_reg0 <= 36'sb100110100100000001111011101110001001;
            sine_reg0   <= 36'sb10011011010100101011101100101100000;
        end
        1624: begin
            cosine_reg0 <= 36'sb100110100010001000000100001011001111;
            sine_reg0   <= 36'sb10011011000000101100010110001000001;
        end
        1625: begin
            cosine_reg0 <= 36'sb100110100000001110011100010101101101;
            sine_reg0   <= 36'sb10011010101100101011011111111100101;
        end
        1626: begin
            cosine_reg0 <= 36'sb100110011110010101000100001110101111;
            sine_reg0   <= 36'sb10011010011000101001001010010110000;
        end
        1627: begin
            cosine_reg0 <= 36'sb100110011100011011111011110111100000;
            sine_reg0   <= 36'sb10011010000100100101010101100000011;
        end
        1628: begin
            cosine_reg0 <= 36'sb100110011010100011000011010001001011;
            sine_reg0   <= 36'sb10011001110000100000000001101000011;
        end
        1629: begin
            cosine_reg0 <= 36'sb100110011000101010011010011100111001;
            sine_reg0   <= 36'sb10011001011100011001001110111010001;
        end
        1630: begin
            cosine_reg0 <= 36'sb100110010110110010000001011011110110;
            sine_reg0   <= 36'sb10011001001000010000111101100010010;
        end
        1631: begin
            cosine_reg0 <= 36'sb100110010100111001111000001111001100;
            sine_reg0   <= 36'sb10011000110100000111001101101101000;
        end
        1632: begin
            cosine_reg0 <= 36'sb100110010011000001111110111000000100;
            sine_reg0   <= 36'sb10011000011111111011111111100111000;
        end
        1633: begin
            cosine_reg0 <= 36'sb100110010001001010010101010111101001;
            sine_reg0   <= 36'sb10011000001011101111010011011100100;
        end
        1634: begin
            cosine_reg0 <= 36'sb100110001111010010111011101111000101;
            sine_reg0   <= 36'sb10010111110111100001001001011010000;
        end
        1635: begin
            cosine_reg0 <= 36'sb100110001101011011110001111111100001;
            sine_reg0   <= 36'sb10010111100011010001100001101100001;
        end
        1636: begin
            cosine_reg0 <= 36'sb100110001011100100111000001010000110;
            sine_reg0   <= 36'sb10010111001111000000011100011111010;
        end
        1637: begin
            cosine_reg0 <= 36'sb100110001001101110001110001111111111;
            sine_reg0   <= 36'sb10010110111010101101111001111111110;
        end
        1638: begin
            cosine_reg0 <= 36'sb100110000111110111110100010010010100;
            sine_reg0   <= 36'sb10010110100110011001111010011010011;
        end
        1639: begin
            cosine_reg0 <= 36'sb100110000110000001101010010010001110;
            sine_reg0   <= 36'sb10010110010010000100011101111011100;
        end
        1640: begin
            cosine_reg0 <= 36'sb100110000100001011110000010000110110;
            sine_reg0   <= 36'sb10010101111101101101100100101111110;
        end
        1641: begin
            cosine_reg0 <= 36'sb100110000010010110000110001111010110;
            sine_reg0   <= 36'sb10010101101001010101001111000011101;
        end
        1642: begin
            cosine_reg0 <= 36'sb100110000000100000101100001110110100;
            sine_reg0   <= 36'sb10010101010100111011011101000011110;
        end
        1643: begin
            cosine_reg0 <= 36'sb100101111110101011100010010000011011;
            sine_reg0   <= 36'sb10010101000000100000001110111100101;
        end
        1644: begin
            cosine_reg0 <= 36'sb100101111100110110101000010101010010;
            sine_reg0   <= 36'sb10010100101100000011100100111011000;
        end
        1645: begin
            cosine_reg0 <= 36'sb100101111011000001111110011110100001;
            sine_reg0   <= 36'sb10010100010111100101011111001011011;
        end
        1646: begin
            cosine_reg0 <= 36'sb100101111001001101100100101101010001;
            sine_reg0   <= 36'sb10010100000011000101111101111010011;
        end
        1647: begin
            cosine_reg0 <= 36'sb100101110111011001011011000010101000;
            sine_reg0   <= 36'sb10010011101110100101000001010100101;
        end
        1648: begin
            cosine_reg0 <= 36'sb100101110101100101100001011111101111;
            sine_reg0   <= 36'sb10010011011010000010101001100110111;
        end
        1649: begin
            cosine_reg0 <= 36'sb100101110011110001111000000101101110;
            sine_reg0   <= 36'sb10010011000101011110110110111101101;
        end
        1650: begin
            cosine_reg0 <= 36'sb100101110001111110011110110101101011;
            sine_reg0   <= 36'sb10010010110000111001101001100101110;
        end
        1651: begin
            cosine_reg0 <= 36'sb100101110000001011010101110000101101;
            sine_reg0   <= 36'sb10010010011100010011000001101011111;
        end
        1652: begin
            cosine_reg0 <= 36'sb100101101110011000011100110111111100;
            sine_reg0   <= 36'sb10010010000111101010111111011100110;
        end
        1653: begin
            cosine_reg0 <= 36'sb100101101100100101110100001100011111;
            sine_reg0   <= 36'sb10010001110011000001100011000100111;
        end
        1654: begin
            cosine_reg0 <= 36'sb100101101010110011011011101111011101;
            sine_reg0   <= 36'sb10010001011110010110101100110001010;
        end
        1655: begin
            cosine_reg0 <= 36'sb100101101001000001010011100001111011;
            sine_reg0   <= 36'sb10010001001001101010011100101110101;
        end
        1656: begin
            cosine_reg0 <= 36'sb100101100111001111011011100101000000;
            sine_reg0   <= 36'sb10010000110100111100110011001001100;
        end
        1657: begin
            cosine_reg0 <= 36'sb100101100101011101110011111001110011;
            sine_reg0   <= 36'sb10010000100000001101110000001111000;
        end
        1658: begin
            cosine_reg0 <= 36'sb100101100011101100011100100001011001;
            sine_reg0   <= 36'sb10010000001011011101010100001011101;
        end
        1659: begin
            cosine_reg0 <= 36'sb100101100001111011010101011100111010;
            sine_reg0   <= 36'sb10001111110110101011011111001100010;
        end
        1660: begin
            cosine_reg0 <= 36'sb100101100000001010011110101101011001;
            sine_reg0   <= 36'sb10001111100001111000010001011101111;
        end
        1661: begin
            cosine_reg0 <= 36'sb100101011110011001111000010011111101;
            sine_reg0   <= 36'sb10001111001101000011101011001101000;
        end
        1662: begin
            cosine_reg0 <= 36'sb100101011100101001100010010001101100;
            sine_reg0   <= 36'sb10001110111000001101101100100110111;
        end
        1663: begin
            cosine_reg0 <= 36'sb100101011010111001011100100111101010;
            sine_reg0   <= 36'sb10001110100011010110010101111000000;
        end
        1664: begin
            cosine_reg0 <= 36'sb100101011001001001100111010110111101;
            sine_reg0   <= 36'sb10001110001110011101100111001101011;
        end
        1665: begin
            cosine_reg0 <= 36'sb100101010111011010000010100000101010;
            sine_reg0   <= 36'sb10001101111001100011100000110100000;
        end
        1666: begin
            cosine_reg0 <= 36'sb100101010101101010101110000101110110;
            sine_reg0   <= 36'sb10001101100100101000000010111000100;
        end
        1667: begin
            cosine_reg0 <= 36'sb100101010011111011101010000111100100;
            sine_reg0   <= 36'sb10001101001111101011001101101000001;
        end
        1668: begin
            cosine_reg0 <= 36'sb100101010010001100110110100110111011;
            sine_reg0   <= 36'sb10001100111010101101000001001111100;
        end
        1669: begin
            cosine_reg0 <= 36'sb100101010000011110010011100100111110;
            sine_reg0   <= 36'sb10001100100101101101011101111011110;
        end
        1670: begin
            cosine_reg0 <= 36'sb100101001110110000000001000010110001;
            sine_reg0   <= 36'sb10001100010000101100100011111001110;
        end
        1671: begin
            cosine_reg0 <= 36'sb100101001101000001111111000001011001;
            sine_reg0   <= 36'sb10001011111011101010010011010110100;
        end
        1672: begin
            cosine_reg0 <= 36'sb100101001011010100001101100001111000;
            sine_reg0   <= 36'sb10001011100110100110101100011110111;
        end
        1673: begin
            cosine_reg0 <= 36'sb100101001001100110101100100101010100;
            sine_reg0   <= 36'sb10001011010001100001101111100000000;
        end
        1674: begin
            cosine_reg0 <= 36'sb100101000111111001011100001100101111;
            sine_reg0   <= 36'sb10001010111100011011011100100110110;
        end
        1675: begin
            cosine_reg0 <= 36'sb100101000110001100011100011001001110;
            sine_reg0   <= 36'sb10001010100111010011110100000000010;
        end
        1676: begin
            cosine_reg0 <= 36'sb100101000100011111101101001011110010;
            sine_reg0   <= 36'sb10001010010010001010110101111001100;
        end
        1677: begin
            cosine_reg0 <= 36'sb100101000010110011001110100101011111;
            sine_reg0   <= 36'sb10001001111101000000100010011111100;
        end
        1678: begin
            cosine_reg0 <= 36'sb100101000001000111000000100111011001;
            sine_reg0   <= 36'sb10001001100111110100111001111111011;
        end
        1679: begin
            cosine_reg0 <= 36'sb100100111111011011000011010010100010;
            sine_reg0   <= 36'sb10001001010010100111111100100110001;
        end
        1680: begin
            cosine_reg0 <= 36'sb100100111101101111010110100111111100;
            sine_reg0   <= 36'sb10001000111101011001101010100000110;
        end
        1681: begin
            cosine_reg0 <= 36'sb100100111100000011111010101000101010;
            sine_reg0   <= 36'sb10001000101000001010000011111100100;
        end
        1682: begin
            cosine_reg0 <= 36'sb100100111010011000101111010101101110;
            sine_reg0   <= 36'sb10001000010010111001001001000110100;
        end
        1683: begin
            cosine_reg0 <= 36'sb100100111000101101110100110000001010;
            sine_reg0   <= 36'sb10000111111101100110111010001011101;
        end
        1684: begin
            cosine_reg0 <= 36'sb100100110111000011001010111001000001;
            sine_reg0   <= 36'sb10000111101000010011010111011001010;
        end
        1685: begin
            cosine_reg0 <= 36'sb100100110101011000110001110001010100;
            sine_reg0   <= 36'sb10000111010010111110100000111100011;
        end
        1686: begin
            cosine_reg0 <= 36'sb100100110011101110101001011010000100;
            sine_reg0   <= 36'sb10000110111101101000010111000010010;
        end
        1687: begin
            cosine_reg0 <= 36'sb100100110010000100110001110100010100;
            sine_reg0   <= 36'sb10000110101000010000111001111000000;
        end
        1688: begin
            cosine_reg0 <= 36'sb100100110000011011001011000001000100;
            sine_reg0   <= 36'sb10000110010010111000001001101010111;
        end
        1689: begin
            cosine_reg0 <= 36'sb100100101110110001110101000001010101;
            sine_reg0   <= 36'sb10000101111101011110000110100111111;
        end
        1690: begin
            cosine_reg0 <= 36'sb100100101101001000101111110110001001;
            sine_reg0   <= 36'sb10000101101000000010110000111100011;
        end
        1691: begin
            cosine_reg0 <= 36'sb100100101011011111111011100000100001;
            sine_reg0   <= 36'sb10000101010010100110001000110101101;
        end
        1692: begin
            cosine_reg0 <= 36'sb100100101001110111011000000001011100;
            sine_reg0   <= 36'sb10000100111101001000001110100000101;
        end
        1693: begin
            cosine_reg0 <= 36'sb100100101000001111000101011001111100;
            sine_reg0   <= 36'sb10000100100111101001000010001010111;
        end
        1694: begin
            cosine_reg0 <= 36'sb100100100110100111000011101011000001;
            sine_reg0   <= 36'sb10000100010010001000100100000001100;
        end
        1695: begin
            cosine_reg0 <= 36'sb100100100100111111010010110101101011;
            sine_reg0   <= 36'sb10000011111100100110110100010001110;
        end
        1696: begin
            cosine_reg0 <= 36'sb100100100011010111110010111010111011;
            sine_reg0   <= 36'sb10000011100111000011110011001001000;
        end
        1697: begin
            cosine_reg0 <= 36'sb100100100001110000100011111011101110;
            sine_reg0   <= 36'sb10000011010001011111100000110100100;
        end
        1698: begin
            cosine_reg0 <= 36'sb100100100000001001100101111001000111;
            sine_reg0   <= 36'sb10000010111011111001111101100001100;
        end
        1699: begin
            cosine_reg0 <= 36'sb100100011110100010111000110100000100;
            sine_reg0   <= 36'sb10000010100110010011001001011101011;
        end
        1700: begin
            cosine_reg0 <= 36'sb100100011100111100011100101101100100;
            sine_reg0   <= 36'sb10000010010000101011000100110101011;
        end
        1701: begin
            cosine_reg0 <= 36'sb100100011011010110010001100110100110;
            sine_reg0   <= 36'sb10000001111011000001101111110110111;
        end
        1702: begin
            cosine_reg0 <= 36'sb100100011001110000010111100000001011;
            sine_reg0   <= 36'sb10000001100101010111001010101111011;
        end
        1703: begin
            cosine_reg0 <= 36'sb100100011000001010101110011011001111;
            sine_reg0   <= 36'sb10000001001111101011010101101100000;
        end
        1704: begin
            cosine_reg0 <= 36'sb100100010110100101010110011000110011;
            sine_reg0   <= 36'sb10000000111001111110010000111010011;
        end
        1705: begin
            cosine_reg0 <= 36'sb100100010101000000001111011001110101;
            sine_reg0   <= 36'sb10000000100100001111111100100111101;
        end
        1706: begin
            cosine_reg0 <= 36'sb100100010011011011011001011111010011;
            sine_reg0   <= 36'sb10000000001110100000011001000001010;
        end
        1707: begin
            cosine_reg0 <= 36'sb100100010001110110110100101010001011;
            sine_reg0   <= 36'sb1111111111000101111100110010100110;
        end
        1708: begin
            cosine_reg0 <= 36'sb100100010000010010100000111011011100;
            sine_reg0   <= 36'sb1111111100010111101100100101111100;
        end
        1709: begin
            cosine_reg0 <= 36'sb100100001110101110011110010100000011;
            sine_reg0   <= 36'sb1111111001101001010010100011111000;
        end
        1710: begin
            cosine_reg0 <= 36'sb100100001101001010101100110100111110;
            sine_reg0   <= 36'sb1111110110111010101110101110000100;
        end
        1711: begin
            cosine_reg0 <= 36'sb100100001011100111001100011111001010;
            sine_reg0   <= 36'sb1111110100001100000001000110001101;
        end
        1712: begin
            cosine_reg0 <= 36'sb100100001010000011111101010011100101;
            sine_reg0   <= 36'sb1111110001011101001001101101111111;
        end
        1713: begin
            cosine_reg0 <= 36'sb100100001000100000111111010011001100;
            sine_reg0   <= 36'sb1111101110101110001000100111000100;
        end
        1714: begin
            cosine_reg0 <= 36'sb100100000110111110010010011110111101;
            sine_reg0   <= 36'sb1111101011111110111101110011001010;
        end
        1715: begin
            cosine_reg0 <= 36'sb100100000101011011110110110111110011;
            sine_reg0   <= 36'sb1111101001001111101001010011111101;
        end
        1716: begin
            cosine_reg0 <= 36'sb100100000011111001101100011110101100;
            sine_reg0   <= 36'sb1111100110100000001011001011000111;
        end
        1717: begin
            cosine_reg0 <= 36'sb100100000010010111110011010100100100;
            sine_reg0   <= 36'sb1111100011110000100011011010010111;
        end
        1718: begin
            cosine_reg0 <= 36'sb100100000000110110001011011010011000;
            sine_reg0   <= 36'sb1111100001000000110010000011011000;
        end
        1719: begin
            cosine_reg0 <= 36'sb100011111111010100110100110001000100;
            sine_reg0   <= 36'sb1111011110010000110111000111110101;
        end
        1720: begin
            cosine_reg0 <= 36'sb100011111101110011101111011001100100;
            sine_reg0   <= 36'sb1111011011100000110010101001011101;
        end
        1721: begin
            cosine_reg0 <= 36'sb100011111100010010111011010100110100;
            sine_reg0   <= 36'sb1111011000110000100100101001111100;
        end
        1722: begin
            cosine_reg0 <= 36'sb100011111010110010011000100011101111;
            sine_reg0   <= 36'sb1111010110000000001101001010111110;
        end
        1723: begin
            cosine_reg0 <= 36'sb100011111001010010000111000111010010;
            sine_reg0   <= 36'sb1111010011001111101100001110010000;
        end
        1724: begin
            cosine_reg0 <= 36'sb100011110111110010000111000000010111;
            sine_reg0   <= 36'sb1111010000011111000001110101011111;
        end
        1725: begin
            cosine_reg0 <= 36'sb100011110110010010011000001111111001;
            sine_reg0   <= 36'sb1111001101101110001110000010010111;
        end
        1726: begin
            cosine_reg0 <= 36'sb100011110100110010111010110110110100;
            sine_reg0   <= 36'sb1111001010111101010000110110100111;
        end
        1727: begin
            cosine_reg0 <= 36'sb100011110011010011101110110110000011;
            sine_reg0   <= 36'sb1111001000001100001010010011111011;
        end
        1728: begin
            cosine_reg0 <= 36'sb100011110001110100110100001110100001;
            sine_reg0   <= 36'sb1111000101011010111010011100000000;
        end
        1729: begin
            cosine_reg0 <= 36'sb100011110000010110001011000001000111;
            sine_reg0   <= 36'sb1111000010101001100001010000100100;
        end
        1730: begin
            cosine_reg0 <= 36'sb100011101110110111110011001110110000;
            sine_reg0   <= 36'sb1110111111110111111110110011010101;
        end
        1731: begin
            cosine_reg0 <= 36'sb100011101101011001101100111000010111;
            sine_reg0   <= 36'sb1110111101000110010011000101111111;
        end
        1732: begin
            cosine_reg0 <= 36'sb100011101011111011110111111110110110;
            sine_reg0   <= 36'sb1110111010010100011110001010010000;
        end
        1733: begin
            cosine_reg0 <= 36'sb100011101010011110010100100011000110;
            sine_reg0   <= 36'sb1110110111100010100000000001110110;
        end
        1734: begin
            cosine_reg0 <= 36'sb100011101001000001000010100110000001;
            sine_reg0   <= 36'sb1110110100110000011000101110011111;
        end
        1735: begin
            cosine_reg0 <= 36'sb100011100111100100000010001000100001;
            sine_reg0   <= 36'sb1110110001111110001000010001111000;
        end
        1736: begin
            cosine_reg0 <= 36'sb100011100110000111010011001011011111;
            sine_reg0   <= 36'sb1110101111001011101110101101110000;
        end
        1737: begin
            cosine_reg0 <= 36'sb100011100100101010110101101111110100;
            sine_reg0   <= 36'sb1110101100011001001100000011110101;
        end
        1738: begin
            cosine_reg0 <= 36'sb100011100011001110101001110110011001;
            sine_reg0   <= 36'sb1110101001100110100000010101110101;
        end
        1739: begin
            cosine_reg0 <= 36'sb100011100001110010101111100000001000;
            sine_reg0   <= 36'sb1110100110110011101011100101011101;
        end
        1740: begin
            cosine_reg0 <= 36'sb100011100000010111000110101101111000;
            sine_reg0   <= 36'sb1110100100000000101101110100011101;
        end
        1741: begin
            cosine_reg0 <= 36'sb100011011110111011101111100000100011;
            sine_reg0   <= 36'sb1110100001001101100111000100100010;
        end
        1742: begin
            cosine_reg0 <= 36'sb100011011101100000101001111001000000;
            sine_reg0   <= 36'sb1110011110011010010111010111011100;
        end
        1743: begin
            cosine_reg0 <= 36'sb100011011100000101110101111000001001;
            sine_reg0   <= 36'sb1110011011100110111110101110111000;
        end
        1744: begin
            cosine_reg0 <= 36'sb100011011010101011010011011110110100;
            sine_reg0   <= 36'sb1110011000110011011101001100100110;
        end
        1745: begin
            cosine_reg0 <= 36'sb100011011001010001000010101101111010;
            sine_reg0   <= 36'sb1110010101111111110010110010010100;
        end
        1746: begin
            cosine_reg0 <= 36'sb100011010111110111000011100110010010;
            sine_reg0   <= 36'sb1110010011001011111111100001110000;
        end
        1747: begin
            cosine_reg0 <= 36'sb100011010110011101010110001000110101;
            sine_reg0   <= 36'sb1110010000011000000011011100101011;
        end
        1748: begin
            cosine_reg0 <= 36'sb100011010101000011111010010110011001;
            sine_reg0   <= 36'sb1110001101100011111110100100110010;
        end
        1749: begin
            cosine_reg0 <= 36'sb100011010011101010110000001111110101;
            sine_reg0   <= 36'sb1110001010101111110000111011110110;
        end
        1750: begin
            cosine_reg0 <= 36'sb100011010010010001110111110110000001;
            sine_reg0   <= 36'sb1110000111111011011010100011100100;
        end
        1751: begin
            cosine_reg0 <= 36'sb100011010000111001010001001001110011;
            sine_reg0   <= 36'sb1110000101000110111011011101101101;
        end
        1752: begin
            cosine_reg0 <= 36'sb100011001111100000111100001100000010;
            sine_reg0   <= 36'sb1110000010010010010011101100000000;
        end
        1753: begin
            cosine_reg0 <= 36'sb100011001110001000111000111101100100;
            sine_reg0   <= 36'sb1101111111011101100011010000001011;
        end
        1754: begin
            cosine_reg0 <= 36'sb100011001100110001000111011111010000;
            sine_reg0   <= 36'sb1101111100101000101010001100000000;
        end
        1755: begin
            cosine_reg0 <= 36'sb100011001011011001100111110001111100;
            sine_reg0   <= 36'sb1101111001110011101000100001001100;
        end
        1756: begin
            cosine_reg0 <= 36'sb100011001010000010011001110110011110;
            sine_reg0   <= 36'sb1101110110111110011110010001100000;
        end
        1757: begin
            cosine_reg0 <= 36'sb100011001000101011011101101101101100;
            sine_reg0   <= 36'sb1101110100001001001011011110101100;
        end
        1758: begin
            cosine_reg0 <= 36'sb100011000111010100110011011000011010;
            sine_reg0   <= 36'sb1101110001010011110000001010011111;
        end
        1759: begin
            cosine_reg0 <= 36'sb100011000101111110011010110111100000;
            sine_reg0   <= 36'sb1101101110011110001100010110101010;
        end
        1760: begin
            cosine_reg0 <= 36'sb100011000100101000010100001011110010;
            sine_reg0   <= 36'sb1101101011101000100000000100111100;
        end
        1761: begin
            cosine_reg0 <= 36'sb100011000011010010011111010110000100;
            sine_reg0   <= 36'sb1101101000110010101011010111000101;
        end
        1762: begin
            cosine_reg0 <= 36'sb100011000001111100111100010111001101;
            sine_reg0   <= 36'sb1101100101111100101110001110110110;
        end
        1763: begin
            cosine_reg0 <= 36'sb100011000000100111101011010000000001;
            sine_reg0   <= 36'sb1101100011000110101000101101111111;
        end
        1764: begin
            cosine_reg0 <= 36'sb100010111111010010101100000001010100;
            sine_reg0   <= 36'sb1101100000010000011010110110001111;
        end
        1765: begin
            cosine_reg0 <= 36'sb100010111101111101111110101011111011;
            sine_reg0   <= 36'sb1101011101011010000100101001011001;
        end
        1766: begin
            cosine_reg0 <= 36'sb100010111100101001100011010000101010;
            sine_reg0   <= 36'sb1101011010100011100110001001001011;
        end
        1767: begin
            cosine_reg0 <= 36'sb100010111011010101011001110000010110;
            sine_reg0   <= 36'sb1101010111101100111111010111010111;
        end
        1768: begin
            cosine_reg0 <= 36'sb100010111010000001100010001011110001;
            sine_reg0   <= 36'sb1101010100110110010000010101101101;
        end
        1769: begin
            cosine_reg0 <= 36'sb100010111000101101111100100011110001;
            sine_reg0   <= 36'sb1101010001111111011001000101111110;
        end
        1770: begin
            cosine_reg0 <= 36'sb100010110111011010101000111001000111;
            sine_reg0   <= 36'sb1101001111001000011001101001111011;
        end
        1771: begin
            cosine_reg0 <= 36'sb100010110110000111100111001100101001;
            sine_reg0   <= 36'sb1101001100010001010010000011010100;
        end
        1772: begin
            cosine_reg0 <= 36'sb100010110100110100110111011111001001;
            sine_reg0   <= 36'sb1101001001011010000010010011111011;
        end
        1773: begin
            cosine_reg0 <= 36'sb100010110011100010011001110001011001;
            sine_reg0   <= 36'sb1101000110100010101010011101100001;
        end
        1774: begin
            cosine_reg0 <= 36'sb100010110010010000001110000100001110;
            sine_reg0   <= 36'sb1101000011101011001010100001110110;
        end
        1775: begin
            cosine_reg0 <= 36'sb100010110000111110010100011000011001;
            sine_reg0   <= 36'sb1101000000110011100010100010101100;
        end
        1776: begin
            cosine_reg0 <= 36'sb100010101111101100101100101110101101;
            sine_reg0   <= 36'sb1100111101111011110010100001110101;
        end
        1777: begin
            cosine_reg0 <= 36'sb100010101110011011010111000111111101;
            sine_reg0   <= 36'sb1100111011000011111010100001000001;
        end
        1778: begin
            cosine_reg0 <= 36'sb100010101101001010010011100100111011;
            sine_reg0   <= 36'sb1100111000001011111010100010000001;
        end
        1779: begin
            cosine_reg0 <= 36'sb100010101011111001100010000110011000;
            sine_reg0   <= 36'sb1100110101010011110010100110101001;
        end
        1780: begin
            cosine_reg0 <= 36'sb100010101010101001000010101101000111;
            sine_reg0   <= 36'sb1100110010011011100010110000101000;
        end
        1781: begin
            cosine_reg0 <= 36'sb100010101001011000110101011001111000;
            sine_reg0   <= 36'sb1100101111100011001011000001110001;
        end
        1782: begin
            cosine_reg0 <= 36'sb100010101000001000111010001101011111;
            sine_reg0   <= 36'sb1100101100101010101011011011110101;
        end
        1783: begin
            cosine_reg0 <= 36'sb100010100110111001010001001000101011;
            sine_reg0   <= 36'sb1100101001110010000100000000100111;
        end
        1784: begin
            cosine_reg0 <= 36'sb100010100101101001111010001100001110;
            sine_reg0   <= 36'sb1100100110111001010100110001110111;
        end
        1785: begin
            cosine_reg0 <= 36'sb100010100100011010110101011000111010;
            sine_reg0   <= 36'sb1100100100000000011101110001011001;
        end
        1786: begin
            cosine_reg0 <= 36'sb100010100011001100000010101111011110;
            sine_reg0   <= 36'sb1100100001000111011111000000111110;
        end
        1787: begin
            cosine_reg0 <= 36'sb100010100001111101100010010000101011;
            sine_reg0   <= 36'sb1100011110001110011000100010010111;
        end
        1788: begin
            cosine_reg0 <= 36'sb100010100000101111010011111101010011;
            sine_reg0   <= 36'sb1100011011010101001010010111011001;
        end
        1789: begin
            cosine_reg0 <= 36'sb100010011111100001010111110110000100;
            sine_reg0   <= 36'sb1100011000011011110100100001110100;
        end
        1790: begin
            cosine_reg0 <= 36'sb100010011110010011101101111011110000;
            sine_reg0   <= 36'sb1100010101100010010111000011011010;
        end
        1791: begin
            cosine_reg0 <= 36'sb100010011101000110010110001111000101;
            sine_reg0   <= 36'sb1100010010101000110001111101111111;
        end
        1792: begin
            cosine_reg0 <= 36'sb100010011011111001010000110000110100;
            sine_reg0   <= 36'sb1100001111101111000101010011010101;
        end
        1793: begin
            cosine_reg0 <= 36'sb100010011010101100011101100001101101;
            sine_reg0   <= 36'sb1100001100110101010001000101001111;
        end
        1794: begin
            cosine_reg0 <= 36'sb100010011001011111111100100010011110;
            sine_reg0   <= 36'sb1100001001111011010101010101011110;
        end
        1795: begin
            cosine_reg0 <= 36'sb100010011000010011101101110011110111;
            sine_reg0   <= 36'sb1100000111000001010010000101110110;
        end
        1796: begin
            cosine_reg0 <= 36'sb100010010111000111110001010110100111;
            sine_reg0   <= 36'sb1100000100000111000111011000001001;
        end
        1797: begin
            cosine_reg0 <= 36'sb100010010101111100000111001011011101;
            sine_reg0   <= 36'sb1100000001001100110101001110001011;
        end
        1798: begin
            cosine_reg0 <= 36'sb100010010100110000101111010011000111;
            sine_reg0   <= 36'sb1011111110010010011011101001101110;
        end
        1799: begin
            cosine_reg0 <= 36'sb100010010011100101101001101110010100;
            sine_reg0   <= 36'sb1011111011010111111010101100100101;
        end
        1800: begin
            cosine_reg0 <= 36'sb100010010010011010110110011101110011;
            sine_reg0   <= 36'sb1011111000011101010010011000100011;
        end
        1801: begin
            cosine_reg0 <= 36'sb100010010001010000010101100010010000;
            sine_reg0   <= 36'sb1011110101100010100010101111011100;
        end
        1802: begin
            cosine_reg0 <= 36'sb100010010000000110000110111100011100;
            sine_reg0   <= 36'sb1011110010100111101011110011000010;
        end
        1803: begin
            cosine_reg0 <= 36'sb100010001110111100001010101101000010;
            sine_reg0   <= 36'sb1011101111101100101101100101001001;
        end
        1804: begin
            cosine_reg0 <= 36'sb100010001101110010100000110100110001;
            sine_reg0   <= 36'sb1011101100110001101000000111100100;
        end
        1805: begin
            cosine_reg0 <= 36'sb100010001100101001001001010100010110;
            sine_reg0   <= 36'sb1011101001110110011011011100000111;
        end
        1806: begin
            cosine_reg0 <= 36'sb100010001011100000000100001100011110;
            sine_reg0   <= 36'sb1011100110111011000111100100100100;
        end
        1807: begin
            cosine_reg0 <= 36'sb100010001010010111010001011101110111;
            sine_reg0   <= 36'sb1011100011111111101100100010110001;
        end
        1808: begin
            cosine_reg0 <= 36'sb100010001001001110110001001001001110;
            sine_reg0   <= 36'sb1011100001000100001010011000011111;
        end
        1809: begin
            cosine_reg0 <= 36'sb100010001000000110100011001111001110;
            sine_reg0   <= 36'sb1011011110001000100001000111100011;
        end
        1810: begin
            cosine_reg0 <= 36'sb100010000110111110100111110000100110;
            sine_reg0   <= 36'sb1011011011001100110000110001110001;
        end
        1811: begin
            cosine_reg0 <= 36'sb100010000101110110111110101110000000;
            sine_reg0   <= 36'sb1011011000010000111001011000111100;
        end
        1812: begin
            cosine_reg0 <= 36'sb100010000100101111101000001000001001;
            sine_reg0   <= 36'sb1011010101010100111010111110111001;
        end
        1813: begin
            cosine_reg0 <= 36'sb100010000011101000100011111111101110;
            sine_reg0   <= 36'sb1011010010011000110101100101011010;
        end
        1814: begin
            cosine_reg0 <= 36'sb100010000010100001110010010101011010;
            sine_reg0   <= 36'sb1011001111011100101001001110010101;
        end
        1815: begin
            cosine_reg0 <= 36'sb100010000001011011010011001001111001;
            sine_reg0   <= 36'sb1011001100100000010101111011011110;
        end
        1816: begin
            cosine_reg0 <= 36'sb100010000000010101000110011101110110;
            sine_reg0   <= 36'sb1011001001100011111011101110101000;
        end
        1817: begin
            cosine_reg0 <= 36'sb100001111111001111001100010001111100;
            sine_reg0   <= 36'sb1011000110100111011010101001100111;
        end
        1818: begin
            cosine_reg0 <= 36'sb100001111110001001100100100110110111;
            sine_reg0   <= 36'sb1011000011101010110010101110010001;
        end
        1819: begin
            cosine_reg0 <= 36'sb100001111101000100001111011101010010;
            sine_reg0   <= 36'sb1011000000101110000011111110011001;
        end
        1820: begin
            cosine_reg0 <= 36'sb100001111011111111001100110101110111;
            sine_reg0   <= 36'sb1010111101110001001110011011110011;
        end
        1821: begin
            cosine_reg0 <= 36'sb100001111010111010011100110001010001;
            sine_reg0   <= 36'sb1010111010110100010010001000010110;
        end
        1822: begin
            cosine_reg0 <= 36'sb100001111001110101111111010000001010;
            sine_reg0   <= 36'sb1010110111110111001111000101110011;
        end
        1823: begin
            cosine_reg0 <= 36'sb100001111000110001110100010011001101;
            sine_reg0   <= 36'sb1010110100111010000101010110000010;
        end
        1824: begin
            cosine_reg0 <= 36'sb100001110111101101111011111011000011;
            sine_reg0   <= 36'sb1010110001111100110100111010110101;
        end
        1825: begin
            cosine_reg0 <= 36'sb100001110110101010010110001000010111;
            sine_reg0   <= 36'sb1010101110111111011101110110000010;
        end
        1826: begin
            cosine_reg0 <= 36'sb100001110101100111000010111011110011;
            sine_reg0   <= 36'sb1010101100000010000000001001011110;
        end
        1827: begin
            cosine_reg0 <= 36'sb100001110100100100000010010101111111;
            sine_reg0   <= 36'sb1010101001000100011011110110111110;
        end
        1828: begin
            cosine_reg0 <= 36'sb100001110011100001010100010111100101;
            sine_reg0   <= 36'sb1010100110000110110001000000010110;
        end
        1829: begin
            cosine_reg0 <= 36'sb100001110010011110111001000001001110;
            sine_reg0   <= 36'sb1010100011001000111111100111011011;
        end
        1830: begin
            cosine_reg0 <= 36'sb100001110001011100110000010011100011;
            sine_reg0   <= 36'sb1010100000001011000111101110000011;
        end
        1831: begin
            cosine_reg0 <= 36'sb100001110000011010111010001111001110;
            sine_reg0   <= 36'sb1010011101001101001001010110000010;
        end
        1832: begin
            cosine_reg0 <= 36'sb100001101111011001010110110100110110;
            sine_reg0   <= 36'sb1010011010001111000100100001001111;
        end
        1833: begin
            cosine_reg0 <= 36'sb100001101110011000000110000101000100;
            sine_reg0   <= 36'sb1010010111010000111001010001011101;
        end
        1834: begin
            cosine_reg0 <= 36'sb100001101101010111001000000000100000;
            sine_reg0   <= 36'sb1010010100010010100111101000100011;
        end
        1835: begin
            cosine_reg0 <= 36'sb100001101100010110011100100111110011;
            sine_reg0   <= 36'sb1010010001010100001111101000010110;
        end
        1836: begin
            cosine_reg0 <= 36'sb100001101011010110000011111011100100;
            sine_reg0   <= 36'sb1010001110010101110001010010101011;
        end
        1837: begin
            cosine_reg0 <= 36'sb100001101010010101111101111100011011;
            sine_reg0   <= 36'sb1010001011010111001100101001010111;
        end
        1838: begin
            cosine_reg0 <= 36'sb100001101001010110001010101011000000;
            sine_reg0   <= 36'sb1010001000011000100001101110010001;
        end
        1839: begin
            cosine_reg0 <= 36'sb100001101000010110101010000111111001;
            sine_reg0   <= 36'sb1010000101011001110000100011001101;
        end
        1840: begin
            cosine_reg0 <= 36'sb100001100111010111011100010011101111;
            sine_reg0   <= 36'sb1010000010011010111001001010000011;
        end
        1841: begin
            cosine_reg0 <= 36'sb100001100110011000100001001111000111;
            sine_reg0   <= 36'sb1001111111011011111011100100100110;
        end
        1842: begin
            cosine_reg0 <= 36'sb100001100101011001111000111010101010;
            sine_reg0   <= 36'sb1001111100011100110111110100101110;
        end
        1843: begin
            cosine_reg0 <= 36'sb100001100100011011100011010110111100;
            sine_reg0   <= 36'sb1001111001011101101101111100001111;
        end
        1844: begin
            cosine_reg0 <= 36'sb100001100011011101100000100100100110;
            sine_reg0   <= 36'sb1001110110011110011101111101000000;
        end
        1845: begin
            cosine_reg0 <= 36'sb100001100010011111110000100100001101;
            sine_reg0   <= 36'sb1001110011011111000111111000110111;
        end
        1846: begin
            cosine_reg0 <= 36'sb100001100001100010010011010110011000;
            sine_reg0   <= 36'sb1001110000011111101011110001101010;
        end
        1847: begin
            cosine_reg0 <= 36'sb100001100000100101001000111011101011;
            sine_reg0   <= 36'sb1001101101100000001001101001001111;
        end
        1848: begin
            cosine_reg0 <= 36'sb100001011111101000010001010100101110;
            sine_reg0   <= 36'sb1001101010100000100001100001011100;
        end
        1849: begin
            cosine_reg0 <= 36'sb100001011110101011101100100010000101;
            sine_reg0   <= 36'sb1001100111100000110011011100000111;
        end
        1850: begin
            cosine_reg0 <= 36'sb100001011101101111011010100100010110;
            sine_reg0   <= 36'sb1001100100100000111111011011000111;
        end
        1851: begin
            cosine_reg0 <= 36'sb100001011100110011011011011100000110;
            sine_reg0   <= 36'sb1001100001100001000101100000010001;
        end
        1852: begin
            cosine_reg0 <= 36'sb100001011011110111101111001001111001;
            sine_reg0   <= 36'sb1001011110100001000101101101011101;
        end
        1853: begin
            cosine_reg0 <= 36'sb100001011010111100010101101110010110;
            sine_reg0   <= 36'sb1001011011100001000000000100100001;
        end
        1854: begin
            cosine_reg0 <= 36'sb100001011010000001001111001010000001;
            sine_reg0   <= 36'sb1001011000100000110100100111010010;
        end
        1855: begin
            cosine_reg0 <= 36'sb100001011001000110011011011101011101;
            sine_reg0   <= 36'sb1001010101100000100011010111101001;
        end
        1856: begin
            cosine_reg0 <= 36'sb100001011000001011111010101001001111;
            sine_reg0   <= 36'sb1001010010100000001100010111011010;
        end
        1857: begin
            cosine_reg0 <= 36'sb100001010111010001101100101101111100;
            sine_reg0   <= 36'sb1001001111011111101111101000011110;
        end
        1858: begin
            cosine_reg0 <= 36'sb100001010110010111110001101100000111;
            sine_reg0   <= 36'sb1001001100011111001101001100101010;
        end
        1859: begin
            cosine_reg0 <= 36'sb100001010101011110001001100100010100;
            sine_reg0   <= 36'sb1001001001011110100101000101110110;
        end
        1860: begin
            cosine_reg0 <= 36'sb100001010100100100110100010111000111;
            sine_reg0   <= 36'sb1001000110011101110111010101111000;
        end
        1861: begin
            cosine_reg0 <= 36'sb100001010011101011110010000101000011;
            sine_reg0   <= 36'sb1001000011011101000011111110100111;
        end
        1862: begin
            cosine_reg0 <= 36'sb100001010010110011000010101110101010;
            sine_reg0   <= 36'sb1001000000011100001011000001111011;
        end
        1863: begin
            cosine_reg0 <= 36'sb100001010001111010100110010100100001;
            sine_reg0   <= 36'sb1000111101011011001100100001101001;
        end
        1864: begin
            cosine_reg0 <= 36'sb100001010001000010011100110111001001;
            sine_reg0   <= 36'sb1000111010011010001000011111101001;
        end
        1865: begin
            cosine_reg0 <= 36'sb100001010000001010100110010111000110;
            sine_reg0   <= 36'sb1000110111011000111110111101110011;
        end
        1866: begin
            cosine_reg0 <= 36'sb100001001111010011000010110100111010;
            sine_reg0   <= 36'sb1000110100010111101111111101111101;
        end
        1867: begin
            cosine_reg0 <= 36'sb100001001110011011110010010001000111;
            sine_reg0   <= 36'sb1000110001010110011011100001111110;
        end
        1868: begin
            cosine_reg0 <= 36'sb100001001101100100110100101100010000;
            sine_reg0   <= 36'sb1000101110010101000001101011101111;
        end
        1869: begin
            cosine_reg0 <= 36'sb100001001100101110001010000110110110;
            sine_reg0   <= 36'sb1000101011010011100010011101000101;
        end
        1870: begin
            cosine_reg0 <= 36'sb100001001011110111110010100001011011;
            sine_reg0   <= 36'sb1000101000010001111101110111111001;
        end
        1871: begin
            cosine_reg0 <= 36'sb100001001011000001101101111100100000;
            sine_reg0   <= 36'sb1000100101010000010011111110000001;
        end
        1872: begin
            cosine_reg0 <= 36'sb100001001010001011111100011000100111;
            sine_reg0   <= 36'sb1000100010001110100100110001010110;
        end
        1873: begin
            cosine_reg0 <= 36'sb100001001001010110011101110110010001;
            sine_reg0   <= 36'sb1000011111001100110000010011101111;
        end
        1874: begin
            cosine_reg0 <= 36'sb100001001000100001010010010101111111;
            sine_reg0   <= 36'sb1000011100001010110110100111000011;
        end
        1875: begin
            cosine_reg0 <= 36'sb100001000111101100011001111000010010;
            sine_reg0   <= 36'sb1000011001001000110111101101001010;
        end
        1876: begin
            cosine_reg0 <= 36'sb100001000110110111110100011101101010;
            sine_reg0   <= 36'sb1000010110000110110011100111111011;
        end
        1877: begin
            cosine_reg0 <= 36'sb100001000110000011100010000110101001;
            sine_reg0   <= 36'sb1000010011000100101010011001001111;
        end
        1878: begin
            cosine_reg0 <= 36'sb100001000101001111100010110011101101;
            sine_reg0   <= 36'sb1000010000000010011100000010111101;
        end
        1879: begin
            cosine_reg0 <= 36'sb100001000100011011110110100101010111;
            sine_reg0   <= 36'sb1000001101000000001000100110111101;
        end
        1880: begin
            cosine_reg0 <= 36'sb100001000011101000011101011100001000;
            sine_reg0   <= 36'sb1000001001111101110000000111000111;
        end
        1881: begin
            cosine_reg0 <= 36'sb100001000010110101010111011000011110;
            sine_reg0   <= 36'sb1000000110111011010010100101010010;
        end
        1882: begin
            cosine_reg0 <= 36'sb100001000010000010100100011010111010;
            sine_reg0   <= 36'sb1000000011111000110000000011010111;
        end
        1883: begin
            cosine_reg0 <= 36'sb100001000001010000000100100011111010;
            sine_reg0   <= 36'sb1000000000110110001000100011001110;
        end
        1884: begin
            cosine_reg0 <= 36'sb100001000000011101110111110011111110;
            sine_reg0   <= 36'sb111111101110011011100000110101110;
        end
        1885: begin
            cosine_reg0 <= 36'sb100000111111101011111110001011100101;
            sine_reg0   <= 36'sb111111010110000101010101111110000;
        end
        1886: begin
            cosine_reg0 <= 36'sb100000111110111010010111101011001101;
            sine_reg0   <= 36'sb111110111101101110100100000001100;
        end
        1887: begin
            cosine_reg0 <= 36'sb100000111110001001000100010011010101;
            sine_reg0   <= 36'sb111110100101010111001011001111010;
        end
        1888: begin
            cosine_reg0 <= 36'sb100000111101011000000100000100011100;
            sine_reg0   <= 36'sb111110001100111111001011110110010;
        end
        1889: begin
            cosine_reg0 <= 36'sb100000111100100111010110111111000000;
            sine_reg0   <= 36'sb111101110100100110100110000101101;
        end
        1890: begin
            cosine_reg0 <= 36'sb100000111011110110111101000011011111;
            sine_reg0   <= 36'sb111101011100001101011010001100011;
        end
        1891: begin
            cosine_reg0 <= 36'sb100000111011000110110110010010010110;
            sine_reg0   <= 36'sb111101000011110011101000011001100;
        end
        1892: begin
            cosine_reg0 <= 36'sb100000111010010111000010101100000011;
            sine_reg0   <= 36'sb111100101011011001010000111100001;
        end
        1893: begin
            cosine_reg0 <= 36'sb100000111001100111100010010001000100;
            sine_reg0   <= 36'sb111100010010111110010100000011010;
        end
        1894: begin
            cosine_reg0 <= 36'sb100000111000111000010101000001110111;
            sine_reg0   <= 36'sb111011111010100010110001111110000;
        end
        1895: begin
            cosine_reg0 <= 36'sb100000111000001001011010111110111000;
            sine_reg0   <= 36'sb111011100010000110101010111011011;
        end
        1896: begin
            cosine_reg0 <= 36'sb100000110111011010110100001000100011;
            sine_reg0   <= 36'sb111011001001101001111111001010100;
        end
        1897: begin
            cosine_reg0 <= 36'sb100000110110101100100000011111010111;
            sine_reg0   <= 36'sb111010110001001100101110111010100;
        end
        1898: begin
            cosine_reg0 <= 36'sb100000110101111110100000000011101111;
            sine_reg0   <= 36'sb111010011000101110111010011010011;
        end
        1899: begin
            cosine_reg0 <= 36'sb100000110101010000110010110110001001;
            sine_reg0   <= 36'sb111010000000010000100001111001001;
        end
        1900: begin
            cosine_reg0 <= 36'sb100000110100100011011000110110111111;
            sine_reg0   <= 36'sb111001100111110001100101100110001;
        end
        1901: begin
            cosine_reg0 <= 36'sb100000110011110110010010000110101110;
            sine_reg0   <= 36'sb111001001111010010000101110000010;
        end
        1902: begin
            cosine_reg0 <= 36'sb100000110011001001011110100101110010;
            sine_reg0   <= 36'sb111000110110110010000010100110110;
        end
        1903: begin
            cosine_reg0 <= 36'sb100000110010011100111110010100100111;
            sine_reg0   <= 36'sb111000011110010001011100011000101;
        end
        1904: begin
            cosine_reg0 <= 36'sb100000110001110000110001010011101000;
            sine_reg0   <= 36'sb111000000101110000010011010101000;
        end
        1905: begin
            cosine_reg0 <= 36'sb100000110001000100110111100011010000;
            sine_reg0   <= 36'sb110111101101001110100111101011000;
        end
        1906: begin
            cosine_reg0 <= 36'sb100000110000011001010001000011111010;
            sine_reg0   <= 36'sb110111010100101100011001101001111;
        end
        1907: begin
            cosine_reg0 <= 36'sb100000101111101101111101110110000010;
            sine_reg0   <= 36'sb110110111100001001101001100000101;
        end
        1908: begin
            cosine_reg0 <= 36'sb100000101111000010111101111010000001;
            sine_reg0   <= 36'sb110110100011100110010111011110100;
        end
        1909: begin
            cosine_reg0 <= 36'sb100000101110011000010001010000010011;
            sine_reg0   <= 36'sb110110001011000010100011110010100;
        end
        1910: begin
            cosine_reg0 <= 36'sb100000101101101101110111111001010010;
            sine_reg0   <= 36'sb110101110010011110001110101011111;
        end
        1911: begin
            cosine_reg0 <= 36'sb100000101101000011110001110101011000;
            sine_reg0   <= 36'sb110101011001111001011000011001110;
        end
        1912: begin
            cosine_reg0 <= 36'sb100000101100011001111111000100111110;
            sine_reg0   <= 36'sb110101000001010100000001001011011;
        end
        1913: begin
            cosine_reg0 <= 36'sb100000101011110000011111101000100000;
            sine_reg0   <= 36'sb110100101000101110001001001111110;
        end
        1914: begin
            cosine_reg0 <= 36'sb100000101011000111010011100000010101;
            sine_reg0   <= 36'sb110100010000000111110000110110001;
        end
        1915: begin
            cosine_reg0 <= 36'sb100000101010011110011010101100111001;
            sine_reg0   <= 36'sb110011110111100000111000001101110;
        end
        1916: begin
            cosine_reg0 <= 36'sb100000101001110101110101001110100011;
            sine_reg0   <= 36'sb110011011110111001011111100101110;
        end
        1917: begin
            cosine_reg0 <= 36'sb100000101001001101100011000101101101;
            sine_reg0   <= 36'sb110011000110010001100111001101001;
        end
        1918: begin
            cosine_reg0 <= 36'sb100000101000100101100100010010110000;
            sine_reg0   <= 36'sb110010101101101001001111010011011;
        end
        1919: begin
            cosine_reg0 <= 36'sb100000100111111101111000110110000101;
            sine_reg0   <= 36'sb110010010101000000011000000111100;
        end
        1920: begin
            cosine_reg0 <= 36'sb100000100111010110100000110000000011;
            sine_reg0   <= 36'sb110001111100010111000001111000110;
        end
        1921: begin
            cosine_reg0 <= 36'sb100000100110101111011100000001000100;
            sine_reg0   <= 36'sb110001100011101101001100110110011;
        end
        1922: begin
            cosine_reg0 <= 36'sb100000100110001000101010101001011111;
            sine_reg0   <= 36'sb110001001011000010111001001111100;
        end
        1923: begin
            cosine_reg0 <= 36'sb100000100101100010001100101001101100;
            sine_reg0   <= 36'sb110000110010011000000111010011011;
        end
        1924: begin
            cosine_reg0 <= 36'sb100000100100111100000010000010000100;
            sine_reg0   <= 36'sb110000011001101100110111010001010;
        end
        1925: begin
            cosine_reg0 <= 36'sb100000100100010110001010110010111100;
            sine_reg0   <= 36'sb110000000001000001001001011000010;
        end
        1926: begin
            cosine_reg0 <= 36'sb100000100011110000100110111100101110;
            sine_reg0   <= 36'sb101111101000010100111101110111101;
        end
        1927: begin
            cosine_reg0 <= 36'sb100000100011001011010110011111110000;
            sine_reg0   <= 36'sb101111001111101000010100111110101;
        end
        1928: begin
            cosine_reg0 <= 36'sb100000100010100110011001011100011001;
            sine_reg0   <= 36'sb101110110110111011001110111100101;
        end
        1929: begin
            cosine_reg0 <= 36'sb100000100010000001101111110010111111;
            sine_reg0   <= 36'sb101110011110001101101100000000101;
        end
        1930: begin
            cosine_reg0 <= 36'sb100000100001011101011001100011111010;
            sine_reg0   <= 36'sb101110000101011111101100011010000;
        end
        1931: begin
            cosine_reg0 <= 36'sb100000100000111001010110101111100000;
            sine_reg0   <= 36'sb101101101100110001010000011000000;
        end
        1932: begin
            cosine_reg0 <= 36'sb100000100000010101100111010110000111;
            sine_reg0   <= 36'sb101101010100000010011000001001111;
        end
        1933: begin
            cosine_reg0 <= 36'sb100000011111110010001011011000000110;
            sine_reg0   <= 36'sb101100111011010011000011111110111;
        end
        1934: begin
            cosine_reg0 <= 36'sb100000011111001111000010110101110001;
            sine_reg0   <= 36'sb101100100010100011010100000110010;
        end
        1935: begin
            cosine_reg0 <= 36'sb100000011110101100001101101111011111;
            sine_reg0   <= 36'sb101100001001110011001000101111001;
        end
        1936: begin
            cosine_reg0 <= 36'sb100000011110001001101100000101100101;
            sine_reg0   <= 36'sb101011110001000010100010001001001;
        end
        1937: begin
            cosine_reg0 <= 36'sb100000011101100111011101111000011000;
            sine_reg0   <= 36'sb101011011000010001100000100011001;
        end
        1938: begin
            cosine_reg0 <= 36'sb100000011101000101100011001000001110;
            sine_reg0   <= 36'sb101010111111100000000100001100101;
        end
        1939: begin
            cosine_reg0 <= 36'sb100000011100100011111011110101011100;
            sine_reg0   <= 36'sb101010100110101110001101010100111;
        end
        1940: begin
            cosine_reg0 <= 36'sb100000011100000010101000000000010101;
            sine_reg0   <= 36'sb101010001101111011111100001011001;
        end
        1941: begin
            cosine_reg0 <= 36'sb100000011011100001100111101001010000;
            sine_reg0   <= 36'sb101001110101001001010000111110110;
        end
        1942: begin
            cosine_reg0 <= 36'sb100000011011000000111010110000100000;
            sine_reg0   <= 36'sb101001011100010110001011111110111;
        end
        1943: begin
            cosine_reg0 <= 36'sb100000011010100000100001010110011001;
            sine_reg0   <= 36'sb101001000011100010101101011011000;
        end
        1944: begin
            cosine_reg0 <= 36'sb100000011010000000011011011011001111;
            sine_reg0   <= 36'sb101000101010101110110101100010010;
        end
        1945: begin
            cosine_reg0 <= 36'sb100000011001100000101000111111010110;
            sine_reg0   <= 36'sb101000010001111010100100100100001;
        end
        1946: begin
            cosine_reg0 <= 36'sb100000011001000001001010000011000010;
            sine_reg0   <= 36'sb100111111001000101111010101111110;
        end
        1947: begin
            cosine_reg0 <= 36'sb100000011000100001111110100110100110;
            sine_reg0   <= 36'sb100111100000010000111000010100011;
        end
        1948: begin
            cosine_reg0 <= 36'sb100000011000000011000110101010010110;
            sine_reg0   <= 36'sb100111000111011011011101100001101;
        end
        1949: begin
            cosine_reg0 <= 36'sb100000010111100100100010001110100011;
            sine_reg0   <= 36'sb100110101110100101101010100110100;
        end
        1950: begin
            cosine_reg0 <= 36'sb100000010111000110010001010011100010;
            sine_reg0   <= 36'sb100110010101101111011111110010100;
        end
        1951: begin
            cosine_reg0 <= 36'sb100000010110101000010011111001100101;
            sine_reg0   <= 36'sb100101111100111000111101010101000;
        end
        1952: begin
            cosine_reg0 <= 36'sb100000010110001010101010000000111111;
            sine_reg0   <= 36'sb100101100100000010000011011101001;
        end
        1953: begin
            cosine_reg0 <= 36'sb100000010101101101010011101010000001;
            sine_reg0   <= 36'sb100101001011001010110010011010011;
        end
        1954: begin
            cosine_reg0 <= 36'sb100000010101010000010000110100111110;
            sine_reg0   <= 36'sb100100110010010011001010011100000;
        end
        1955: begin
            cosine_reg0 <= 36'sb100000010100110011100001100010000111;
            sine_reg0   <= 36'sb100100011001011011001011110001011;
        end
        1956: begin
            cosine_reg0 <= 36'sb100000010100010111000101110001101111;
            sine_reg0   <= 36'sb100100000000100010110110101001111;
        end
        1957: begin
            cosine_reg0 <= 36'sb100000010011111010111101100100000111;
            sine_reg0   <= 36'sb100011100111101010001011010100110;
        end
        1958: begin
            cosine_reg0 <= 36'sb100000010011011111001000111001100001;
            sine_reg0   <= 36'sb100011001110110001001010000001100;
        end
        1959: begin
            cosine_reg0 <= 36'sb100000010011000011100111110010001100;
            sine_reg0   <= 36'sb100010110101110111110010111111011;
        end
        1960: begin
            cosine_reg0 <= 36'sb100000010010101000011010001110011100;
            sine_reg0   <= 36'sb100010011100111110000110011101110;
        end
        1961: begin
            cosine_reg0 <= 36'sb100000010010001101100000001110011111;
            sine_reg0   <= 36'sb100010000100000100000100101011111;
        end
        1962: begin
            cosine_reg0 <= 36'sb100000010001110010111001110010100111;
            sine_reg0   <= 36'sb100001101011001001101101111001011;
        end
        1963: begin
            cosine_reg0 <= 36'sb100000010001011000100110111011000101;
            sine_reg0   <= 36'sb100001010010001111000010010101011;
        end
        1964: begin
            cosine_reg0 <= 36'sb100000010000111110100111101000001000;
            sine_reg0   <= 36'sb100000111001010100000010001111100;
        end
        1965: begin
            cosine_reg0 <= 36'sb100000010000100100111011111010000000;
            sine_reg0   <= 36'sb100000100000011000101101110110110;
        end
        1966: begin
            cosine_reg0 <= 36'sb100000010000001011100011110000111110;
            sine_reg0   <= 36'sb100000000111011101000101011010111;
        end
        1967: begin
            cosine_reg0 <= 36'sb100000001111110010011111001101010001;
            sine_reg0   <= 36'sb11111101110100001001001001011000;
        end
        1968: begin
            cosine_reg0 <= 36'sb100000001111011001101110001111001001;
            sine_reg0   <= 36'sb11111010101100100111001010110101;
        end
        1969: begin
            cosine_reg0 <= 36'sb100000001111000001010000110110110100;
            sine_reg0   <= 36'sb11110111100101000010110001101001;
        end
        1970: begin
            cosine_reg0 <= 36'sb100000001110101001000111000100100010;
            sine_reg0   <= 36'sb11110100011101011011111111101111;
        end
        1971: begin
            cosine_reg0 <= 36'sb100000001110010001010000111000100001;
            sine_reg0   <= 36'sb11110001010101110010110111000010;
        end
        1972: begin
            cosine_reg0 <= 36'sb100000001101111001101110010011000001;
            sine_reg0   <= 36'sb11101110001110000111011001011101;
        end
        1973: begin
            cosine_reg0 <= 36'sb100000001101100010011111010100010000;
            sine_reg0   <= 36'sb11101011000110011001101000111100;
        end
        1974: begin
            cosine_reg0 <= 36'sb100000001101001011100011111100011101;
            sine_reg0   <= 36'sb11100111111110101001100111011001;
        end
        1975: begin
            cosine_reg0 <= 36'sb100000001100110100111100001011110100;
            sine_reg0   <= 36'sb11100100110110110111010110110001;
        end
        1976: begin
            cosine_reg0 <= 36'sb100000001100011110101000000010100110;
            sine_reg0   <= 36'sb11100001101111000010111000111101;
        end
        1977: begin
            cosine_reg0 <= 36'sb100000001100001000100111100000111110;
            sine_reg0   <= 36'sb11011110100111001100001111111001;
        end
        1978: begin
            cosine_reg0 <= 36'sb100000001011110010111010100111001011;
            sine_reg0   <= 36'sb11011011011111010011011101100010;
        end
        1979: begin
            cosine_reg0 <= 36'sb100000001011011101100001010101011010;
            sine_reg0   <= 36'sb11011000010111011000100011110001;
        end
        1980: begin
            cosine_reg0 <= 36'sb100000001011001000011011101011111000;
            sine_reg0   <= 36'sb11010101001111011011100100100010;
        end
        1981: begin
            cosine_reg0 <= 36'sb100000001010110011101001101010110011;
            sine_reg0   <= 36'sb11010010000111011100100001110001;
        end
        1982: begin
            cosine_reg0 <= 36'sb100000001010011111001011010010010111;
            sine_reg0   <= 36'sb11001110111111011011011101011001;
        end
        1983: begin
            cosine_reg0 <= 36'sb100000001010001011000000100010110001;
            sine_reg0   <= 36'sb11001011110111011000011001010101;
        end
        1984: begin
            cosine_reg0 <= 36'sb100000001001110111001001011100001101;
            sine_reg0   <= 36'sb11001000101111010011010111100001;
        end
        1985: begin
            cosine_reg0 <= 36'sb100000001001100011100101111110110111;
            sine_reg0   <= 36'sb11000101100111001100011001111000;
        end
        1986: begin
            cosine_reg0 <= 36'sb100000001001010000010110001010111100;
            sine_reg0   <= 36'sb11000010011111000011100010010110;
        end
        1987: begin
            cosine_reg0 <= 36'sb100000001000111101011010000000100111;
            sine_reg0   <= 36'sb10111111010110111000110010110110;
        end
        1988: begin
            cosine_reg0 <= 36'sb100000001000101010110001100000000101;
            sine_reg0   <= 36'sb10111100001110101100001101010011;
        end
        1989: begin
            cosine_reg0 <= 36'sb100000001000011000011100101001011111;
            sine_reg0   <= 36'sb10111001000110011101110011101001;
        end
        1990: begin
            cosine_reg0 <= 36'sb100000001000000110011011011101000011;
            sine_reg0   <= 36'sb10110101111110001101100111110100;
        end
        1991: begin
            cosine_reg0 <= 36'sb100000000111110100101101111010111011;
            sine_reg0   <= 36'sb10110010110101111011101011101110;
        end
        1992: begin
            cosine_reg0 <= 36'sb100000000111100011010100000011010010;
            sine_reg0   <= 36'sb10101111101101101000000001010101;
        end
        1993: begin
            cosine_reg0 <= 36'sb100000000111010010001101110110010010;
            sine_reg0   <= 36'sb10101100100101010010101010100010;
        end
        1994: begin
            cosine_reg0 <= 36'sb100000000111000001011011010100000111;
            sine_reg0   <= 36'sb10101001011100111011101001010010;
        end
        1995: begin
            cosine_reg0 <= 36'sb100000000110110000111100011100111010;
            sine_reg0   <= 36'sb10100110010100100010111111100001;
        end
        1996: begin
            cosine_reg0 <= 36'sb100000000110100000110001010000110101;
            sine_reg0   <= 36'sb10100011001100001000101111001001;
        end
        1997: begin
            cosine_reg0 <= 36'sb100000000110010000111001110000000100;
            sine_reg0   <= 36'sb10100000000011101100111010000111;
        end
        1998: begin
            cosine_reg0 <= 36'sb100000000110000001010101111010101111;
            sine_reg0   <= 36'sb10011100111011001111100010010110;
        end
        1999: begin
            cosine_reg0 <= 36'sb100000000101110010000101110001000000;
            sine_reg0   <= 36'sb10011001110010110000101001110010;
        end
        2000: begin
            cosine_reg0 <= 36'sb100000000101100011001001010011000001;
            sine_reg0   <= 36'sb10010110101010010000010010010110;
        end
        2001: begin
            cosine_reg0 <= 36'sb100000000101010100100000100000111010;
            sine_reg0   <= 36'sb10010011100001101110011101111111;
        end
        2002: begin
            cosine_reg0 <= 36'sb100000000101000110001011011010110101;
            sine_reg0   <= 36'sb10010000011001001011001110100111;
        end
        2003: begin
            cosine_reg0 <= 36'sb100000000100111000001010000000111011;
            sine_reg0   <= 36'sb10001101010000100110100110001011;
        end
        2004: begin
            cosine_reg0 <= 36'sb100000000100101010011100010011010011;
            sine_reg0   <= 36'sb10001010001000000000100110100111;
        end
        2005: begin
            cosine_reg0 <= 36'sb100000000100011101000010010010001000;
            sine_reg0   <= 36'sb10000110111111011001010001110101;
        end
        2006: begin
            cosine_reg0 <= 36'sb100000000100001111111011111101100000;
            sine_reg0   <= 36'sb10000011110110110000101001110010;
        end
        2007: begin
            cosine_reg0 <= 36'sb100000000100000011001001010101100101;
            sine_reg0   <= 36'sb10000000101110000110110000011010;
        end
        2008: begin
            cosine_reg0 <= 36'sb100000000011110110101010011010011101;
            sine_reg0   <= 36'sb1111101100101011011100111101000;
        end
        2009: begin
            cosine_reg0 <= 36'sb100000000011101010011111001100010001;
            sine_reg0   <= 36'sb1111010011100101111010001011000;
        end
        2010: begin
            cosine_reg0 <= 36'sb100000000011011110100111101011001001;
            sine_reg0   <= 36'sb1110111010100000001101111100110;
        end
        2011: begin
            cosine_reg0 <= 36'sb100000000011010011000011110111001010;
            sine_reg0   <= 36'sb1110100001011010011000100001110;
        end
        2012: begin
            cosine_reg0 <= 36'sb100000000011000111110011110000011110;
            sine_reg0   <= 36'sb1110001000010100011010001001011;
        end
        2013: begin
            cosine_reg0 <= 36'sb100000000010111100110111010111001001;
            sine_reg0   <= 36'sb1101101111001110010011000011010;
        end
        2014: begin
            cosine_reg0 <= 36'sb100000000010110010001110101011010101;
            sine_reg0   <= 36'sb1101010110001000000011011110101;
        end
        2015: begin
            cosine_reg0 <= 36'sb100000000010100111111001101101000101;
            sine_reg0   <= 36'sb1100111101000001101011101011010;
        end
        2016: begin
            cosine_reg0 <= 36'sb100000000010011101111000011100100011;
            sine_reg0   <= 36'sb1100100011111011001011111000100;
        end
        2017: begin
            cosine_reg0 <= 36'sb100000000010010100001010111001110010;
            sine_reg0   <= 36'sb1100001010110100100100010101111;
        end
        2018: begin
            cosine_reg0 <= 36'sb100000000010001010110001000100111010;
            sine_reg0   <= 36'sb1011110001101101110101010010110;
        end
        2019: begin
            cosine_reg0 <= 36'sb100000000010000001101010111110000000;
            sine_reg0   <= 36'sb1011011000100110111110111110110;
        end
        2020: begin
            cosine_reg0 <= 36'sb100000000001111000111000100101001010;
            sine_reg0   <= 36'sb1010111111100000000001101001010;
        end
        2021: begin
            cosine_reg0 <= 36'sb100000000001110000011001111010011101;
            sine_reg0   <= 36'sb1010100110011000111101100001111;
        end
        2022: begin
            cosine_reg0 <= 36'sb100000000001101000001110111101111111;
            sine_reg0   <= 36'sb1010001101010001110010111000000;
        end
        2023: begin
            cosine_reg0 <= 36'sb100000000001100000010111101111110100;
            sine_reg0   <= 36'sb1001110100001010100001111011001;
        end
        2024: begin
            cosine_reg0 <= 36'sb100000000001011000110100010000000001;
            sine_reg0   <= 36'sb1001011011000011001010111010110;
        end
        2025: begin
            cosine_reg0 <= 36'sb100000000001010001100100011110101100;
            sine_reg0   <= 36'sb1001000001111011101110000110100;
        end
        2026: begin
            cosine_reg0 <= 36'sb100000000001001010101000011011111000;
            sine_reg0   <= 36'sb1000101000110100001011101101101;
        end
        2027: begin
            cosine_reg0 <= 36'sb100000000001000100000000000111101001;
            sine_reg0   <= 36'sb1000001111101100100011111111110;
        end
        2028: begin
            cosine_reg0 <= 36'sb100000000000111101101011100010000101;
            sine_reg0   <= 36'sb111110110100100110111001100100;
        end
        2029: begin
            cosine_reg0 <= 36'sb100000000000110111101010101011001110;
            sine_reg0   <= 36'sb111011101011101000101100011001;
        end
        2030: begin
            cosine_reg0 <= 36'sb100000000000110001111101100011001000;
            sine_reg0   <= 36'sb111000100010101001111010011010;
        end
        2031: begin
            cosine_reg0 <= 36'sb100000000000101100100100001001111000;
            sine_reg0   <= 36'sb110101011001101010100101100011;
        end
        2032: begin
            cosine_reg0 <= 36'sb100000000000100111011110011111100000;
            sine_reg0   <= 36'sb110010010000101010101111101111;
        end
        2033: begin
            cosine_reg0 <= 36'sb100000000000100010101100100100000011;
            sine_reg0   <= 36'sb101111000111101010011010111100;
        end
        2034: begin
            cosine_reg0 <= 36'sb100000000000011110001110010111100101;
            sine_reg0   <= 36'sb101011111110101001101001000100;
        end
        2035: begin
            cosine_reg0 <= 36'sb100000000000011010000011111010001000;
            sine_reg0   <= 36'sb101000110101101000011100000100;
        end
        2036: begin
            cosine_reg0 <= 36'sb100000000000010110001101001011101110;
            sine_reg0   <= 36'sb100101101100100110110101111000;
        end
        2037: begin
            cosine_reg0 <= 36'sb100000000000010010101010001100011011;
            sine_reg0   <= 36'sb100010100011100100111000011011;
        end
        2038: begin
            cosine_reg0 <= 36'sb100000000000001111011010111100010000;
            sine_reg0   <= 36'sb11111011010100010100101101011;
        end
        2039: begin
            cosine_reg0 <= 36'sb100000000000001100011111011011001111;
            sine_reg0   <= 36'sb11100010001011111111111100010;
        end
        2040: begin
            cosine_reg0 <= 36'sb100000000000001001110111101001011010;
            sine_reg0   <= 36'sb11001001000011101000111111101;
        end
        2041: begin
            cosine_reg0 <= 36'sb100000000000000111100011100110110011;
            sine_reg0   <= 36'sb10101111111011010000000111000;
        end
        2042: begin
            cosine_reg0 <= 36'sb100000000000000101100011010011011011;
            sine_reg0   <= 36'sb10010110110010110101100001110;
        end
        2043: begin
            cosine_reg0 <= 36'sb100000000000000011110110101111010100;
            sine_reg0   <= 36'sb1111101101010011001011111101;
        end
        2044: begin
            cosine_reg0 <= 36'sb100000000000000010011101111010011101;
            sine_reg0   <= 36'sb1100100100001111100001111111;
        end
        2045: begin
            cosine_reg0 <= 36'sb100000000000000001011000110100111001;
            sine_reg0   <= 36'sb1001011011001011110000010001;
        end
        2046: begin
            cosine_reg0 <= 36'sb100000000000000000100111011110101000;
            sine_reg0   <= 36'sb110010010000111111000110000;
        end
        2047: begin
            cosine_reg0 <= 36'sb100000000000000000001001110111101011;
            sine_reg0   <= 36'sb11001001000011111101010110;
        end
        2048: begin
            cosine_reg0 <= 36'sb100000000000000000000000000000000001;
            sine_reg0   <= 36'sb0;
        end
        2049: begin
            cosine_reg0 <= 36'sb100000000000000000001001110111101011;
            sine_reg0   <= 36'sb111111111100110110111100000010101010;
        end
        2050: begin
            cosine_reg0 <= 36'sb100000000000000000100111011110101000;
            sine_reg0   <= 36'sb111111111001101101111000000111010000;
        end
        2051: begin
            cosine_reg0 <= 36'sb100000000000000001011000110100111001;
            sine_reg0   <= 36'sb111111110110100100110100001111101111;
        end
        2052: begin
            cosine_reg0 <= 36'sb100000000000000010011101111010011101;
            sine_reg0   <= 36'sb111111110011011011110000011110000001;
        end
        2053: begin
            cosine_reg0 <= 36'sb100000000000000011110110101111010100;
            sine_reg0   <= 36'sb111111110000010010101100110100000011;
        end
        2054: begin
            cosine_reg0 <= 36'sb100000000000000101100011010011011011;
            sine_reg0   <= 36'sb111111101101001001101001010011110010;
        end
        2055: begin
            cosine_reg0 <= 36'sb100000000000000111100011100110110011;
            sine_reg0   <= 36'sb111111101010000000100101111111001000;
        end
        2056: begin
            cosine_reg0 <= 36'sb100000000000001001110111101001011010;
            sine_reg0   <= 36'sb111111100110110111100010111000000011;
        end
        2057: begin
            cosine_reg0 <= 36'sb100000000000001100011111011011001111;
            sine_reg0   <= 36'sb111111100011101110100000000000011110;
        end
        2058: begin
            cosine_reg0 <= 36'sb100000000000001111011010111100010000;
            sine_reg0   <= 36'sb111111100000100101011101011010010101;
        end
        2059: begin
            cosine_reg0 <= 36'sb100000000000010010101010001100011011;
            sine_reg0   <= 36'sb111111011101011100011011000111100101;
        end
        2060: begin
            cosine_reg0 <= 36'sb100000000000010110001101001011101110;
            sine_reg0   <= 36'sb111111011010010011011001001010001000;
        end
        2061: begin
            cosine_reg0 <= 36'sb100000000000011010000011111010001000;
            sine_reg0   <= 36'sb111111010111001010010111100011111100;
        end
        2062: begin
            cosine_reg0 <= 36'sb100000000000011110001110010111100101;
            sine_reg0   <= 36'sb111111010100000001010110010110111100;
        end
        2063: begin
            cosine_reg0 <= 36'sb100000000000100010101100100100000011;
            sine_reg0   <= 36'sb111111010000111000010101100101000100;
        end
        2064: begin
            cosine_reg0 <= 36'sb100000000000100111011110011111100000;
            sine_reg0   <= 36'sb111111001101101111010101010000010001;
        end
        2065: begin
            cosine_reg0 <= 36'sb100000000000101100100100001001111000;
            sine_reg0   <= 36'sb111111001010100110010101011010011101;
        end
        2066: begin
            cosine_reg0 <= 36'sb100000000000110001111101100011001000;
            sine_reg0   <= 36'sb111111000111011101010110000101100110;
        end
        2067: begin
            cosine_reg0 <= 36'sb100000000000110111101010101011001110;
            sine_reg0   <= 36'sb111111000100010100010111010011100111;
        end
        2068: begin
            cosine_reg0 <= 36'sb100000000000111101101011100010000101;
            sine_reg0   <= 36'sb111111000001001011011001000110011100;
        end
        2069: begin
            cosine_reg0 <= 36'sb100000000001000100000000000111101001;
            sine_reg0   <= 36'sb111110111110000010011011100000000010;
        end
        2070: begin
            cosine_reg0 <= 36'sb100000000001001010101000011011111000;
            sine_reg0   <= 36'sb111110111010111001011110100010010011;
        end
        2071: begin
            cosine_reg0 <= 36'sb100000000001010001100100011110101100;
            sine_reg0   <= 36'sb111110110111110000100010001111001100;
        end
        2072: begin
            cosine_reg0 <= 36'sb100000000001011000110100010000000001;
            sine_reg0   <= 36'sb111110110100100111100110101000101010;
        end
        2073: begin
            cosine_reg0 <= 36'sb100000000001100000010111101111110100;
            sine_reg0   <= 36'sb111110110001011110101011110000100111;
        end
        2074: begin
            cosine_reg0 <= 36'sb100000000001101000001110111101111111;
            sine_reg0   <= 36'sb111110101110010101110001101001000000;
        end
        2075: begin
            cosine_reg0 <= 36'sb100000000001110000011001111010011101;
            sine_reg0   <= 36'sb111110101011001100111000010011110001;
        end
        2076: begin
            cosine_reg0 <= 36'sb100000000001111000111000100101001010;
            sine_reg0   <= 36'sb111110101000000011111111110010110110;
        end
        2077: begin
            cosine_reg0 <= 36'sb100000000010000001101010111110000000;
            sine_reg0   <= 36'sb111110100100111011001000001000001010;
        end
        2078: begin
            cosine_reg0 <= 36'sb100000000010001010110001000100111010;
            sine_reg0   <= 36'sb111110100001110010010001010101101010;
        end
        2079: begin
            cosine_reg0 <= 36'sb100000000010010100001010111001110010;
            sine_reg0   <= 36'sb111110011110101001011011011101010001;
        end
        2080: begin
            cosine_reg0 <= 36'sb100000000010011101111000011100100011;
            sine_reg0   <= 36'sb111110011011100000100110100000111100;
        end
        2081: begin
            cosine_reg0 <= 36'sb100000000010100111111001101101000101;
            sine_reg0   <= 36'sb111110011000010111110010100010100110;
        end
        2082: begin
            cosine_reg0 <= 36'sb100000000010110010001110101011010101;
            sine_reg0   <= 36'sb111110010101001110111111100100001011;
        end
        2083: begin
            cosine_reg0 <= 36'sb100000000010111100110111010111001001;
            sine_reg0   <= 36'sb111110010010000110001101100111100110;
        end
        2084: begin
            cosine_reg0 <= 36'sb100000000011000111110011110000011110;
            sine_reg0   <= 36'sb111110001110111101011100101110110101;
        end
        2085: begin
            cosine_reg0 <= 36'sb100000000011010011000011110111001010;
            sine_reg0   <= 36'sb111110001011110100101100111011110010;
        end
        2086: begin
            cosine_reg0 <= 36'sb100000000011011110100111101011001001;
            sine_reg0   <= 36'sb111110001000101011111110010000011010;
        end
        2087: begin
            cosine_reg0 <= 36'sb100000000011101010011111001100010001;
            sine_reg0   <= 36'sb111110000101100011010000101110101000;
        end
        2088: begin
            cosine_reg0 <= 36'sb100000000011110110101010011010011101;
            sine_reg0   <= 36'sb111110000010011010100100011000011000;
        end
        2089: begin
            cosine_reg0 <= 36'sb100000000100000011001001010101100101;
            sine_reg0   <= 36'sb111101111111010001111001001111100110;
        end
        2090: begin
            cosine_reg0 <= 36'sb100000000100001111111011111101100000;
            sine_reg0   <= 36'sb111101111100001001001111010110001110;
        end
        2091: begin
            cosine_reg0 <= 36'sb100000000100011101000010010010001000;
            sine_reg0   <= 36'sb111101111001000000100110101110001011;
        end
        2092: begin
            cosine_reg0 <= 36'sb100000000100101010011100010011010011;
            sine_reg0   <= 36'sb111101110101110111111111011001011001;
        end
        2093: begin
            cosine_reg0 <= 36'sb100000000100111000001010000000111011;
            sine_reg0   <= 36'sb111101110010101111011001011001110101;
        end
        2094: begin
            cosine_reg0 <= 36'sb100000000101000110001011011010110101;
            sine_reg0   <= 36'sb111101101111100110110100110001011001;
        end
        2095: begin
            cosine_reg0 <= 36'sb100000000101010100100000100000111010;
            sine_reg0   <= 36'sb111101101100011110010001100010000001;
        end
        2096: begin
            cosine_reg0 <= 36'sb100000000101100011001001010011000001;
            sine_reg0   <= 36'sb111101101001010101101111101101101010;
        end
        2097: begin
            cosine_reg0 <= 36'sb100000000101110010000101110001000000;
            sine_reg0   <= 36'sb111101100110001101001111010110001110;
        end
        2098: begin
            cosine_reg0 <= 36'sb100000000110000001010101111010101111;
            sine_reg0   <= 36'sb111101100011000100110000011101101010;
        end
        2099: begin
            cosine_reg0 <= 36'sb100000000110010000111001110000000100;
            sine_reg0   <= 36'sb111101011111111100010011000101111001;
        end
        2100: begin
            cosine_reg0 <= 36'sb100000000110100000110001010000110101;
            sine_reg0   <= 36'sb111101011100110011110111010000110111;
        end
        2101: begin
            cosine_reg0 <= 36'sb100000000110110000111100011100111010;
            sine_reg0   <= 36'sb111101011001101011011101000000011111;
        end
        2102: begin
            cosine_reg0 <= 36'sb100000000111000001011011010100000111;
            sine_reg0   <= 36'sb111101010110100011000100010110101110;
        end
        2103: begin
            cosine_reg0 <= 36'sb100000000111010010001101110110010010;
            sine_reg0   <= 36'sb111101010011011010101101010101011110;
        end
        2104: begin
            cosine_reg0 <= 36'sb100000000111100011010100000011010010;
            sine_reg0   <= 36'sb111101010000010010010111111110101011;
        end
        2105: begin
            cosine_reg0 <= 36'sb100000000111110100101101111010111011;
            sine_reg0   <= 36'sb111101001101001010000100010100010010;
        end
        2106: begin
            cosine_reg0 <= 36'sb100000001000000110011011011101000011;
            sine_reg0   <= 36'sb111101001010000001110010011000001100;
        end
        2107: begin
            cosine_reg0 <= 36'sb100000001000011000011100101001011111;
            sine_reg0   <= 36'sb111101000110111001100010001100010111;
        end
        2108: begin
            cosine_reg0 <= 36'sb100000001000101010110001100000000101;
            sine_reg0   <= 36'sb111101000011110001010011110010101101;
        end
        2109: begin
            cosine_reg0 <= 36'sb100000001000111101011010000000100111;
            sine_reg0   <= 36'sb111101000000101001000111001101001010;
        end
        2110: begin
            cosine_reg0 <= 36'sb100000001001010000010110001010111100;
            sine_reg0   <= 36'sb111100111101100000111100011101101010;
        end
        2111: begin
            cosine_reg0 <= 36'sb100000001001100011100101111110110111;
            sine_reg0   <= 36'sb111100111010011000110011100110001000;
        end
        2112: begin
            cosine_reg0 <= 36'sb100000001001110111001001011100001101;
            sine_reg0   <= 36'sb111100110111010000101100101000011111;
        end
        2113: begin
            cosine_reg0 <= 36'sb100000001010001011000000100010110001;
            sine_reg0   <= 36'sb111100110100001000100111100110101011;
        end
        2114: begin
            cosine_reg0 <= 36'sb100000001010011111001011010010010111;
            sine_reg0   <= 36'sb111100110001000000100100100010100111;
        end
        2115: begin
            cosine_reg0 <= 36'sb100000001010110011101001101010110011;
            sine_reg0   <= 36'sb111100101101111000100011011110001111;
        end
        2116: begin
            cosine_reg0 <= 36'sb100000001011001000011011101011111000;
            sine_reg0   <= 36'sb111100101010110000100100011011011110;
        end
        2117: begin
            cosine_reg0 <= 36'sb100000001011011101100001010101011010;
            sine_reg0   <= 36'sb111100100111101000100111011100001111;
        end
        2118: begin
            cosine_reg0 <= 36'sb100000001011110010111010100111001011;
            sine_reg0   <= 36'sb111100100100100000101100100010011110;
        end
        2119: begin
            cosine_reg0 <= 36'sb100000001100001000100111100000111110;
            sine_reg0   <= 36'sb111100100001011000110011110000000111;
        end
        2120: begin
            cosine_reg0 <= 36'sb100000001100011110101000000010100110;
            sine_reg0   <= 36'sb111100011110010000111101000111000011;
        end
        2121: begin
            cosine_reg0 <= 36'sb100000001100110100111100001011110100;
            sine_reg0   <= 36'sb111100011011001001001000101001001111;
        end
        2122: begin
            cosine_reg0 <= 36'sb100000001101001011100011111100011101;
            sine_reg0   <= 36'sb111100011000000001010110011000100111;
        end
        2123: begin
            cosine_reg0 <= 36'sb100000001101100010011111010100010000;
            sine_reg0   <= 36'sb111100010100111001100110010111000100;
        end
        2124: begin
            cosine_reg0 <= 36'sb100000001101111001101110010011000001;
            sine_reg0   <= 36'sb111100010001110001111000100110100011;
        end
        2125: begin
            cosine_reg0 <= 36'sb100000001110010001010000111000100001;
            sine_reg0   <= 36'sb111100001110101010001101001000111110;
        end
        2126: begin
            cosine_reg0 <= 36'sb100000001110101001000111000100100010;
            sine_reg0   <= 36'sb111100001011100010100100000000010001;
        end
        2127: begin
            cosine_reg0 <= 36'sb100000001111000001010000110110110100;
            sine_reg0   <= 36'sb111100001000011010111101001110010111;
        end
        2128: begin
            cosine_reg0 <= 36'sb100000001111011001101110001111001001;
            sine_reg0   <= 36'sb111100000101010011011000110101001011;
        end
        2129: begin
            cosine_reg0 <= 36'sb100000001111110010011111001101010001;
            sine_reg0   <= 36'sb111100000010001011110110110110101000;
        end
        2130: begin
            cosine_reg0 <= 36'sb100000010000001011100011110000111110;
            sine_reg0   <= 36'sb111011111111000100010111010100101001;
        end
        2131: begin
            cosine_reg0 <= 36'sb100000010000100100111011111010000000;
            sine_reg0   <= 36'sb111011111011111100111010010001001010;
        end
        2132: begin
            cosine_reg0 <= 36'sb100000010000111110100111101000001000;
            sine_reg0   <= 36'sb111011111000110101011111101110000100;
        end
        2133: begin
            cosine_reg0 <= 36'sb100000010001011000100110111011000101;
            sine_reg0   <= 36'sb111011110101101110000111101101010101;
        end
        2134: begin
            cosine_reg0 <= 36'sb100000010001110010111001110010100111;
            sine_reg0   <= 36'sb111011110010100110110010010000110101;
        end
        2135: begin
            cosine_reg0 <= 36'sb100000010010001101100000001110011111;
            sine_reg0   <= 36'sb111011101111011111011111011010100001;
        end
        2136: begin
            cosine_reg0 <= 36'sb100000010010101000011010001110011100;
            sine_reg0   <= 36'sb111011101100011000001111001100010010;
        end
        2137: begin
            cosine_reg0 <= 36'sb100000010011000011100111110010001100;
            sine_reg0   <= 36'sb111011101001010001000001101000000101;
        end
        2138: begin
            cosine_reg0 <= 36'sb100000010011011111001000111001100001;
            sine_reg0   <= 36'sb111011100110001001110110101111110100;
        end
        2139: begin
            cosine_reg0 <= 36'sb100000010011111010111101100100000111;
            sine_reg0   <= 36'sb111011100011000010101110100101011010;
        end
        2140: begin
            cosine_reg0 <= 36'sb100000010100010111000101110001101111;
            sine_reg0   <= 36'sb111011011111111011101001001010110001;
        end
        2141: begin
            cosine_reg0 <= 36'sb100000010100110011100001100010000111;
            sine_reg0   <= 36'sb111011011100110100100110100001110101;
        end
        2142: begin
            cosine_reg0 <= 36'sb100000010101010000010000110100111110;
            sine_reg0   <= 36'sb111011011001101101100110101100100000;
        end
        2143: begin
            cosine_reg0 <= 36'sb100000010101101101010011101010000001;
            sine_reg0   <= 36'sb111011010110100110101001101100101101;
        end
        2144: begin
            cosine_reg0 <= 36'sb100000010110001010101010000000111111;
            sine_reg0   <= 36'sb111011010011011111101111100100010111;
        end
        2145: begin
            cosine_reg0 <= 36'sb100000010110101000010011111001100101;
            sine_reg0   <= 36'sb111011010000011000111000010101011000;
        end
        2146: begin
            cosine_reg0 <= 36'sb100000010111000110010001010011100010;
            sine_reg0   <= 36'sb111011001101010010000100000001101100;
        end
        2147: begin
            cosine_reg0 <= 36'sb100000010111100100100010001110100011;
            sine_reg0   <= 36'sb111011001010001011010010101011001100;
        end
        2148: begin
            cosine_reg0 <= 36'sb100000011000000011000110101010010110;
            sine_reg0   <= 36'sb111011000111000100100100010011110011;
        end
        2149: begin
            cosine_reg0 <= 36'sb100000011000100001111110100110100110;
            sine_reg0   <= 36'sb111011000011111101111000111101011101;
        end
        2150: begin
            cosine_reg0 <= 36'sb100000011001000001001010000011000010;
            sine_reg0   <= 36'sb111011000000110111010000101010000010;
        end
        2151: begin
            cosine_reg0 <= 36'sb100000011001100000101000111111010110;
            sine_reg0   <= 36'sb111010111101110000101011011011011111;
        end
        2152: begin
            cosine_reg0 <= 36'sb100000011010000000011011011011001111;
            sine_reg0   <= 36'sb111010111010101010001001010011101110;
        end
        2153: begin
            cosine_reg0 <= 36'sb100000011010100000100001010110011001;
            sine_reg0   <= 36'sb111010110111100011101010010100101000;
        end
        2154: begin
            cosine_reg0 <= 36'sb100000011011000000111010110000100000;
            sine_reg0   <= 36'sb111010110100011101001110100000001001;
        end
        2155: begin
            cosine_reg0 <= 36'sb100000011011100001100111101001010000;
            sine_reg0   <= 36'sb111010110001010110110101111000001010;
        end
        2156: begin
            cosine_reg0 <= 36'sb100000011100000010101000000000010101;
            sine_reg0   <= 36'sb111010101110010000100000011110100111;
        end
        2157: begin
            cosine_reg0 <= 36'sb100000011100100011111011110101011100;
            sine_reg0   <= 36'sb111010101011001010001110010101011001;
        end
        2158: begin
            cosine_reg0 <= 36'sb100000011101000101100011001000001110;
            sine_reg0   <= 36'sb111010101000000011111111011110011011;
        end
        2159: begin
            cosine_reg0 <= 36'sb100000011101100111011101111000011000;
            sine_reg0   <= 36'sb111010100100111101110011111011100111;
        end
        2160: begin
            cosine_reg0 <= 36'sb100000011110001001101100000101100101;
            sine_reg0   <= 36'sb111010100001110111101011101110110111;
        end
        2161: begin
            cosine_reg0 <= 36'sb100000011110101100001101101111011111;
            sine_reg0   <= 36'sb111010011110110001100110111010000111;
        end
        2162: begin
            cosine_reg0 <= 36'sb100000011111001111000010110101110001;
            sine_reg0   <= 36'sb111010011011101011100101011111001110;
        end
        2163: begin
            cosine_reg0 <= 36'sb100000011111110010001011011000000110;
            sine_reg0   <= 36'sb111010011000100101100111100000001001;
        end
        2164: begin
            cosine_reg0 <= 36'sb100000100000010101100111010110000111;
            sine_reg0   <= 36'sb111010010101011111101100111110110001;
        end
        2165: begin
            cosine_reg0 <= 36'sb100000100000111001010110101111100000;
            sine_reg0   <= 36'sb111010010010011001110101111101000000;
        end
        2166: begin
            cosine_reg0 <= 36'sb100000100001011101011001100011111010;
            sine_reg0   <= 36'sb111010001111010100000010011100110000;
        end
        2167: begin
            cosine_reg0 <= 36'sb100000100010000001101111110010111111;
            sine_reg0   <= 36'sb111010001100001110010010011111111011;
        end
        2168: begin
            cosine_reg0 <= 36'sb100000100010100110011001011100011001;
            sine_reg0   <= 36'sb111010001001001000100110001000011011;
        end
        2169: begin
            cosine_reg0 <= 36'sb100000100011001011010110011111110000;
            sine_reg0   <= 36'sb111010000110000010111101011000001011;
        end
        2170: begin
            cosine_reg0 <= 36'sb100000100011110000100110111100101110;
            sine_reg0   <= 36'sb111010000010111101011000010001000011;
        end
        2171: begin
            cosine_reg0 <= 36'sb100000100100010110001010110010111100;
            sine_reg0   <= 36'sb111001111111110111110110110100111110;
        end
        2172: begin
            cosine_reg0 <= 36'sb100000100100111100000010000010000100;
            sine_reg0   <= 36'sb111001111100110010011001000101110110;
        end
        2173: begin
            cosine_reg0 <= 36'sb100000100101100010001100101001101100;
            sine_reg0   <= 36'sb111001111001101100111111000101100101;
        end
        2174: begin
            cosine_reg0 <= 36'sb100000100110001000101010101001011111;
            sine_reg0   <= 36'sb111001110110100111101000110110000100;
        end
        2175: begin
            cosine_reg0 <= 36'sb100000100110101111011100000001000100;
            sine_reg0   <= 36'sb111001110011100010010110011001001101;
        end
        2176: begin
            cosine_reg0 <= 36'sb100000100111010110100000110000000011;
            sine_reg0   <= 36'sb111001110000011101000111110000111010;
        end
        2177: begin
            cosine_reg0 <= 36'sb100000100111111101111000110110000101;
            sine_reg0   <= 36'sb111001101101010111111100111111000100;
        end
        2178: begin
            cosine_reg0 <= 36'sb100000101000100101100100010010110000;
            sine_reg0   <= 36'sb111001101010010010110110000101100101;
        end
        2179: begin
            cosine_reg0 <= 36'sb100000101001001101100011000101101101;
            sine_reg0   <= 36'sb111001100111001101110011000110010111;
        end
        2180: begin
            cosine_reg0 <= 36'sb100000101001110101110101001110100011;
            sine_reg0   <= 36'sb111001100100001000110100000011010010;
        end
        2181: begin
            cosine_reg0 <= 36'sb100000101010011110011010101100111001;
            sine_reg0   <= 36'sb111001100001000011111000111110010010;
        end
        2182: begin
            cosine_reg0 <= 36'sb100000101011000111010011100000010101;
            sine_reg0   <= 36'sb111001011101111111000001111001001111;
        end
        2183: begin
            cosine_reg0 <= 36'sb100000101011110000011111101000100000;
            sine_reg0   <= 36'sb111001011010111010001110110110000010;
        end
        2184: begin
            cosine_reg0 <= 36'sb100000101100011001111111000100111110;
            sine_reg0   <= 36'sb111001010111110101011111110110100101;
        end
        2185: begin
            cosine_reg0 <= 36'sb100000101101000011110001110101011000;
            sine_reg0   <= 36'sb111001010100110000110100111100110010;
        end
        2186: begin
            cosine_reg0 <= 36'sb100000101101101101110111111001010010;
            sine_reg0   <= 36'sb111001010001101100001110001010100001;
        end
        2187: begin
            cosine_reg0 <= 36'sb100000101110011000010001010000010011;
            sine_reg0   <= 36'sb111001001110100111101011100001101100;
        end
        2188: begin
            cosine_reg0 <= 36'sb100000101111000010111101111010000001;
            sine_reg0   <= 36'sb111001001011100011001101000100001100;
        end
        2189: begin
            cosine_reg0 <= 36'sb100000101111101101111101110110000010;
            sine_reg0   <= 36'sb111001001000011110110010110011111011;
        end
        2190: begin
            cosine_reg0 <= 36'sb100000110000011001010001000011111010;
            sine_reg0   <= 36'sb111001000101011010011100110010110001;
        end
        2191: begin
            cosine_reg0 <= 36'sb100000110001000100110111100011010000;
            sine_reg0   <= 36'sb111001000010010110001011000010101000;
        end
        2192: begin
            cosine_reg0 <= 36'sb100000110001110000110001010011101000;
            sine_reg0   <= 36'sb111000111111010001111101100101011000;
        end
        2193: begin
            cosine_reg0 <= 36'sb100000110010011100111110010100100111;
            sine_reg0   <= 36'sb111000111100001101110100011100111011;
        end
        2194: begin
            cosine_reg0 <= 36'sb100000110011001001011110100101110010;
            sine_reg0   <= 36'sb111000111001001001101111101011001010;
        end
        2195: begin
            cosine_reg0 <= 36'sb100000110011110110010010000110101110;
            sine_reg0   <= 36'sb111000110110000101101111010001111110;
        end
        2196: begin
            cosine_reg0 <= 36'sb100000110100100011011000110110111111;
            sine_reg0   <= 36'sb111000110011000001110011010011001111;
        end
        2197: begin
            cosine_reg0 <= 36'sb100000110101010000110010110110001001;
            sine_reg0   <= 36'sb111000101111111101111011110000110111;
        end
        2198: begin
            cosine_reg0 <= 36'sb100000110101111110100000000011101111;
            sine_reg0   <= 36'sb111000101100111010001000101100101101;
        end
        2199: begin
            cosine_reg0 <= 36'sb100000110110101100100000011111010111;
            sine_reg0   <= 36'sb111000101001110110011010001000101100;
        end
        2200: begin
            cosine_reg0 <= 36'sb100000110111011010110100001000100011;
            sine_reg0   <= 36'sb111000100110110010110000000110101100;
        end
        2201: begin
            cosine_reg0 <= 36'sb100000111000001001011010111110111000;
            sine_reg0   <= 36'sb111000100011101111001010101000100101;
        end
        2202: begin
            cosine_reg0 <= 36'sb100000111000111000010101000001110111;
            sine_reg0   <= 36'sb111000100000101011101001110000010000;
        end
        2203: begin
            cosine_reg0 <= 36'sb100000111001100111100010010001000100;
            sine_reg0   <= 36'sb111000011101101000001101011111100110;
        end
        2204: begin
            cosine_reg0 <= 36'sb100000111010010111000010101100000011;
            sine_reg0   <= 36'sb111000011010100100110101111000011111;
        end
        2205: begin
            cosine_reg0 <= 36'sb100000111011000110110110010010010110;
            sine_reg0   <= 36'sb111000010111100001100010111100110100;
        end
        2206: begin
            cosine_reg0 <= 36'sb100000111011110110111101000011011111;
            sine_reg0   <= 36'sb111000010100011110010100101110011101;
        end
        2207: begin
            cosine_reg0 <= 36'sb100000111100100111010110111111000000;
            sine_reg0   <= 36'sb111000010001011011001011001111010011;
        end
        2208: begin
            cosine_reg0 <= 36'sb100000111101011000000100000100011100;
            sine_reg0   <= 36'sb111000001110011000000110100001001110;
        end
        2209: begin
            cosine_reg0 <= 36'sb100000111110001001000100010011010101;
            sine_reg0   <= 36'sb111000001011010101000110100110000110;
        end
        2210: begin
            cosine_reg0 <= 36'sb100000111110111010010111101011001101;
            sine_reg0   <= 36'sb111000001000010010001011011111110100;
        end
        2211: begin
            cosine_reg0 <= 36'sb100000111111101011111110001011100101;
            sine_reg0   <= 36'sb111000000101001111010101010000010000;
        end
        2212: begin
            cosine_reg0 <= 36'sb100001000000011101110111110011111110;
            sine_reg0   <= 36'sb111000000010001100100011111001010010;
        end
        2213: begin
            cosine_reg0 <= 36'sb100001000001010000000100100011111010;
            sine_reg0   <= 36'sb110111111111001001110111011100110010;
        end
        2214: begin
            cosine_reg0 <= 36'sb100001000010000010100100011010111010;
            sine_reg0   <= 36'sb110111111100000111001111111100101001;
        end
        2215: begin
            cosine_reg0 <= 36'sb100001000010110101010111011000011110;
            sine_reg0   <= 36'sb110111111001000100101101011010101110;
        end
        2216: begin
            cosine_reg0 <= 36'sb100001000011101000011101011100001000;
            sine_reg0   <= 36'sb110111110110000010001111111000111001;
        end
        2217: begin
            cosine_reg0 <= 36'sb100001000100011011110110100101010111;
            sine_reg0   <= 36'sb110111110010111111110111011001000011;
        end
        2218: begin
            cosine_reg0 <= 36'sb100001000101001111100010110011101101;
            sine_reg0   <= 36'sb110111101111111101100011111101000011;
        end
        2219: begin
            cosine_reg0 <= 36'sb100001000110000011100010000110101001;
            sine_reg0   <= 36'sb110111101100111011010101100110110001;
        end
        2220: begin
            cosine_reg0 <= 36'sb100001000110110111110100011101101010;
            sine_reg0   <= 36'sb110111101001111001001100011000000101;
        end
        2221: begin
            cosine_reg0 <= 36'sb100001000111101100011001111000010010;
            sine_reg0   <= 36'sb110111100110110111001000010010110110;
        end
        2222: begin
            cosine_reg0 <= 36'sb100001001000100001010010010101111111;
            sine_reg0   <= 36'sb110111100011110101001001011000111101;
        end
        2223: begin
            cosine_reg0 <= 36'sb100001001001010110011101110110010001;
            sine_reg0   <= 36'sb110111100000110011001111101100010001;
        end
        2224: begin
            cosine_reg0 <= 36'sb100001001010001011111100011000100111;
            sine_reg0   <= 36'sb110111011101110001011011001110101010;
        end
        2225: begin
            cosine_reg0 <= 36'sb100001001011000001101101111100100000;
            sine_reg0   <= 36'sb110111011010101111101100000001111111;
        end
        2226: begin
            cosine_reg0 <= 36'sb100001001011110111110010100001011011;
            sine_reg0   <= 36'sb110111010111101110000010001000000111;
        end
        2227: begin
            cosine_reg0 <= 36'sb100001001100101110001010000110110110;
            sine_reg0   <= 36'sb110111010100101100011101100010111011;
        end
        2228: begin
            cosine_reg0 <= 36'sb100001001101100100110100101100010000;
            sine_reg0   <= 36'sb110111010001101010111110010100010001;
        end
        2229: begin
            cosine_reg0 <= 36'sb100001001110011011110010010001000111;
            sine_reg0   <= 36'sb110111001110101001100100011110000010;
        end
        2230: begin
            cosine_reg0 <= 36'sb100001001111010011000010110100111010;
            sine_reg0   <= 36'sb110111001011101000010000000010000011;
        end
        2231: begin
            cosine_reg0 <= 36'sb100001010000001010100110010111000110;
            sine_reg0   <= 36'sb110111001000100111000001000010001101;
        end
        2232: begin
            cosine_reg0 <= 36'sb100001010001000010011100110111001001;
            sine_reg0   <= 36'sb110111000101100101110111100000010111;
        end
        2233: begin
            cosine_reg0 <= 36'sb100001010001111010100110010100100001;
            sine_reg0   <= 36'sb110111000010100100110011011110010111;
        end
        2234: begin
            cosine_reg0 <= 36'sb100001010010110011000010101110101010;
            sine_reg0   <= 36'sb110110111111100011110100111110000101;
        end
        2235: begin
            cosine_reg0 <= 36'sb100001010011101011110010000101000011;
            sine_reg0   <= 36'sb110110111100100010111100000001011001;
        end
        2236: begin
            cosine_reg0 <= 36'sb100001010100100100110100010111000111;
            sine_reg0   <= 36'sb110110111001100010001000101010001000;
        end
        2237: begin
            cosine_reg0 <= 36'sb100001010101011110001001100100010100;
            sine_reg0   <= 36'sb110110110110100001011010111010001010;
        end
        2238: begin
            cosine_reg0 <= 36'sb100001010110010111110001101100000111;
            sine_reg0   <= 36'sb110110110011100000110010110011010110;
        end
        2239: begin
            cosine_reg0 <= 36'sb100001010111010001101100101101111100;
            sine_reg0   <= 36'sb110110110000100000010000010111100010;
        end
        2240: begin
            cosine_reg0 <= 36'sb100001011000001011111010101001001111;
            sine_reg0   <= 36'sb110110101101011111110011101000100110;
        end
        2241: begin
            cosine_reg0 <= 36'sb100001011001000110011011011101011101;
            sine_reg0   <= 36'sb110110101010011111011100101000010111;
        end
        2242: begin
            cosine_reg0 <= 36'sb100001011010000001001111001010000001;
            sine_reg0   <= 36'sb110110100111011111001011011000101110;
        end
        2243: begin
            cosine_reg0 <= 36'sb100001011010111100010101101110010110;
            sine_reg0   <= 36'sb110110100100011110111111111011011111;
        end
        2244: begin
            cosine_reg0 <= 36'sb100001011011110111101111001001111001;
            sine_reg0   <= 36'sb110110100001011110111010010010100011;
        end
        2245: begin
            cosine_reg0 <= 36'sb100001011100110011011011011100000110;
            sine_reg0   <= 36'sb110110011110011110111010011111101111;
        end
        2246: begin
            cosine_reg0 <= 36'sb100001011101101111011010100100010110;
            sine_reg0   <= 36'sb110110011011011111000000100100111001;
        end
        2247: begin
            cosine_reg0 <= 36'sb100001011110101011101100100010000101;
            sine_reg0   <= 36'sb110110011000011111001100100011111001;
        end
        2248: begin
            cosine_reg0 <= 36'sb100001011111101000010001010100101110;
            sine_reg0   <= 36'sb110110010101011111011110011110100100;
        end
        2249: begin
            cosine_reg0 <= 36'sb100001100000100101001000111011101011;
            sine_reg0   <= 36'sb110110010010011111110110010110110001;
        end
        2250: begin
            cosine_reg0 <= 36'sb100001100001100010010011010110011000;
            sine_reg0   <= 36'sb110110001111100000010100001110010110;
        end
        2251: begin
            cosine_reg0 <= 36'sb100001100010011111110000100100001101;
            sine_reg0   <= 36'sb110110001100100000111000000111001001;
        end
        2252: begin
            cosine_reg0 <= 36'sb100001100011011101100000100100100110;
            sine_reg0   <= 36'sb110110001001100001100010000011000000;
        end
        2253: begin
            cosine_reg0 <= 36'sb100001100100011011100011010110111100;
            sine_reg0   <= 36'sb110110000110100010010010000011110001;
        end
        2254: begin
            cosine_reg0 <= 36'sb100001100101011001111000111010101010;
            sine_reg0   <= 36'sb110110000011100011001000001011010010;
        end
        2255: begin
            cosine_reg0 <= 36'sb100001100110011000100001001111000111;
            sine_reg0   <= 36'sb110110000000100100000100011011011010;
        end
        2256: begin
            cosine_reg0 <= 36'sb100001100111010111011100010011101111;
            sine_reg0   <= 36'sb110101111101100101000110110101111101;
        end
        2257: begin
            cosine_reg0 <= 36'sb100001101000010110101010000111111001;
            sine_reg0   <= 36'sb110101111010100110001111011100110011;
        end
        2258: begin
            cosine_reg0 <= 36'sb100001101001010110001010101011000000;
            sine_reg0   <= 36'sb110101110111100111011110010001101111;
        end
        2259: begin
            cosine_reg0 <= 36'sb100001101010010101111101111100011011;
            sine_reg0   <= 36'sb110101110100101000110011010110101001;
        end
        2260: begin
            cosine_reg0 <= 36'sb100001101011010110000011111011100100;
            sine_reg0   <= 36'sb110101110001101010001110101101010101;
        end
        2261: begin
            cosine_reg0 <= 36'sb100001101100010110011100100111110011;
            sine_reg0   <= 36'sb110101101110101011110000010111101010;
        end
        2262: begin
            cosine_reg0 <= 36'sb100001101101010111001000000000100000;
            sine_reg0   <= 36'sb110101101011101101011000010111011101;
        end
        2263: begin
            cosine_reg0 <= 36'sb100001101110011000000110000101000100;
            sine_reg0   <= 36'sb110101101000101111000110101110100011;
        end
        2264: begin
            cosine_reg0 <= 36'sb100001101111011001010110110100110110;
            sine_reg0   <= 36'sb110101100101110000111011011110110001;
        end
        2265: begin
            cosine_reg0 <= 36'sb100001110000011010111010001111001110;
            sine_reg0   <= 36'sb110101100010110010110110101001111110;
        end
        2266: begin
            cosine_reg0 <= 36'sb100001110001011100110000010011100011;
            sine_reg0   <= 36'sb110101011111110100111000010001111101;
        end
        2267: begin
            cosine_reg0 <= 36'sb100001110010011110111001000001001110;
            sine_reg0   <= 36'sb110101011100110111000000011000100101;
        end
        2268: begin
            cosine_reg0 <= 36'sb100001110011100001010100010111100101;
            sine_reg0   <= 36'sb110101011001111001001110111111101010;
        end
        2269: begin
            cosine_reg0 <= 36'sb100001110100100100000010010101111111;
            sine_reg0   <= 36'sb110101010110111011100100001001000010;
        end
        2270: begin
            cosine_reg0 <= 36'sb100001110101100111000010111011110011;
            sine_reg0   <= 36'sb110101010011111101111111110110100010;
        end
        2271: begin
            cosine_reg0 <= 36'sb100001110110101010010110001000010111;
            sine_reg0   <= 36'sb110101010001000000100010001001111110;
        end
        2272: begin
            cosine_reg0 <= 36'sb100001110111101101111011111011000011;
            sine_reg0   <= 36'sb110101001110000011001011000101001011;
        end
        2273: begin
            cosine_reg0 <= 36'sb100001111000110001110100010011001101;
            sine_reg0   <= 36'sb110101001011000101111010101001111110;
        end
        2274: begin
            cosine_reg0 <= 36'sb100001111001110101111111010000001010;
            sine_reg0   <= 36'sb110101001000001000110000111010001101;
        end
        2275: begin
            cosine_reg0 <= 36'sb100001111010111010011100110001010001;
            sine_reg0   <= 36'sb110101000101001011101101110111101010;
        end
        2276: begin
            cosine_reg0 <= 36'sb100001111011111111001100110101110111;
            sine_reg0   <= 36'sb110101000010001110110001100100001101;
        end
        2277: begin
            cosine_reg0 <= 36'sb100001111101000100001111011101010010;
            sine_reg0   <= 36'sb110100111111010001111100000001100111;
        end
        2278: begin
            cosine_reg0 <= 36'sb100001111110001001100100100110110111;
            sine_reg0   <= 36'sb110100111100010101001101010001101111;
        end
        2279: begin
            cosine_reg0 <= 36'sb100001111111001111001100010001111100;
            sine_reg0   <= 36'sb110100111001011000100101010110011001;
        end
        2280: begin
            cosine_reg0 <= 36'sb100010000000010101000110011101110110;
            sine_reg0   <= 36'sb110100110110011100000100010001011000;
        end
        2281: begin
            cosine_reg0 <= 36'sb100010000001011011010011001001111001;
            sine_reg0   <= 36'sb110100110011011111101010000100100010;
        end
        2282: begin
            cosine_reg0 <= 36'sb100010000010100001110010010101011010;
            sine_reg0   <= 36'sb110100110000100011010110110001101011;
        end
        2283: begin
            cosine_reg0 <= 36'sb100010000011101000100011111111101110;
            sine_reg0   <= 36'sb110100101101100111001010011010100110;
        end
        2284: begin
            cosine_reg0 <= 36'sb100010000100101111101000001000001001;
            sine_reg0   <= 36'sb110100101010101011000101000001000111;
        end
        2285: begin
            cosine_reg0 <= 36'sb100010000101110110111110101110000000;
            sine_reg0   <= 36'sb110100100111101111000110100111000100;
        end
        2286: begin
            cosine_reg0 <= 36'sb100010000110111110100111110000100110;
            sine_reg0   <= 36'sb110100100100110011001111001110001111;
        end
        2287: begin
            cosine_reg0 <= 36'sb100010001000000110100011001111001110;
            sine_reg0   <= 36'sb110100100001110111011110111000011101;
        end
        2288: begin
            cosine_reg0 <= 36'sb100010001001001110110001001001001110;
            sine_reg0   <= 36'sb110100011110111011110101100111100001;
        end
        2289: begin
            cosine_reg0 <= 36'sb100010001010010111010001011101110111;
            sine_reg0   <= 36'sb110100011100000000010011011101001111;
        end
        2290: begin
            cosine_reg0 <= 36'sb100010001011100000000100001100011110;
            sine_reg0   <= 36'sb110100011001000100111000011011011100;
        end
        2291: begin
            cosine_reg0 <= 36'sb100010001100101001001001010100010110;
            sine_reg0   <= 36'sb110100010110001001100100100011111001;
        end
        2292: begin
            cosine_reg0 <= 36'sb100010001101110010100000110100110001;
            sine_reg0   <= 36'sb110100010011001110010111111000011100;
        end
        2293: begin
            cosine_reg0 <= 36'sb100010001110111100001010101101000010;
            sine_reg0   <= 36'sb110100010000010011010010011010110111;
        end
        2294: begin
            cosine_reg0 <= 36'sb100010010000000110000110111100011100;
            sine_reg0   <= 36'sb110100001101011000010100001100111110;
        end
        2295: begin
            cosine_reg0 <= 36'sb100010010001010000010101100010010000;
            sine_reg0   <= 36'sb110100001010011101011101010000100100;
        end
        2296: begin
            cosine_reg0 <= 36'sb100010010010011010110110011101110011;
            sine_reg0   <= 36'sb110100000111100010101101100111011101;
        end
        2297: begin
            cosine_reg0 <= 36'sb100010010011100101101001101110010100;
            sine_reg0   <= 36'sb110100000100101000000101010011011011;
        end
        2298: begin
            cosine_reg0 <= 36'sb100010010100110000101111010011000111;
            sine_reg0   <= 36'sb110100000001101101100100010110010010;
        end
        2299: begin
            cosine_reg0 <= 36'sb100010010101111100000111001011011101;
            sine_reg0   <= 36'sb110011111110110011001010110001110101;
        end
        2300: begin
            cosine_reg0 <= 36'sb100010010111000111110001010110100111;
            sine_reg0   <= 36'sb110011111011111000111000100111110111;
        end
        2301: begin
            cosine_reg0 <= 36'sb100010011000010011101101110011110111;
            sine_reg0   <= 36'sb110011111000111110101101111010001010;
        end
        2302: begin
            cosine_reg0 <= 36'sb100010011001011111111100100010011110;
            sine_reg0   <= 36'sb110011110110000100101010101010100010;
        end
        2303: begin
            cosine_reg0 <= 36'sb100010011010101100011101100001101101;
            sine_reg0   <= 36'sb110011110011001010101110111010110001;
        end
        2304: begin
            cosine_reg0 <= 36'sb100010011011111001010000110000110100;
            sine_reg0   <= 36'sb110011110000010000111010101100101011;
        end
        2305: begin
            cosine_reg0 <= 36'sb100010011101000110010110001111000101;
            sine_reg0   <= 36'sb110011101101010111001110000010000001;
        end
        2306: begin
            cosine_reg0 <= 36'sb100010011110010011101101111011110000;
            sine_reg0   <= 36'sb110011101010011101101000111100100110;
        end
        2307: begin
            cosine_reg0 <= 36'sb100010011111100001010111110110000100;
            sine_reg0   <= 36'sb110011100111100100001011011110001100;
        end
        2308: begin
            cosine_reg0 <= 36'sb100010100000101111010011111101010011;
            sine_reg0   <= 36'sb110011100100101010110101101000100111;
        end
        2309: begin
            cosine_reg0 <= 36'sb100010100001111101100010010000101011;
            sine_reg0   <= 36'sb110011100001110001100111011101101001;
        end
        2310: begin
            cosine_reg0 <= 36'sb100010100011001100000010101111011110;
            sine_reg0   <= 36'sb110011011110111000100000111111000010;
        end
        2311: begin
            cosine_reg0 <= 36'sb100010100100011010110101011000111010;
            sine_reg0   <= 36'sb110011011011111111100010001110100111;
        end
        2312: begin
            cosine_reg0 <= 36'sb100010100101101001111010001100001110;
            sine_reg0   <= 36'sb110011011001000110101011001110001001;
        end
        2313: begin
            cosine_reg0 <= 36'sb100010100110111001010001001000101011;
            sine_reg0   <= 36'sb110011010110001101111011111111011001;
        end
        2314: begin
            cosine_reg0 <= 36'sb100010101000001000111010001101011111;
            sine_reg0   <= 36'sb110011010011010101010100100100001011;
        end
        2315: begin
            cosine_reg0 <= 36'sb100010101001011000110101011001111000;
            sine_reg0   <= 36'sb110011010000011100110100111110001111;
        end
        2316: begin
            cosine_reg0 <= 36'sb100010101010101001000010101101000111;
            sine_reg0   <= 36'sb110011001101100100011101001111011000;
        end
        2317: begin
            cosine_reg0 <= 36'sb100010101011111001100010000110011000;
            sine_reg0   <= 36'sb110011001010101100001101011001010111;
        end
        2318: begin
            cosine_reg0 <= 36'sb100010101101001010010011100100111011;
            sine_reg0   <= 36'sb110011000111110100000101011101111111;
        end
        2319: begin
            cosine_reg0 <= 36'sb100010101110011011010111000111111101;
            sine_reg0   <= 36'sb110011000100111100000101011110111111;
        end
        2320: begin
            cosine_reg0 <= 36'sb100010101111101100101100101110101101;
            sine_reg0   <= 36'sb110011000010000100001101011110001011;
        end
        2321: begin
            cosine_reg0 <= 36'sb100010110000111110010100011000011001;
            sine_reg0   <= 36'sb110010111111001100011101011101010100;
        end
        2322: begin
            cosine_reg0 <= 36'sb100010110010010000001110000100001110;
            sine_reg0   <= 36'sb110010111100010100110101011110001010;
        end
        2323: begin
            cosine_reg0 <= 36'sb100010110011100010011001110001011001;
            sine_reg0   <= 36'sb110010111001011101010101100010011111;
        end
        2324: begin
            cosine_reg0 <= 36'sb100010110100110100110111011111001001;
            sine_reg0   <= 36'sb110010110110100101111101101100000101;
        end
        2325: begin
            cosine_reg0 <= 36'sb100010110110000111100111001100101001;
            sine_reg0   <= 36'sb110010110011101110101101111100101100;
        end
        2326: begin
            cosine_reg0 <= 36'sb100010110111011010101000111001000111;
            sine_reg0   <= 36'sb110010110000110111100110010110000101;
        end
        2327: begin
            cosine_reg0 <= 36'sb100010111000101101111100100011110001;
            sine_reg0   <= 36'sb110010101110000000100110111010000010;
        end
        2328: begin
            cosine_reg0 <= 36'sb100010111010000001100010001011110001;
            sine_reg0   <= 36'sb110010101011001001101111101010010011;
        end
        2329: begin
            cosine_reg0 <= 36'sb100010111011010101011001110000010110;
            sine_reg0   <= 36'sb110010101000010011000000101000101001;
        end
        2330: begin
            cosine_reg0 <= 36'sb100010111100101001100011010000101010;
            sine_reg0   <= 36'sb110010100101011100011001110110110101;
        end
        2331: begin
            cosine_reg0 <= 36'sb100010111101111101111110101011111011;
            sine_reg0   <= 36'sb110010100010100101111011010110100111;
        end
        2332: begin
            cosine_reg0 <= 36'sb100010111111010010101100000001010100;
            sine_reg0   <= 36'sb110010011111101111100101001001110001;
        end
        2333: begin
            cosine_reg0 <= 36'sb100011000000100111101011010000000001;
            sine_reg0   <= 36'sb110010011100111001010111010010000001;
        end
        2334: begin
            cosine_reg0 <= 36'sb100011000001111100111100010111001101;
            sine_reg0   <= 36'sb110010011010000011010001110001001010;
        end
        2335: begin
            cosine_reg0 <= 36'sb100011000011010010011111010110000100;
            sine_reg0   <= 36'sb110010010111001101010100101000111011;
        end
        2336: begin
            cosine_reg0 <= 36'sb100011000100101000010100001011110010;
            sine_reg0   <= 36'sb110010010100010111011111111011000100;
        end
        2337: begin
            cosine_reg0 <= 36'sb100011000101111110011010110111100000;
            sine_reg0   <= 36'sb110010010001100001110011101001010110;
        end
        2338: begin
            cosine_reg0 <= 36'sb100011000111010100110011011000011010;
            sine_reg0   <= 36'sb110010001110101100001111110101100001;
        end
        2339: begin
            cosine_reg0 <= 36'sb100011001000101011011101101101101100;
            sine_reg0   <= 36'sb110010001011110110110100100001010100;
        end
        2340: begin
            cosine_reg0 <= 36'sb100011001010000010011001110110011110;
            sine_reg0   <= 36'sb110010001001000001100001101110100000;
        end
        2341: begin
            cosine_reg0 <= 36'sb100011001011011001100111110001111100;
            sine_reg0   <= 36'sb110010000110001100010111011110110100;
        end
        2342: begin
            cosine_reg0 <= 36'sb100011001100110001000111011111010000;
            sine_reg0   <= 36'sb110010000011010111010101110100000000;
        end
        2343: begin
            cosine_reg0 <= 36'sb100011001110001000111000111101100100;
            sine_reg0   <= 36'sb110010000000100010011100101111110101;
        end
        2344: begin
            cosine_reg0 <= 36'sb100011001111100000111100001100000010;
            sine_reg0   <= 36'sb110001111101101101101100010100000000;
        end
        2345: begin
            cosine_reg0 <= 36'sb100011010000111001010001001001110011;
            sine_reg0   <= 36'sb110001111010111001000100100010010011;
        end
        2346: begin
            cosine_reg0 <= 36'sb100011010010010001110111110110000001;
            sine_reg0   <= 36'sb110001111000000100100101011100011100;
        end
        2347: begin
            cosine_reg0 <= 36'sb100011010011101010110000001111110101;
            sine_reg0   <= 36'sb110001110101010000001111000100001010;
        end
        2348: begin
            cosine_reg0 <= 36'sb100011010101000011111010010110011001;
            sine_reg0   <= 36'sb110001110010011100000001011011001110;
        end
        2349: begin
            cosine_reg0 <= 36'sb100011010110011101010110001000110101;
            sine_reg0   <= 36'sb110001101111100111111100100011010101;
        end
        2350: begin
            cosine_reg0 <= 36'sb100011010111110111000011100110010010;
            sine_reg0   <= 36'sb110001101100110100000000011110010000;
        end
        2351: begin
            cosine_reg0 <= 36'sb100011011001010001000010101101111010;
            sine_reg0   <= 36'sb110001101010000000001101001101101100;
        end
        2352: begin
            cosine_reg0 <= 36'sb100011011010101011010011011110110100;
            sine_reg0   <= 36'sb110001100111001100100010110011011010;
        end
        2353: begin
            cosine_reg0 <= 36'sb100011011100000101110101111000001001;
            sine_reg0   <= 36'sb110001100100011001000001010001001000;
        end
        2354: begin
            cosine_reg0 <= 36'sb100011011101100000101001111001000000;
            sine_reg0   <= 36'sb110001100001100101101000101000100100;
        end
        2355: begin
            cosine_reg0 <= 36'sb100011011110111011101111100000100011;
            sine_reg0   <= 36'sb110001011110110010011000111011011110;
        end
        2356: begin
            cosine_reg0 <= 36'sb100011100000010111000110101101111000;
            sine_reg0   <= 36'sb110001011011111111010010001011100011;
        end
        2357: begin
            cosine_reg0 <= 36'sb100011100001110010101111100000001000;
            sine_reg0   <= 36'sb110001011001001100010100011010100011;
        end
        2358: begin
            cosine_reg0 <= 36'sb100011100011001110101001110110011001;
            sine_reg0   <= 36'sb110001010110011001011111101010001011;
        end
        2359: begin
            cosine_reg0 <= 36'sb100011100100101010110101101111110100;
            sine_reg0   <= 36'sb110001010011100110110011111100001011;
        end
        2360: begin
            cosine_reg0 <= 36'sb100011100110000111010011001011011111;
            sine_reg0   <= 36'sb110001010000110100010001010010010000;
        end
        2361: begin
            cosine_reg0 <= 36'sb100011100111100100000010001000100001;
            sine_reg0   <= 36'sb110001001110000001110111101110001000;
        end
        2362: begin
            cosine_reg0 <= 36'sb100011101001000001000010100110000001;
            sine_reg0   <= 36'sb110001001011001111100111010001100001;
        end
        2363: begin
            cosine_reg0 <= 36'sb100011101010011110010100100011000110;
            sine_reg0   <= 36'sb110001001000011101011111111110001010;
        end
        2364: begin
            cosine_reg0 <= 36'sb100011101011111011110111111110110110;
            sine_reg0   <= 36'sb110001000101101011100001110101110000;
        end
        2365: begin
            cosine_reg0 <= 36'sb100011101101011001101100111000010111;
            sine_reg0   <= 36'sb110001000010111001101100111010000001;
        end
        2366: begin
            cosine_reg0 <= 36'sb100011101110110111110011001110110000;
            sine_reg0   <= 36'sb110001000000001000000001001100101011;
        end
        2367: begin
            cosine_reg0 <= 36'sb100011110000010110001011000001000111;
            sine_reg0   <= 36'sb110000111101010110011110101111011100;
        end
        2368: begin
            cosine_reg0 <= 36'sb100011110001110100110100001110100001;
            sine_reg0   <= 36'sb110000111010100101000101100100000000;
        end
        2369: begin
            cosine_reg0 <= 36'sb100011110011010011101110110110000011;
            sine_reg0   <= 36'sb110000110111110011110101101100000101;
        end
        2370: begin
            cosine_reg0 <= 36'sb100011110100110010111010110110110100;
            sine_reg0   <= 36'sb110000110101000010101111001001011001;
        end
        2371: begin
            cosine_reg0 <= 36'sb100011110110010010011000001111111001;
            sine_reg0   <= 36'sb110000110010010001110001111101101001;
        end
        2372: begin
            cosine_reg0 <= 36'sb100011110111110010000111000000010111;
            sine_reg0   <= 36'sb110000101111100000111110001010100001;
        end
        2373: begin
            cosine_reg0 <= 36'sb100011111001010010000111000111010010;
            sine_reg0   <= 36'sb110000101100110000010011110001110000;
        end
        2374: begin
            cosine_reg0 <= 36'sb100011111010110010011000100011101111;
            sine_reg0   <= 36'sb110000101001111111110010110101000010;
        end
        2375: begin
            cosine_reg0 <= 36'sb100011111100010010111011010100110100;
            sine_reg0   <= 36'sb110000100111001111011011010110000100;
        end
        2376: begin
            cosine_reg0 <= 36'sb100011111101110011101111011001100100;
            sine_reg0   <= 36'sb110000100100011111001101010110100011;
        end
        2377: begin
            cosine_reg0 <= 36'sb100011111111010100110100110001000100;
            sine_reg0   <= 36'sb110000100001101111001000111000001011;
        end
        2378: begin
            cosine_reg0 <= 36'sb100100000000110110001011011010011000;
            sine_reg0   <= 36'sb110000011110111111001101111100101000;
        end
        2379: begin
            cosine_reg0 <= 36'sb100100000010010111110011010100100100;
            sine_reg0   <= 36'sb110000011100001111011100100101101001;
        end
        2380: begin
            cosine_reg0 <= 36'sb100100000011111001101100011110101100;
            sine_reg0   <= 36'sb110000011001011111110100110100111001;
        end
        2381: begin
            cosine_reg0 <= 36'sb100100000101011011110110110111110011;
            sine_reg0   <= 36'sb110000010110110000010110101100000011;
        end
        2382: begin
            cosine_reg0 <= 36'sb100100000110111110010010011110111101;
            sine_reg0   <= 36'sb110000010100000001000010001100110110;
        end
        2383: begin
            cosine_reg0 <= 36'sb100100001000100000111111010011001100;
            sine_reg0   <= 36'sb110000010001010001110111011000111100;
        end
        2384: begin
            cosine_reg0 <= 36'sb100100001010000011111101010011100101;
            sine_reg0   <= 36'sb110000001110100010110110010010000001;
        end
        2385: begin
            cosine_reg0 <= 36'sb100100001011100111001100011111001010;
            sine_reg0   <= 36'sb110000001011110011111110111001110011;
        end
        2386: begin
            cosine_reg0 <= 36'sb100100001101001010101100110100111110;
            sine_reg0   <= 36'sb110000001001000101010001010001111100;
        end
        2387: begin
            cosine_reg0 <= 36'sb100100001110101110011110010100000011;
            sine_reg0   <= 36'sb110000000110010110101101011100001000;
        end
        2388: begin
            cosine_reg0 <= 36'sb100100010000010010100000111011011100;
            sine_reg0   <= 36'sb110000000011101000010011011010000100;
        end
        2389: begin
            cosine_reg0 <= 36'sb100100010001110110110100101010001011;
            sine_reg0   <= 36'sb110000000000111010000011001101011010;
        end
        2390: begin
            cosine_reg0 <= 36'sb100100010011011011011001011111010011;
            sine_reg0   <= 36'sb101111111110001011111100110111110110;
        end
        2391: begin
            cosine_reg0 <= 36'sb100100010101000000001111011001110101;
            sine_reg0   <= 36'sb101111111011011110000000011011000011;
        end
        2392: begin
            cosine_reg0 <= 36'sb100100010110100101010110011000110011;
            sine_reg0   <= 36'sb101111111000110000001101111000101101;
        end
        2393: begin
            cosine_reg0 <= 36'sb100100011000001010101110011011001111;
            sine_reg0   <= 36'sb101111110110000010100101010010100000;
        end
        2394: begin
            cosine_reg0 <= 36'sb100100011001110000010111100000001011;
            sine_reg0   <= 36'sb101111110011010101000110101010000101;
        end
        2395: begin
            cosine_reg0 <= 36'sb100100011011010110010001100110100110;
            sine_reg0   <= 36'sb101111110000100111110010000001001001;
        end
        2396: begin
            cosine_reg0 <= 36'sb100100011100111100011100101101100100;
            sine_reg0   <= 36'sb101111101101111010100111011001010101;
        end
        2397: begin
            cosine_reg0 <= 36'sb100100011110100010111000110100000100;
            sine_reg0   <= 36'sb101111101011001101100110110100010101;
        end
        2398: begin
            cosine_reg0 <= 36'sb100100100000001001100101111001000111;
            sine_reg0   <= 36'sb101111101000100000110000010011110100;
        end
        2399: begin
            cosine_reg0 <= 36'sb100100100001110000100011111011101110;
            sine_reg0   <= 36'sb101111100101110100000011111001011100;
        end
        2400: begin
            cosine_reg0 <= 36'sb100100100011010111110010111010111011;
            sine_reg0   <= 36'sb101111100011000111100001100110111000;
        end
        2401: begin
            cosine_reg0 <= 36'sb100100100100111111010010110101101011;
            sine_reg0   <= 36'sb101111100000011011001001011101110010;
        end
        2402: begin
            cosine_reg0 <= 36'sb100100100110100111000011101011000001;
            sine_reg0   <= 36'sb101111011101101110111011011111110100;
        end
        2403: begin
            cosine_reg0 <= 36'sb100100101000001111000101011001111100;
            sine_reg0   <= 36'sb101111011011000010110111101110101001;
        end
        2404: begin
            cosine_reg0 <= 36'sb100100101001110111011000000001011100;
            sine_reg0   <= 36'sb101111011000010110111110001011111011;
        end
        2405: begin
            cosine_reg0 <= 36'sb100100101011011111111011100000100001;
            sine_reg0   <= 36'sb101111010101101011001110111001010011;
        end
        2406: begin
            cosine_reg0 <= 36'sb100100101101001000101111110110001001;
            sine_reg0   <= 36'sb101111010010111111101001111000011101;
        end
        2407: begin
            cosine_reg0 <= 36'sb100100101110110001110101000001010101;
            sine_reg0   <= 36'sb101111010000010100001111001011000001;
        end
        2408: begin
            cosine_reg0 <= 36'sb100100110000011011001011000001000100;
            sine_reg0   <= 36'sb101111001101101000111110110010101001;
        end
        2409: begin
            cosine_reg0 <= 36'sb100100110010000100110001110100010100;
            sine_reg0   <= 36'sb101111001010111101111000110001000000;
        end
        2410: begin
            cosine_reg0 <= 36'sb100100110011101110101001011010000100;
            sine_reg0   <= 36'sb101111001000010010111101000111101110;
        end
        2411: begin
            cosine_reg0 <= 36'sb100100110101011000110001110001010100;
            sine_reg0   <= 36'sb101111000101101000001011111000011101;
        end
        2412: begin
            cosine_reg0 <= 36'sb100100110111000011001010111001000001;
            sine_reg0   <= 36'sb101111000010111101100101000100110110;
        end
        2413: begin
            cosine_reg0 <= 36'sb100100111000101101110100110000001010;
            sine_reg0   <= 36'sb101111000000010011001000101110100011;
        end
        2414: begin
            cosine_reg0 <= 36'sb100100111010011000101111010101101110;
            sine_reg0   <= 36'sb101110111101101000110110110111001100;
        end
        2415: begin
            cosine_reg0 <= 36'sb100100111100000011111010101000101010;
            sine_reg0   <= 36'sb101110111010111110101111100000011100;
        end
        2416: begin
            cosine_reg0 <= 36'sb100100111101101111010110100111111100;
            sine_reg0   <= 36'sb101110111000010100110010101011111010;
        end
        2417: begin
            cosine_reg0 <= 36'sb100100111111011011000011010010100010;
            sine_reg0   <= 36'sb101110110101101011000000011011001111;
        end
        2418: begin
            cosine_reg0 <= 36'sb100101000001000111000000100111011001;
            sine_reg0   <= 36'sb101110110011000001011000110000000101;
        end
        2419: begin
            cosine_reg0 <= 36'sb100101000010110011001110100101011111;
            sine_reg0   <= 36'sb101110110000010111111011101100000100;
        end
        2420: begin
            cosine_reg0 <= 36'sb100101000100011111101101001011110010;
            sine_reg0   <= 36'sb101110101101101110101001010000110100;
        end
        2421: begin
            cosine_reg0 <= 36'sb100101000110001100011100011001001110;
            sine_reg0   <= 36'sb101110101011000101100001011111111110;
        end
        2422: begin
            cosine_reg0 <= 36'sb100101000111111001011100001100101111;
            sine_reg0   <= 36'sb101110101000011100100100011011001010;
        end
        2423: begin
            cosine_reg0 <= 36'sb100101001001100110101100100101010100;
            sine_reg0   <= 36'sb101110100101110011110010000100000000;
        end
        2424: begin
            cosine_reg0 <= 36'sb100101001011010100001101100001111000;
            sine_reg0   <= 36'sb101110100011001011001010011100001001;
        end
        2425: begin
            cosine_reg0 <= 36'sb100101001101000001111111000001011001;
            sine_reg0   <= 36'sb101110100000100010101101100101001100;
        end
        2426: begin
            cosine_reg0 <= 36'sb100101001110110000000001000010110001;
            sine_reg0   <= 36'sb101110011101111010011011100000110010;
        end
        2427: begin
            cosine_reg0 <= 36'sb100101010000011110010011100100111110;
            sine_reg0   <= 36'sb101110011011010010010100010000100010;
        end
        2428: begin
            cosine_reg0 <= 36'sb100101010010001100110110100110111011;
            sine_reg0   <= 36'sb101110011000101010010111110110000100;
        end
        2429: begin
            cosine_reg0 <= 36'sb100101010011111011101010000111100100;
            sine_reg0   <= 36'sb101110010110000010100110010010111111;
        end
        2430: begin
            cosine_reg0 <= 36'sb100101010101101010101110000101110110;
            sine_reg0   <= 36'sb101110010011011010111111101000111100;
        end
        2431: begin
            cosine_reg0 <= 36'sb100101010111011010000010100000101010;
            sine_reg0   <= 36'sb101110010000110011100011111001100000;
        end
        2432: begin
            cosine_reg0 <= 36'sb100101011001001001100111010110111101;
            sine_reg0   <= 36'sb101110001110001100010011000110010101;
        end
        2433: begin
            cosine_reg0 <= 36'sb100101011010111001011100100111101010;
            sine_reg0   <= 36'sb101110001011100101001101010001000000;
        end
        2434: begin
            cosine_reg0 <= 36'sb100101011100101001100010010001101100;
            sine_reg0   <= 36'sb101110001000111110010010011011001001;
        end
        2435: begin
            cosine_reg0 <= 36'sb100101011110011001111000010011111101;
            sine_reg0   <= 36'sb101110000110010111100010100110011000;
        end
        2436: begin
            cosine_reg0 <= 36'sb100101100000001010011110101101011001;
            sine_reg0   <= 36'sb101110000011110000111101110100010001;
        end
        2437: begin
            cosine_reg0 <= 36'sb100101100001111011010101011100111010;
            sine_reg0   <= 36'sb101110000001001010100100000110011110;
        end
        2438: begin
            cosine_reg0 <= 36'sb100101100011101100011100100001011001;
            sine_reg0   <= 36'sb101101111110100100010101011110100011;
        end
        2439: begin
            cosine_reg0 <= 36'sb100101100101011101110011111001110011;
            sine_reg0   <= 36'sb101101111011111110010001111110001000;
        end
        2440: begin
            cosine_reg0 <= 36'sb100101100111001111011011100101000000;
            sine_reg0   <= 36'sb101101111001011000011001100110110100;
        end
        2441: begin
            cosine_reg0 <= 36'sb100101101001000001010011100001111011;
            sine_reg0   <= 36'sb101101110110110010101100011010001011;
        end
        2442: begin
            cosine_reg0 <= 36'sb100101101010110011011011101111011101;
            sine_reg0   <= 36'sb101101110100001101001010011001110110;
        end
        2443: begin
            cosine_reg0 <= 36'sb100101101100100101110100001100011111;
            sine_reg0   <= 36'sb101101110001100111110011100111011001;
        end
        2444: begin
            cosine_reg0 <= 36'sb100101101110011000011100110111111100;
            sine_reg0   <= 36'sb101101101111000010101000000100011010;
        end
        2445: begin
            cosine_reg0 <= 36'sb100101110000001011010101110000101101;
            sine_reg0   <= 36'sb101101101100011101100111110010100001;
        end
        2446: begin
            cosine_reg0 <= 36'sb100101110001111110011110110101101011;
            sine_reg0   <= 36'sb101101101001111000110010110011010010;
        end
        2447: begin
            cosine_reg0 <= 36'sb100101110011110001111000000101101110;
            sine_reg0   <= 36'sb101101100111010100001001001000010011;
        end
        2448: begin
            cosine_reg0 <= 36'sb100101110101100101100001011111101111;
            sine_reg0   <= 36'sb101101100100101111101010110011001001;
        end
        2449: begin
            cosine_reg0 <= 36'sb100101110111011001011011000010101000;
            sine_reg0   <= 36'sb101101100010001011010111110101011011;
        end
        2450: begin
            cosine_reg0 <= 36'sb100101111001001101100100101101010001;
            sine_reg0   <= 36'sb101101011111100111010000010000101101;
        end
        2451: begin
            cosine_reg0 <= 36'sb100101111011000001111110011110100001;
            sine_reg0   <= 36'sb101101011101000011010100000110100101;
        end
        2452: begin
            cosine_reg0 <= 36'sb100101111100110110101000010101010010;
            sine_reg0   <= 36'sb101101011010011111100011011000101000;
        end
        2453: begin
            cosine_reg0 <= 36'sb100101111110101011100010010000011011;
            sine_reg0   <= 36'sb101101010111111011111110001000011011;
        end
        2454: begin
            cosine_reg0 <= 36'sb100110000000100000101100001110110100;
            sine_reg0   <= 36'sb101101010101011000100100010111100010;
        end
        2455: begin
            cosine_reg0 <= 36'sb100110000010010110000110001111010110;
            sine_reg0   <= 36'sb101101010010110101010110000111100011;
        end
        2456: begin
            cosine_reg0 <= 36'sb100110000100001011110000010000110110;
            sine_reg0   <= 36'sb101101010000010010010011011010000010;
        end
        2457: begin
            cosine_reg0 <= 36'sb100110000110000001101010010010001110;
            sine_reg0   <= 36'sb101101001101101111011100010000100100;
        end
        2458: begin
            cosine_reg0 <= 36'sb100110000111110111110100010010010100;
            sine_reg0   <= 36'sb101101001011001100110000101100101101;
        end
        2459: begin
            cosine_reg0 <= 36'sb100110001001101110001110001111111111;
            sine_reg0   <= 36'sb101101001000101010010000110000000010;
        end
        2460: begin
            cosine_reg0 <= 36'sb100110001011100100111000001010000110;
            sine_reg0   <= 36'sb101101000110000111111100011100000110;
        end
        2461: begin
            cosine_reg0 <= 36'sb100110001101011011110001111111100001;
            sine_reg0   <= 36'sb101101000011100101110011110010011111;
        end
        2462: begin
            cosine_reg0 <= 36'sb100110001111010010111011101111000101;
            sine_reg0   <= 36'sb101101000001000011110110110100110000;
        end
        2463: begin
            cosine_reg0 <= 36'sb100110010001001010010101010111101001;
            sine_reg0   <= 36'sb101100111110100010000101100100011100;
        end
        2464: begin
            cosine_reg0 <= 36'sb100110010011000001111110111000000100;
            sine_reg0   <= 36'sb101100111100000000100000000011001000;
        end
        2465: begin
            cosine_reg0 <= 36'sb100110010100111001111000001111001100;
            sine_reg0   <= 36'sb101100111001011111000110010010011000;
        end
        2466: begin
            cosine_reg0 <= 36'sb100110010110110010000001011011110110;
            sine_reg0   <= 36'sb101100110110111101111000010011101110;
        end
        2467: begin
            cosine_reg0 <= 36'sb100110011000101010011010011100111001;
            sine_reg0   <= 36'sb101100110100011100110110001000101111;
        end
        2468: begin
            cosine_reg0 <= 36'sb100110011010100011000011010001001011;
            sine_reg0   <= 36'sb101100110001111011111111110010111101;
        end
        2469: begin
            cosine_reg0 <= 36'sb100110011100011011111011110111100000;
            sine_reg0   <= 36'sb101100101111011011010101010011111101;
        end
        2470: begin
            cosine_reg0 <= 36'sb100110011110010101000100001110101111;
            sine_reg0   <= 36'sb101100101100111010110110101101010000;
        end
        2471: begin
            cosine_reg0 <= 36'sb100110100000001110011100010101101101;
            sine_reg0   <= 36'sb101100101010011010100100000000011011;
        end
        2472: begin
            cosine_reg0 <= 36'sb100110100010001000000100001011001111;
            sine_reg0   <= 36'sb101100100111111010011101001110111111;
        end
        2473: begin
            cosine_reg0 <= 36'sb100110100100000001111011101110001001;
            sine_reg0   <= 36'sb101100100101011010100010011010100000;
        end
        2474: begin
            cosine_reg0 <= 36'sb100110100101111100000010111101010001;
            sine_reg0   <= 36'sb101100100010111010110011100100100000;
        end
        2475: begin
            cosine_reg0 <= 36'sb100110100111110110011001110111011100;
            sine_reg0   <= 36'sb101100100000011011010000101110100010;
        end
        2476: begin
            cosine_reg0 <= 36'sb100110101001110001000000011011011101;
            sine_reg0   <= 36'sb101100011101111011111001111010001001;
        end
        2477: begin
            cosine_reg0 <= 36'sb100110101011101011110110101000001010;
            sine_reg0   <= 36'sb101100011011011100101111001000110101;
        end
        2478: begin
            cosine_reg0 <= 36'sb100110101101100110111100011100010110;
            sine_reg0   <= 36'sb101100011000111101110000011100001011;
        end
        2479: begin
            cosine_reg0 <= 36'sb100110101111100010010001110110110101;
            sine_reg0   <= 36'sb101100010110011110111101110101101011;
        end
        2480: begin
            cosine_reg0 <= 36'sb100110110001011101110110110110011100;
            sine_reg0   <= 36'sb101100010100000000010111010110111001;
        end
        2481: begin
            cosine_reg0 <= 36'sb100110110011011001101011011001111110;
            sine_reg0   <= 36'sb101100010001100001111101000001010100;
        end
        2482: begin
            cosine_reg0 <= 36'sb100110110101010101101111100000001111;
            sine_reg0   <= 36'sb101100001111000011101110110110100000;
        end
        2483: begin
            cosine_reg0 <= 36'sb100110110111010010000011001000000011;
            sine_reg0   <= 36'sb101100001100100101101100110111111110;
        end
        2484: begin
            cosine_reg0 <= 36'sb100110111001001110100110010000001100;
            sine_reg0   <= 36'sb101100001010000111110111000111001111;
        end
        2485: begin
            cosine_reg0 <= 36'sb100110111011001011011000110111011101;
            sine_reg0   <= 36'sb101100000111101010001101100101110101;
        end
        2486: begin
            cosine_reg0 <= 36'sb100110111101001000011010111100101011;
            sine_reg0   <= 36'sb101100000101001100110000010101010001;
        end
        2487: begin
            cosine_reg0 <= 36'sb100110111111000101101100011110100111;
            sine_reg0   <= 36'sb101100000010101111011111010111000100;
        end
        2488: begin
            cosine_reg0 <= 36'sb100111000001000011001101011100000101;
            sine_reg0   <= 36'sb101100000000010010011010101100101111;
        end
        2489: begin
            cosine_reg0 <= 36'sb100111000011000000111101110011110111;
            sine_reg0   <= 36'sb101011111101110101100010010111110011;
        end
        2490: begin
            cosine_reg0 <= 36'sb100111000100111110111101100100101111;
            sine_reg0   <= 36'sb101011111011011000110110011001110001;
        end
        2491: begin
            cosine_reg0 <= 36'sb100111000110111101001100101101011111;
            sine_reg0   <= 36'sb101011111000111100010110110100001010;
        end
        2492: begin
            cosine_reg0 <= 36'sb100111001000111011101011001100111011;
            sine_reg0   <= 36'sb101011110110100000000011101000011101;
        end
        2493: begin
            cosine_reg0 <= 36'sb100111001010111010011001000001110100;
            sine_reg0   <= 36'sb101011110100000011111100111000001100;
        end
        2494: begin
            cosine_reg0 <= 36'sb100111001100111001010110001010111011;
            sine_reg0   <= 36'sb101011110001101000000010100100110110;
        end
        2495: begin
            cosine_reg0 <= 36'sb100111001110111000100010100111000010;
            sine_reg0   <= 36'sb101011101111001100010100101111111100;
        end
        2496: begin
            cosine_reg0 <= 36'sb100111010000110111111110010100111100;
            sine_reg0   <= 36'sb101011101100110000110011011010111110;
        end
        2497: begin
            cosine_reg0 <= 36'sb100111010010110111101001010011011000;
            sine_reg0   <= 36'sb101011101010010101011110100111011100;
        end
        2498: begin
            cosine_reg0 <= 36'sb100111010100110111100011100001001001;
            sine_reg0   <= 36'sb101011100111111010010110010110110110;
        end
        2499: begin
            cosine_reg0 <= 36'sb100111010110110111101100111101000000;
            sine_reg0   <= 36'sb101011100101011111011010101010101011;
        end
        2500: begin
            cosine_reg0 <= 36'sb100111011000111000000101100101101101;
            sine_reg0   <= 36'sb101011100011000100101011100100011011;
        end
        2501: begin
            cosine_reg0 <= 36'sb100111011010111000101101011010000010;
            sine_reg0   <= 36'sb101011100000101010001001000101100101;
        end
        2502: begin
            cosine_reg0 <= 36'sb100111011100111001100100011000101111;
            sine_reg0   <= 36'sb101011011110001111110011001111101000;
        end
        2503: begin
            cosine_reg0 <= 36'sb100111011110111010101010100000100100;
            sine_reg0   <= 36'sb101011011011110101101010000100000101;
        end
        2504: begin
            cosine_reg0 <= 36'sb100111100000111011111111110000010010;
            sine_reg0   <= 36'sb101011011001011011101101100100011010;
        end
        2505: begin
            cosine_reg0 <= 36'sb100111100010111101100100000110101010;
            sine_reg0   <= 36'sb101011010111000001111101110010000101;
        end
        2506: begin
            cosine_reg0 <= 36'sb100111100100111111010111100010011010;
            sine_reg0   <= 36'sb101011010100101000011010101110100111;
        end
        2507: begin
            cosine_reg0 <= 36'sb100111100111000001011010000010010100;
            sine_reg0   <= 36'sb101011010010001111000100011011011101;
        end
        2508: begin
            cosine_reg0 <= 36'sb100111101001000011101011100101000110;
            sine_reg0   <= 36'sb101011001111110101111010111010000110;
        end
        2509: begin
            cosine_reg0 <= 36'sb100111101011000110001100001001100010;
            sine_reg0   <= 36'sb101011001101011100111110001100000000;
        end
        2510: begin
            cosine_reg0 <= 36'sb100111101101001000111011101110010101;
            sine_reg0   <= 36'sb101011001011000100001110010010101010;
        end
        2511: begin
            cosine_reg0 <= 36'sb100111101111001011111010010010010000;
            sine_reg0   <= 36'sb101011001000101011101011001111100011;
        end
        2512: begin
            cosine_reg0 <= 36'sb100111110001001111000111110100000001;
            sine_reg0   <= 36'sb101011000110010011010101000100001000;
        end
        2513: begin
            cosine_reg0 <= 36'sb100111110011010010100100010010011000;
            sine_reg0   <= 36'sb101011000011111011001011110001110111;
        end
        2514: begin
            cosine_reg0 <= 36'sb100111110101010110001111101100000011;
            sine_reg0   <= 36'sb101011000001100011001111011010001101;
        end
        2515: begin
            cosine_reg0 <= 36'sb100111110111011010001001111111110010;
            sine_reg0   <= 36'sb101010111111001011011111111110101010;
        end
        2516: begin
            cosine_reg0 <= 36'sb100111111001011110010011001100010011;
            sine_reg0   <= 36'sb101010111100110011111101100000101010;
        end
        2517: begin
            cosine_reg0 <= 36'sb100111111011100010101011010000010101;
            sine_reg0   <= 36'sb101010111010011100101000000001101011;
        end
        2518: begin
            cosine_reg0 <= 36'sb100111111101100111010010001010100101;
            sine_reg0   <= 36'sb101010111000000101011111100011001010;
        end
        2519: begin
            cosine_reg0 <= 36'sb100111111111101100000111111001110011;
            sine_reg0   <= 36'sb101010110101101110100100000110100101;
        end
        2520: begin
            cosine_reg0 <= 36'sb101000000001110001001100011100101011;
            sine_reg0   <= 36'sb101010110011010111110101101101011000;
        end
        2521: begin
            cosine_reg0 <= 36'sb101000000011110110011111110001111100;
            sine_reg0   <= 36'sb101010110001000001010100011001000000;
        end
        2522: begin
            cosine_reg0 <= 36'sb101000000101111100000001111000010101;
            sine_reg0   <= 36'sb101010101110101011000000001010111011;
        end
        2523: begin
            cosine_reg0 <= 36'sb101000001000000001110010101110100001;
            sine_reg0   <= 36'sb101010101100010100111001000100100101;
        end
        2524: begin
            cosine_reg0 <= 36'sb101000001010000111110010010011010000;
            sine_reg0   <= 36'sb101010101001111110111111000111011011;
        end
        2525: begin
            cosine_reg0 <= 36'sb101000001100001110000000100101001110;
            sine_reg0   <= 36'sb101010100111101001010010010100111001;
        end
        2526: begin
            cosine_reg0 <= 36'sb101000001110010100011101100011001000;
            sine_reg0   <= 36'sb101010100101010011110010101110011011;
        end
        2527: begin
            cosine_reg0 <= 36'sb101000010000011011001001001011101100;
            sine_reg0   <= 36'sb101010100010111110100000010101011110;
        end
        2528: begin
            cosine_reg0 <= 36'sb101000010010100010000011011101100110;
            sine_reg0   <= 36'sb101010100000101001011011001011011101;
        end
        2529: begin
            cosine_reg0 <= 36'sb101000010100101001001100010111100100;
            sine_reg0   <= 36'sb101010011110010100100011010001110110;
        end
        2530: begin
            cosine_reg0 <= 36'sb101000010110110000100011111000010001;
            sine_reg0   <= 36'sb101010011011111111111000101010000011;
        end
        2531: begin
            cosine_reg0 <= 36'sb101000011000111000001001111110011011;
            sine_reg0   <= 36'sb101010011001101011011011010101100000;
        end
        2532: begin
            cosine_reg0 <= 36'sb101000011010111111111110101000101101;
            sine_reg0   <= 36'sb101010010111010111001011010101101001;
        end
        2533: begin
            cosine_reg0 <= 36'sb101000011101001000000001110101110100;
            sine_reg0   <= 36'sb101010010101000011001000101011111010;
        end
        2534: begin
            cosine_reg0 <= 36'sb101000011111010000010011100100011101;
            sine_reg0   <= 36'sb101010010010101111010011011001101101;
        end
        2535: begin
            cosine_reg0 <= 36'sb101000100001011000110011110011010010;
            sine_reg0   <= 36'sb101010010000011011101011100000011110;
        end
        2536: begin
            cosine_reg0 <= 36'sb101000100011100001100010100001000000;
            sine_reg0   <= 36'sb101010001110001000010001000001100111;
        end
        2537: begin
            cosine_reg0 <= 36'sb101000100101101010011111101100010010;
            sine_reg0   <= 36'sb101010001011110101000011111110100101;
        end
        2538: begin
            cosine_reg0 <= 36'sb101000100111110011101011010011110101;
            sine_reg0   <= 36'sb101010001001100010000100011000110001;
        end
        2539: begin
            cosine_reg0 <= 36'sb101000101001111101000101010110010010;
            sine_reg0   <= 36'sb101010000111001111010010010001100111;
        end
        2540: begin
            cosine_reg0 <= 36'sb101000101100000110101101110010010111;
            sine_reg0   <= 36'sb101010000100111100101101101010100000;
        end
        2541: begin
            cosine_reg0 <= 36'sb101000101110010000100100100110101100;
            sine_reg0   <= 36'sb101010000010101010010110100100110111;
        end
        2542: begin
            cosine_reg0 <= 36'sb101000110000011010101001110001111111;
            sine_reg0   <= 36'sb101010000000011000001101000010000111;
        end
        2543: begin
            cosine_reg0 <= 36'sb101000110010100100111101010010111001;
            sine_reg0   <= 36'sb101001111110000110010001000011101010;
        end
        2544: begin
            cosine_reg0 <= 36'sb101000110100101111011111001000000101;
            sine_reg0   <= 36'sb101001111011110100100010101010111001;
        end
        2545: begin
            cosine_reg0 <= 36'sb101000110110111010001111010000001101;
            sine_reg0   <= 36'sb101001111001100011000001111001001111;
        end
        2546: begin
            cosine_reg0 <= 36'sb101000111001000101001101101001111101;
            sine_reg0   <= 36'sb101001110111010001101110110000000110;
        end
        2547: begin
            cosine_reg0 <= 36'sb101000111011010000011010010011111110;
            sine_reg0   <= 36'sb101001110101000000101001010000110110;
        end
        2548: begin
            cosine_reg0 <= 36'sb101000111101011011110101001100111011;
            sine_reg0   <= 36'sb101001110010101111110001011100111010;
        end
        2549: begin
            cosine_reg0 <= 36'sb101000111111100111011110010011011101;
            sine_reg0   <= 36'sb101001110000011111000111010101101010;
        end
        2550: begin
            cosine_reg0 <= 36'sb101001000001110011010101100110001110;
            sine_reg0   <= 36'sb101001101110001110101010111100100001;
        end
        2551: begin
            cosine_reg0 <= 36'sb101001000011111111011011000011111001;
            sine_reg0   <= 36'sb101001101011111110011100010010110111;
        end
        2552: begin
            cosine_reg0 <= 36'sb101001000110001011101110101011000110;
            sine_reg0   <= 36'sb101001101001101110011011011010000101;
        end
        2553: begin
            cosine_reg0 <= 36'sb101001001000011000010000011010011111;
            sine_reg0   <= 36'sb101001100111011110101000010011100011;
        end
        2554: begin
            cosine_reg0 <= 36'sb101001001010100101000000010000101110;
            sine_reg0   <= 36'sb101001100101001111000011000000101100;
        end
        2555: begin
            cosine_reg0 <= 36'sb101001001100110001111110001100011011;
            sine_reg0   <= 36'sb101001100010111111101011100010110111;
        end
        2556: begin
            cosine_reg0 <= 36'sb101001001110111111001010001100010000;
            sine_reg0   <= 36'sb101001100000110000100001111011011100;
        end
        2557: begin
            cosine_reg0 <= 36'sb101001010001001100100100001110110110;
            sine_reg0   <= 36'sb101001011110100001100110001011110101;
        end
        2558: begin
            cosine_reg0 <= 36'sb101001010011011010001100010010110101;
            sine_reg0   <= 36'sb101001011100010010111000010101011000;
        end
        2559: begin
            cosine_reg0 <= 36'sb101001010101101000000010010110110110;
            sine_reg0   <= 36'sb101001011010000100011000011001011111;
        end
        2560: begin
            cosine_reg0 <= 36'sb101001010111110110000110011001100001;
            sine_reg0   <= 36'sb101001010111110110000110011001100001;
        end
        2561: begin
            cosine_reg0 <= 36'sb101001011010000100011000011001011111;
            sine_reg0   <= 36'sb101001010101101000000010010110110110;
        end
        2562: begin
            cosine_reg0 <= 36'sb101001011100010010111000010101011000;
            sine_reg0   <= 36'sb101001010011011010001100010010110101;
        end
        2563: begin
            cosine_reg0 <= 36'sb101001011110100001100110001011110101;
            sine_reg0   <= 36'sb101001010001001100100100001110110110;
        end
        2564: begin
            cosine_reg0 <= 36'sb101001100000110000100001111011011100;
            sine_reg0   <= 36'sb101001001110111111001010001100010000;
        end
        2565: begin
            cosine_reg0 <= 36'sb101001100010111111101011100010110111;
            sine_reg0   <= 36'sb101001001100110001111110001100011011;
        end
        2566: begin
            cosine_reg0 <= 36'sb101001100101001111000011000000101100;
            sine_reg0   <= 36'sb101001001010100101000000010000101110;
        end
        2567: begin
            cosine_reg0 <= 36'sb101001100111011110101000010011100011;
            sine_reg0   <= 36'sb101001001000011000010000011010011111;
        end
        2568: begin
            cosine_reg0 <= 36'sb101001101001101110011011011010000101;
            sine_reg0   <= 36'sb101001000110001011101110101011000110;
        end
        2569: begin
            cosine_reg0 <= 36'sb101001101011111110011100010010110111;
            sine_reg0   <= 36'sb101001000011111111011011000011111001;
        end
        2570: begin
            cosine_reg0 <= 36'sb101001101110001110101010111100100001;
            sine_reg0   <= 36'sb101001000001110011010101100110001110;
        end
        2571: begin
            cosine_reg0 <= 36'sb101001110000011111000111010101101010;
            sine_reg0   <= 36'sb101000111111100111011110010011011101;
        end
        2572: begin
            cosine_reg0 <= 36'sb101001110010101111110001011100111010;
            sine_reg0   <= 36'sb101000111101011011110101001100111011;
        end
        2573: begin
            cosine_reg0 <= 36'sb101001110101000000101001010000110110;
            sine_reg0   <= 36'sb101000111011010000011010010011111110;
        end
        2574: begin
            cosine_reg0 <= 36'sb101001110111010001101110110000000110;
            sine_reg0   <= 36'sb101000111001000101001101101001111101;
        end
        2575: begin
            cosine_reg0 <= 36'sb101001111001100011000001111001001111;
            sine_reg0   <= 36'sb101000110110111010001111010000001101;
        end
        2576: begin
            cosine_reg0 <= 36'sb101001111011110100100010101010111001;
            sine_reg0   <= 36'sb101000110100101111011111001000000101;
        end
        2577: begin
            cosine_reg0 <= 36'sb101001111110000110010001000011101010;
            sine_reg0   <= 36'sb101000110010100100111101010010111001;
        end
        2578: begin
            cosine_reg0 <= 36'sb101010000000011000001101000010000111;
            sine_reg0   <= 36'sb101000110000011010101001110001111111;
        end
        2579: begin
            cosine_reg0 <= 36'sb101010000010101010010110100100110111;
            sine_reg0   <= 36'sb101000101110010000100100100110101100;
        end
        2580: begin
            cosine_reg0 <= 36'sb101010000100111100101101101010100000;
            sine_reg0   <= 36'sb101000101100000110101101110010010111;
        end
        2581: begin
            cosine_reg0 <= 36'sb101010000111001111010010010001100111;
            sine_reg0   <= 36'sb101000101001111101000101010110010010;
        end
        2582: begin
            cosine_reg0 <= 36'sb101010001001100010000100011000110001;
            sine_reg0   <= 36'sb101000100111110011101011010011110101;
        end
        2583: begin
            cosine_reg0 <= 36'sb101010001011110101000011111110100101;
            sine_reg0   <= 36'sb101000100101101010011111101100010010;
        end
        2584: begin
            cosine_reg0 <= 36'sb101010001110001000010001000001100111;
            sine_reg0   <= 36'sb101000100011100001100010100001000000;
        end
        2585: begin
            cosine_reg0 <= 36'sb101010010000011011101011100000011110;
            sine_reg0   <= 36'sb101000100001011000110011110011010010;
        end
        2586: begin
            cosine_reg0 <= 36'sb101010010010101111010011011001101101;
            sine_reg0   <= 36'sb101000011111010000010011100100011101;
        end
        2587: begin
            cosine_reg0 <= 36'sb101010010101000011001000101011111010;
            sine_reg0   <= 36'sb101000011101001000000001110101110100;
        end
        2588: begin
            cosine_reg0 <= 36'sb101010010111010111001011010101101001;
            sine_reg0   <= 36'sb101000011010111111111110101000101101;
        end
        2589: begin
            cosine_reg0 <= 36'sb101010011001101011011011010101100000;
            sine_reg0   <= 36'sb101000011000111000001001111110011011;
        end
        2590: begin
            cosine_reg0 <= 36'sb101010011011111111111000101010000011;
            sine_reg0   <= 36'sb101000010110110000100011111000010001;
        end
        2591: begin
            cosine_reg0 <= 36'sb101010011110010100100011010001110110;
            sine_reg0   <= 36'sb101000010100101001001100010111100100;
        end
        2592: begin
            cosine_reg0 <= 36'sb101010100000101001011011001011011101;
            sine_reg0   <= 36'sb101000010010100010000011011101100110;
        end
        2593: begin
            cosine_reg0 <= 36'sb101010100010111110100000010101011110;
            sine_reg0   <= 36'sb101000010000011011001001001011101100;
        end
        2594: begin
            cosine_reg0 <= 36'sb101010100101010011110010101110011011;
            sine_reg0   <= 36'sb101000001110010100011101100011001000;
        end
        2595: begin
            cosine_reg0 <= 36'sb101010100111101001010010010100111001;
            sine_reg0   <= 36'sb101000001100001110000000100101001110;
        end
        2596: begin
            cosine_reg0 <= 36'sb101010101001111110111111000111011011;
            sine_reg0   <= 36'sb101000001010000111110010010011010000;
        end
        2597: begin
            cosine_reg0 <= 36'sb101010101100010100111001000100100101;
            sine_reg0   <= 36'sb101000001000000001110010101110100001;
        end
        2598: begin
            cosine_reg0 <= 36'sb101010101110101011000000001010111011;
            sine_reg0   <= 36'sb101000000101111100000001111000010101;
        end
        2599: begin
            cosine_reg0 <= 36'sb101010110001000001010100011001000000;
            sine_reg0   <= 36'sb101000000011110110011111110001111100;
        end
        2600: begin
            cosine_reg0 <= 36'sb101010110011010111110101101101011000;
            sine_reg0   <= 36'sb101000000001110001001100011100101011;
        end
        2601: begin
            cosine_reg0 <= 36'sb101010110101101110100100000110100101;
            sine_reg0   <= 36'sb100111111111101100000111111001110011;
        end
        2602: begin
            cosine_reg0 <= 36'sb101010111000000101011111100011001010;
            sine_reg0   <= 36'sb100111111101100111010010001010100101;
        end
        2603: begin
            cosine_reg0 <= 36'sb101010111010011100101000000001101011;
            sine_reg0   <= 36'sb100111111011100010101011010000010101;
        end
        2604: begin
            cosine_reg0 <= 36'sb101010111100110011111101100000101010;
            sine_reg0   <= 36'sb100111111001011110010011001100010011;
        end
        2605: begin
            cosine_reg0 <= 36'sb101010111111001011011111111110101010;
            sine_reg0   <= 36'sb100111110111011010001001111111110010;
        end
        2606: begin
            cosine_reg0 <= 36'sb101011000001100011001111011010001101;
            sine_reg0   <= 36'sb100111110101010110001111101100000011;
        end
        2607: begin
            cosine_reg0 <= 36'sb101011000011111011001011110001110111;
            sine_reg0   <= 36'sb100111110011010010100100010010011000;
        end
        2608: begin
            cosine_reg0 <= 36'sb101011000110010011010101000100001000;
            sine_reg0   <= 36'sb100111110001001111000111110100000001;
        end
        2609: begin
            cosine_reg0 <= 36'sb101011001000101011101011001111100011;
            sine_reg0   <= 36'sb100111101111001011111010010010010000;
        end
        2610: begin
            cosine_reg0 <= 36'sb101011001011000100001110010010101010;
            sine_reg0   <= 36'sb100111101101001000111011101110010101;
        end
        2611: begin
            cosine_reg0 <= 36'sb101011001101011100111110001100000000;
            sine_reg0   <= 36'sb100111101011000110001100001001100010;
        end
        2612: begin
            cosine_reg0 <= 36'sb101011001111110101111010111010000110;
            sine_reg0   <= 36'sb100111101001000011101011100101000110;
        end
        2613: begin
            cosine_reg0 <= 36'sb101011010010001111000100011011011101;
            sine_reg0   <= 36'sb100111100111000001011010000010010100;
        end
        2614: begin
            cosine_reg0 <= 36'sb101011010100101000011010101110100111;
            sine_reg0   <= 36'sb100111100100111111010111100010011010;
        end
        2615: begin
            cosine_reg0 <= 36'sb101011010111000001111101110010000101;
            sine_reg0   <= 36'sb100111100010111101100100000110101010;
        end
        2616: begin
            cosine_reg0 <= 36'sb101011011001011011101101100100011010;
            sine_reg0   <= 36'sb100111100000111011111111110000010010;
        end
        2617: begin
            cosine_reg0 <= 36'sb101011011011110101101010000100000101;
            sine_reg0   <= 36'sb100111011110111010101010100000100100;
        end
        2618: begin
            cosine_reg0 <= 36'sb101011011110001111110011001111101000;
            sine_reg0   <= 36'sb100111011100111001100100011000101111;
        end
        2619: begin
            cosine_reg0 <= 36'sb101011100000101010001001000101100101;
            sine_reg0   <= 36'sb100111011010111000101101011010000010;
        end
        2620: begin
            cosine_reg0 <= 36'sb101011100011000100101011100100011011;
            sine_reg0   <= 36'sb100111011000111000000101100101101101;
        end
        2621: begin
            cosine_reg0 <= 36'sb101011100101011111011010101010101011;
            sine_reg0   <= 36'sb100111010110110111101100111101000000;
        end
        2622: begin
            cosine_reg0 <= 36'sb101011100111111010010110010110110110;
            sine_reg0   <= 36'sb100111010100110111100011100001001001;
        end
        2623: begin
            cosine_reg0 <= 36'sb101011101010010101011110100111011100;
            sine_reg0   <= 36'sb100111010010110111101001010011011000;
        end
        2624: begin
            cosine_reg0 <= 36'sb101011101100110000110011011010111110;
            sine_reg0   <= 36'sb100111010000110111111110010100111100;
        end
        2625: begin
            cosine_reg0 <= 36'sb101011101111001100010100101111111100;
            sine_reg0   <= 36'sb100111001110111000100010100111000010;
        end
        2626: begin
            cosine_reg0 <= 36'sb101011110001101000000010100100110110;
            sine_reg0   <= 36'sb100111001100111001010110001010111011;
        end
        2627: begin
            cosine_reg0 <= 36'sb101011110100000011111100111000001100;
            sine_reg0   <= 36'sb100111001010111010011001000001110100;
        end
        2628: begin
            cosine_reg0 <= 36'sb101011110110100000000011101000011101;
            sine_reg0   <= 36'sb100111001000111011101011001100111011;
        end
        2629: begin
            cosine_reg0 <= 36'sb101011111000111100010110110100001010;
            sine_reg0   <= 36'sb100111000110111101001100101101011111;
        end
        2630: begin
            cosine_reg0 <= 36'sb101011111011011000110110011001110001;
            sine_reg0   <= 36'sb100111000100111110111101100100101111;
        end
        2631: begin
            cosine_reg0 <= 36'sb101011111101110101100010010111110011;
            sine_reg0   <= 36'sb100111000011000000111101110011110111;
        end
        2632: begin
            cosine_reg0 <= 36'sb101100000000010010011010101100101111;
            sine_reg0   <= 36'sb100111000001000011001101011100000101;
        end
        2633: begin
            cosine_reg0 <= 36'sb101100000010101111011111010111000100;
            sine_reg0   <= 36'sb100110111111000101101100011110100111;
        end
        2634: begin
            cosine_reg0 <= 36'sb101100000101001100110000010101010001;
            sine_reg0   <= 36'sb100110111101001000011010111100101011;
        end
        2635: begin
            cosine_reg0 <= 36'sb101100000111101010001101100101110101;
            sine_reg0   <= 36'sb100110111011001011011000110111011101;
        end
        2636: begin
            cosine_reg0 <= 36'sb101100001010000111110111000111001111;
            sine_reg0   <= 36'sb100110111001001110100110010000001100;
        end
        2637: begin
            cosine_reg0 <= 36'sb101100001100100101101100110111111110;
            sine_reg0   <= 36'sb100110110111010010000011001000000011;
        end
        2638: begin
            cosine_reg0 <= 36'sb101100001111000011101110110110100000;
            sine_reg0   <= 36'sb100110110101010101101111100000001111;
        end
        2639: begin
            cosine_reg0 <= 36'sb101100010001100001111101000001010100;
            sine_reg0   <= 36'sb100110110011011001101011011001111110;
        end
        2640: begin
            cosine_reg0 <= 36'sb101100010100000000010111010110111001;
            sine_reg0   <= 36'sb100110110001011101110110110110011100;
        end
        2641: begin
            cosine_reg0 <= 36'sb101100010110011110111101110101101011;
            sine_reg0   <= 36'sb100110101111100010010001110110110101;
        end
        2642: begin
            cosine_reg0 <= 36'sb101100011000111101110000011100001011;
            sine_reg0   <= 36'sb100110101101100110111100011100010110;
        end
        2643: begin
            cosine_reg0 <= 36'sb101100011011011100101111001000110101;
            sine_reg0   <= 36'sb100110101011101011110110101000001010;
        end
        2644: begin
            cosine_reg0 <= 36'sb101100011101111011111001111010001001;
            sine_reg0   <= 36'sb100110101001110001000000011011011101;
        end
        2645: begin
            cosine_reg0 <= 36'sb101100100000011011010000101110100010;
            sine_reg0   <= 36'sb100110100111110110011001110111011100;
        end
        2646: begin
            cosine_reg0 <= 36'sb101100100010111010110011100100100000;
            sine_reg0   <= 36'sb100110100101111100000010111101010001;
        end
        2647: begin
            cosine_reg0 <= 36'sb101100100101011010100010011010100000;
            sine_reg0   <= 36'sb100110100100000001111011101110001001;
        end
        2648: begin
            cosine_reg0 <= 36'sb101100100111111010011101001110111111;
            sine_reg0   <= 36'sb100110100010001000000100001011001111;
        end
        2649: begin
            cosine_reg0 <= 36'sb101100101010011010100100000000011011;
            sine_reg0   <= 36'sb100110100000001110011100010101101101;
        end
        2650: begin
            cosine_reg0 <= 36'sb101100101100111010110110101101010000;
            sine_reg0   <= 36'sb100110011110010101000100001110101111;
        end
        2651: begin
            cosine_reg0 <= 36'sb101100101111011011010101010011111101;
            sine_reg0   <= 36'sb100110011100011011111011110111100000;
        end
        2652: begin
            cosine_reg0 <= 36'sb101100110001111011111111110010111101;
            sine_reg0   <= 36'sb100110011010100011000011010001001011;
        end
        2653: begin
            cosine_reg0 <= 36'sb101100110100011100110110001000101111;
            sine_reg0   <= 36'sb100110011000101010011010011100111001;
        end
        2654: begin
            cosine_reg0 <= 36'sb101100110110111101111000010011101110;
            sine_reg0   <= 36'sb100110010110110010000001011011110110;
        end
        2655: begin
            cosine_reg0 <= 36'sb101100111001011111000110010010011000;
            sine_reg0   <= 36'sb100110010100111001111000001111001100;
        end
        2656: begin
            cosine_reg0 <= 36'sb101100111100000000100000000011001000;
            sine_reg0   <= 36'sb100110010011000001111110111000000100;
        end
        2657: begin
            cosine_reg0 <= 36'sb101100111110100010000101100100011100;
            sine_reg0   <= 36'sb100110010001001010010101010111101001;
        end
        2658: begin
            cosine_reg0 <= 36'sb101101000001000011110110110100110000;
            sine_reg0   <= 36'sb100110001111010010111011101111000101;
        end
        2659: begin
            cosine_reg0 <= 36'sb101101000011100101110011110010011111;
            sine_reg0   <= 36'sb100110001101011011110001111111100001;
        end
        2660: begin
            cosine_reg0 <= 36'sb101101000110000111111100011100000110;
            sine_reg0   <= 36'sb100110001011100100111000001010000110;
        end
        2661: begin
            cosine_reg0 <= 36'sb101101001000101010010000110000000010;
            sine_reg0   <= 36'sb100110001001101110001110001111111111;
        end
        2662: begin
            cosine_reg0 <= 36'sb101101001011001100110000101100101101;
            sine_reg0   <= 36'sb100110000111110111110100010010010100;
        end
        2663: begin
            cosine_reg0 <= 36'sb101101001101101111011100010000100100;
            sine_reg0   <= 36'sb100110000110000001101010010010001110;
        end
        2664: begin
            cosine_reg0 <= 36'sb101101010000010010010011011010000010;
            sine_reg0   <= 36'sb100110000100001011110000010000110110;
        end
        2665: begin
            cosine_reg0 <= 36'sb101101010010110101010110000111100011;
            sine_reg0   <= 36'sb100110000010010110000110001111010110;
        end
        2666: begin
            cosine_reg0 <= 36'sb101101010101011000100100010111100010;
            sine_reg0   <= 36'sb100110000000100000101100001110110100;
        end
        2667: begin
            cosine_reg0 <= 36'sb101101010111111011111110001000011011;
            sine_reg0   <= 36'sb100101111110101011100010010000011011;
        end
        2668: begin
            cosine_reg0 <= 36'sb101101011010011111100011011000101000;
            sine_reg0   <= 36'sb100101111100110110101000010101010010;
        end
        2669: begin
            cosine_reg0 <= 36'sb101101011101000011010100000110100101;
            sine_reg0   <= 36'sb100101111011000001111110011110100001;
        end
        2670: begin
            cosine_reg0 <= 36'sb101101011111100111010000010000101101;
            sine_reg0   <= 36'sb100101111001001101100100101101010001;
        end
        2671: begin
            cosine_reg0 <= 36'sb101101100010001011010111110101011011;
            sine_reg0   <= 36'sb100101110111011001011011000010101000;
        end
        2672: begin
            cosine_reg0 <= 36'sb101101100100101111101010110011001001;
            sine_reg0   <= 36'sb100101110101100101100001011111101111;
        end
        2673: begin
            cosine_reg0 <= 36'sb101101100111010100001001001000010011;
            sine_reg0   <= 36'sb100101110011110001111000000101101110;
        end
        2674: begin
            cosine_reg0 <= 36'sb101101101001111000110010110011010010;
            sine_reg0   <= 36'sb100101110001111110011110110101101011;
        end
        2675: begin
            cosine_reg0 <= 36'sb101101101100011101100111110010100001;
            sine_reg0   <= 36'sb100101110000001011010101110000101101;
        end
        2676: begin
            cosine_reg0 <= 36'sb101101101111000010101000000100011010;
            sine_reg0   <= 36'sb100101101110011000011100110111111100;
        end
        2677: begin
            cosine_reg0 <= 36'sb101101110001100111110011100111011001;
            sine_reg0   <= 36'sb100101101100100101110100001100011111;
        end
        2678: begin
            cosine_reg0 <= 36'sb101101110100001101001010011001110110;
            sine_reg0   <= 36'sb100101101010110011011011101111011101;
        end
        2679: begin
            cosine_reg0 <= 36'sb101101110110110010101100011010001011;
            sine_reg0   <= 36'sb100101101001000001010011100001111011;
        end
        2680: begin
            cosine_reg0 <= 36'sb101101111001011000011001100110110100;
            sine_reg0   <= 36'sb100101100111001111011011100101000000;
        end
        2681: begin
            cosine_reg0 <= 36'sb101101111011111110010001111110001000;
            sine_reg0   <= 36'sb100101100101011101110011111001110011;
        end
        2682: begin
            cosine_reg0 <= 36'sb101101111110100100010101011110100011;
            sine_reg0   <= 36'sb100101100011101100011100100001011001;
        end
        2683: begin
            cosine_reg0 <= 36'sb101110000001001010100100000110011110;
            sine_reg0   <= 36'sb100101100001111011010101011100111010;
        end
        2684: begin
            cosine_reg0 <= 36'sb101110000011110000111101110100010001;
            sine_reg0   <= 36'sb100101100000001010011110101101011001;
        end
        2685: begin
            cosine_reg0 <= 36'sb101110000110010111100010100110011000;
            sine_reg0   <= 36'sb100101011110011001111000010011111101;
        end
        2686: begin
            cosine_reg0 <= 36'sb101110001000111110010010011011001001;
            sine_reg0   <= 36'sb100101011100101001100010010001101100;
        end
        2687: begin
            cosine_reg0 <= 36'sb101110001011100101001101010001000000;
            sine_reg0   <= 36'sb100101011010111001011100100111101010;
        end
        2688: begin
            cosine_reg0 <= 36'sb101110001110001100010011000110010101;
            sine_reg0   <= 36'sb100101011001001001100111010110111101;
        end
        2689: begin
            cosine_reg0 <= 36'sb101110010000110011100011111001100000;
            sine_reg0   <= 36'sb100101010111011010000010100000101010;
        end
        2690: begin
            cosine_reg0 <= 36'sb101110010011011010111111101000111100;
            sine_reg0   <= 36'sb100101010101101010101110000101110110;
        end
        2691: begin
            cosine_reg0 <= 36'sb101110010110000010100110010010111111;
            sine_reg0   <= 36'sb100101010011111011101010000111100100;
        end
        2692: begin
            cosine_reg0 <= 36'sb101110011000101010010111110110000100;
            sine_reg0   <= 36'sb100101010010001100110110100110111011;
        end
        2693: begin
            cosine_reg0 <= 36'sb101110011011010010010100010000100010;
            sine_reg0   <= 36'sb100101010000011110010011100100111110;
        end
        2694: begin
            cosine_reg0 <= 36'sb101110011101111010011011100000110010;
            sine_reg0   <= 36'sb100101001110110000000001000010110001;
        end
        2695: begin
            cosine_reg0 <= 36'sb101110100000100010101101100101001100;
            sine_reg0   <= 36'sb100101001101000001111111000001011001;
        end
        2696: begin
            cosine_reg0 <= 36'sb101110100011001011001010011100001001;
            sine_reg0   <= 36'sb100101001011010100001101100001111000;
        end
        2697: begin
            cosine_reg0 <= 36'sb101110100101110011110010000100000000;
            sine_reg0   <= 36'sb100101001001100110101100100101010100;
        end
        2698: begin
            cosine_reg0 <= 36'sb101110101000011100100100011011001010;
            sine_reg0   <= 36'sb100101000111111001011100001100101111;
        end
        2699: begin
            cosine_reg0 <= 36'sb101110101011000101100001011111111110;
            sine_reg0   <= 36'sb100101000110001100011100011001001110;
        end
        2700: begin
            cosine_reg0 <= 36'sb101110101101101110101001010000110100;
            sine_reg0   <= 36'sb100101000100011111101101001011110010;
        end
        2701: begin
            cosine_reg0 <= 36'sb101110110000010111111011101100000100;
            sine_reg0   <= 36'sb100101000010110011001110100101011111;
        end
        2702: begin
            cosine_reg0 <= 36'sb101110110011000001011000110000000101;
            sine_reg0   <= 36'sb100101000001000111000000100111011001;
        end
        2703: begin
            cosine_reg0 <= 36'sb101110110101101011000000011011001111;
            sine_reg0   <= 36'sb100100111111011011000011010010100010;
        end
        2704: begin
            cosine_reg0 <= 36'sb101110111000010100110010101011111010;
            sine_reg0   <= 36'sb100100111101101111010110100111111100;
        end
        2705: begin
            cosine_reg0 <= 36'sb101110111010111110101111100000011100;
            sine_reg0   <= 36'sb100100111100000011111010101000101010;
        end
        2706: begin
            cosine_reg0 <= 36'sb101110111101101000110110110111001100;
            sine_reg0   <= 36'sb100100111010011000101111010101101110;
        end
        2707: begin
            cosine_reg0 <= 36'sb101111000000010011001000101110100011;
            sine_reg0   <= 36'sb100100111000101101110100110000001010;
        end
        2708: begin
            cosine_reg0 <= 36'sb101111000010111101100101000100110110;
            sine_reg0   <= 36'sb100100110111000011001010111001000001;
        end
        2709: begin
            cosine_reg0 <= 36'sb101111000101101000001011111000011101;
            sine_reg0   <= 36'sb100100110101011000110001110001010100;
        end
        2710: begin
            cosine_reg0 <= 36'sb101111001000010010111101000111101110;
            sine_reg0   <= 36'sb100100110011101110101001011010000100;
        end
        2711: begin
            cosine_reg0 <= 36'sb101111001010111101111000110001000000;
            sine_reg0   <= 36'sb100100110010000100110001110100010100;
        end
        2712: begin
            cosine_reg0 <= 36'sb101111001101101000111110110010101001;
            sine_reg0   <= 36'sb100100110000011011001011000001000100;
        end
        2713: begin
            cosine_reg0 <= 36'sb101111010000010100001111001011000001;
            sine_reg0   <= 36'sb100100101110110001110101000001010101;
        end
        2714: begin
            cosine_reg0 <= 36'sb101111010010111111101001111000011101;
            sine_reg0   <= 36'sb100100101101001000101111110110001001;
        end
        2715: begin
            cosine_reg0 <= 36'sb101111010101101011001110111001010011;
            sine_reg0   <= 36'sb100100101011011111111011100000100001;
        end
        2716: begin
            cosine_reg0 <= 36'sb101111011000010110111110001011111011;
            sine_reg0   <= 36'sb100100101001110111011000000001011100;
        end
        2717: begin
            cosine_reg0 <= 36'sb101111011011000010110111101110101001;
            sine_reg0   <= 36'sb100100101000001111000101011001111100;
        end
        2718: begin
            cosine_reg0 <= 36'sb101111011101101110111011011111110100;
            sine_reg0   <= 36'sb100100100110100111000011101011000001;
        end
        2719: begin
            cosine_reg0 <= 36'sb101111100000011011001001011101110010;
            sine_reg0   <= 36'sb100100100100111111010010110101101011;
        end
        2720: begin
            cosine_reg0 <= 36'sb101111100011000111100001100110111000;
            sine_reg0   <= 36'sb100100100011010111110010111010111011;
        end
        2721: begin
            cosine_reg0 <= 36'sb101111100101110100000011111001011100;
            sine_reg0   <= 36'sb100100100001110000100011111011101110;
        end
        2722: begin
            cosine_reg0 <= 36'sb101111101000100000110000010011110100;
            sine_reg0   <= 36'sb100100100000001001100101111001000111;
        end
        2723: begin
            cosine_reg0 <= 36'sb101111101011001101100110110100010101;
            sine_reg0   <= 36'sb100100011110100010111000110100000100;
        end
        2724: begin
            cosine_reg0 <= 36'sb101111101101111010100111011001010101;
            sine_reg0   <= 36'sb100100011100111100011100101101100100;
        end
        2725: begin
            cosine_reg0 <= 36'sb101111110000100111110010000001001001;
            sine_reg0   <= 36'sb100100011011010110010001100110100110;
        end
        2726: begin
            cosine_reg0 <= 36'sb101111110011010101000110101010000101;
            sine_reg0   <= 36'sb100100011001110000010111100000001011;
        end
        2727: begin
            cosine_reg0 <= 36'sb101111110110000010100101010010100000;
            sine_reg0   <= 36'sb100100011000001010101110011011001111;
        end
        2728: begin
            cosine_reg0 <= 36'sb101111111000110000001101111000101101;
            sine_reg0   <= 36'sb100100010110100101010110011000110011;
        end
        2729: begin
            cosine_reg0 <= 36'sb101111111011011110000000011011000011;
            sine_reg0   <= 36'sb100100010101000000001111011001110101;
        end
        2730: begin
            cosine_reg0 <= 36'sb101111111110001011111100110111110110;
            sine_reg0   <= 36'sb100100010011011011011001011111010011;
        end
        2731: begin
            cosine_reg0 <= 36'sb110000000000111010000011001101011010;
            sine_reg0   <= 36'sb100100010001110110110100101010001011;
        end
        2732: begin
            cosine_reg0 <= 36'sb110000000011101000010011011010000100;
            sine_reg0   <= 36'sb100100010000010010100000111011011100;
        end
        2733: begin
            cosine_reg0 <= 36'sb110000000110010110101101011100001000;
            sine_reg0   <= 36'sb100100001110101110011110010100000011;
        end
        2734: begin
            cosine_reg0 <= 36'sb110000001001000101010001010001111100;
            sine_reg0   <= 36'sb100100001101001010101100110100111110;
        end
        2735: begin
            cosine_reg0 <= 36'sb110000001011110011111110111001110011;
            sine_reg0   <= 36'sb100100001011100111001100011111001010;
        end
        2736: begin
            cosine_reg0 <= 36'sb110000001110100010110110010010000001;
            sine_reg0   <= 36'sb100100001010000011111101010011100101;
        end
        2737: begin
            cosine_reg0 <= 36'sb110000010001010001110111011000111100;
            sine_reg0   <= 36'sb100100001000100000111111010011001100;
        end
        2738: begin
            cosine_reg0 <= 36'sb110000010100000001000010001100110110;
            sine_reg0   <= 36'sb100100000110111110010010011110111101;
        end
        2739: begin
            cosine_reg0 <= 36'sb110000010110110000010110101100000011;
            sine_reg0   <= 36'sb100100000101011011110110110111110011;
        end
        2740: begin
            cosine_reg0 <= 36'sb110000011001011111110100110100111001;
            sine_reg0   <= 36'sb100100000011111001101100011110101100;
        end
        2741: begin
            cosine_reg0 <= 36'sb110000011100001111011100100101101001;
            sine_reg0   <= 36'sb100100000010010111110011010100100100;
        end
        2742: begin
            cosine_reg0 <= 36'sb110000011110111111001101111100101000;
            sine_reg0   <= 36'sb100100000000110110001011011010011000;
        end
        2743: begin
            cosine_reg0 <= 36'sb110000100001101111001000111000001011;
            sine_reg0   <= 36'sb100011111111010100110100110001000100;
        end
        2744: begin
            cosine_reg0 <= 36'sb110000100100011111001101010110100011;
            sine_reg0   <= 36'sb100011111101110011101111011001100100;
        end
        2745: begin
            cosine_reg0 <= 36'sb110000100111001111011011010110000100;
            sine_reg0   <= 36'sb100011111100010010111011010100110100;
        end
        2746: begin
            cosine_reg0 <= 36'sb110000101001111111110010110101000010;
            sine_reg0   <= 36'sb100011111010110010011000100011101111;
        end
        2747: begin
            cosine_reg0 <= 36'sb110000101100110000010011110001110000;
            sine_reg0   <= 36'sb100011111001010010000111000111010010;
        end
        2748: begin
            cosine_reg0 <= 36'sb110000101111100000111110001010100001;
            sine_reg0   <= 36'sb100011110111110010000111000000010111;
        end
        2749: begin
            cosine_reg0 <= 36'sb110000110010010001110001111101101001;
            sine_reg0   <= 36'sb100011110110010010011000001111111001;
        end
        2750: begin
            cosine_reg0 <= 36'sb110000110101000010101111001001011001;
            sine_reg0   <= 36'sb100011110100110010111010110110110100;
        end
        2751: begin
            cosine_reg0 <= 36'sb110000110111110011110101101100000101;
            sine_reg0   <= 36'sb100011110011010011101110110110000011;
        end
        2752: begin
            cosine_reg0 <= 36'sb110000111010100101000101100100000000;
            sine_reg0   <= 36'sb100011110001110100110100001110100001;
        end
        2753: begin
            cosine_reg0 <= 36'sb110000111101010110011110101111011100;
            sine_reg0   <= 36'sb100011110000010110001011000001000111;
        end
        2754: begin
            cosine_reg0 <= 36'sb110001000000001000000001001100101011;
            sine_reg0   <= 36'sb100011101110110111110011001110110000;
        end
        2755: begin
            cosine_reg0 <= 36'sb110001000010111001101100111010000001;
            sine_reg0   <= 36'sb100011101101011001101100111000010111;
        end
        2756: begin
            cosine_reg0 <= 36'sb110001000101101011100001110101110000;
            sine_reg0   <= 36'sb100011101011111011110111111110110110;
        end
        2757: begin
            cosine_reg0 <= 36'sb110001001000011101011111111110001010;
            sine_reg0   <= 36'sb100011101010011110010100100011000110;
        end
        2758: begin
            cosine_reg0 <= 36'sb110001001011001111100111010001100001;
            sine_reg0   <= 36'sb100011101001000001000010100110000001;
        end
        2759: begin
            cosine_reg0 <= 36'sb110001001110000001110111101110001000;
            sine_reg0   <= 36'sb100011100111100100000010001000100001;
        end
        2760: begin
            cosine_reg0 <= 36'sb110001010000110100010001010010010000;
            sine_reg0   <= 36'sb100011100110000111010011001011011111;
        end
        2761: begin
            cosine_reg0 <= 36'sb110001010011100110110011111100001011;
            sine_reg0   <= 36'sb100011100100101010110101101111110100;
        end
        2762: begin
            cosine_reg0 <= 36'sb110001010110011001011111101010001011;
            sine_reg0   <= 36'sb100011100011001110101001110110011001;
        end
        2763: begin
            cosine_reg0 <= 36'sb110001011001001100010100011010100011;
            sine_reg0   <= 36'sb100011100001110010101111100000001000;
        end
        2764: begin
            cosine_reg0 <= 36'sb110001011011111111010010001011100011;
            sine_reg0   <= 36'sb100011100000010111000110101101111000;
        end
        2765: begin
            cosine_reg0 <= 36'sb110001011110110010011000111011011110;
            sine_reg0   <= 36'sb100011011110111011101111100000100011;
        end
        2766: begin
            cosine_reg0 <= 36'sb110001100001100101101000101000100100;
            sine_reg0   <= 36'sb100011011101100000101001111001000000;
        end
        2767: begin
            cosine_reg0 <= 36'sb110001100100011001000001010001001000;
            sine_reg0   <= 36'sb100011011100000101110101111000001001;
        end
        2768: begin
            cosine_reg0 <= 36'sb110001100111001100100010110011011010;
            sine_reg0   <= 36'sb100011011010101011010011011110110100;
        end
        2769: begin
            cosine_reg0 <= 36'sb110001101010000000001101001101101100;
            sine_reg0   <= 36'sb100011011001010001000010101101111010;
        end
        2770: begin
            cosine_reg0 <= 36'sb110001101100110100000000011110010000;
            sine_reg0   <= 36'sb100011010111110111000011100110010010;
        end
        2771: begin
            cosine_reg0 <= 36'sb110001101111100111111100100011010101;
            sine_reg0   <= 36'sb100011010110011101010110001000110101;
        end
        2772: begin
            cosine_reg0 <= 36'sb110001110010011100000001011011001110;
            sine_reg0   <= 36'sb100011010101000011111010010110011001;
        end
        2773: begin
            cosine_reg0 <= 36'sb110001110101010000001111000100001010;
            sine_reg0   <= 36'sb100011010011101010110000001111110101;
        end
        2774: begin
            cosine_reg0 <= 36'sb110001111000000100100101011100011100;
            sine_reg0   <= 36'sb100011010010010001110111110110000001;
        end
        2775: begin
            cosine_reg0 <= 36'sb110001111010111001000100100010010011;
            sine_reg0   <= 36'sb100011010000111001010001001001110011;
        end
        2776: begin
            cosine_reg0 <= 36'sb110001111101101101101100010100000000;
            sine_reg0   <= 36'sb100011001111100000111100001100000010;
        end
        2777: begin
            cosine_reg0 <= 36'sb110010000000100010011100101111110101;
            sine_reg0   <= 36'sb100011001110001000111000111101100100;
        end
        2778: begin
            cosine_reg0 <= 36'sb110010000011010111010101110100000000;
            sine_reg0   <= 36'sb100011001100110001000111011111010000;
        end
        2779: begin
            cosine_reg0 <= 36'sb110010000110001100010111011110110100;
            sine_reg0   <= 36'sb100011001011011001100111110001111100;
        end
        2780: begin
            cosine_reg0 <= 36'sb110010001001000001100001101110100000;
            sine_reg0   <= 36'sb100011001010000010011001110110011110;
        end
        2781: begin
            cosine_reg0 <= 36'sb110010001011110110110100100001010100;
            sine_reg0   <= 36'sb100011001000101011011101101101101100;
        end
        2782: begin
            cosine_reg0 <= 36'sb110010001110101100001111110101100001;
            sine_reg0   <= 36'sb100011000111010100110011011000011010;
        end
        2783: begin
            cosine_reg0 <= 36'sb110010010001100001110011101001010110;
            sine_reg0   <= 36'sb100011000101111110011010110111100000;
        end
        2784: begin
            cosine_reg0 <= 36'sb110010010100010111011111111011000100;
            sine_reg0   <= 36'sb100011000100101000010100001011110010;
        end
        2785: begin
            cosine_reg0 <= 36'sb110010010111001101010100101000111011;
            sine_reg0   <= 36'sb100011000011010010011111010110000100;
        end
        2786: begin
            cosine_reg0 <= 36'sb110010011010000011010001110001001010;
            sine_reg0   <= 36'sb100011000001111100111100010111001101;
        end
        2787: begin
            cosine_reg0 <= 36'sb110010011100111001010111010010000001;
            sine_reg0   <= 36'sb100011000000100111101011010000000001;
        end
        2788: begin
            cosine_reg0 <= 36'sb110010011111101111100101001001110001;
            sine_reg0   <= 36'sb100010111111010010101100000001010100;
        end
        2789: begin
            cosine_reg0 <= 36'sb110010100010100101111011010110100111;
            sine_reg0   <= 36'sb100010111101111101111110101011111011;
        end
        2790: begin
            cosine_reg0 <= 36'sb110010100101011100011001110110110101;
            sine_reg0   <= 36'sb100010111100101001100011010000101010;
        end
        2791: begin
            cosine_reg0 <= 36'sb110010101000010011000000101000101001;
            sine_reg0   <= 36'sb100010111011010101011001110000010110;
        end
        2792: begin
            cosine_reg0 <= 36'sb110010101011001001101111101010010011;
            sine_reg0   <= 36'sb100010111010000001100010001011110001;
        end
        2793: begin
            cosine_reg0 <= 36'sb110010101110000000100110111010000010;
            sine_reg0   <= 36'sb100010111000101101111100100011110001;
        end
        2794: begin
            cosine_reg0 <= 36'sb110010110000110111100110010110000101;
            sine_reg0   <= 36'sb100010110111011010101000111001000111;
        end
        2795: begin
            cosine_reg0 <= 36'sb110010110011101110101101111100101100;
            sine_reg0   <= 36'sb100010110110000111100111001100101001;
        end
        2796: begin
            cosine_reg0 <= 36'sb110010110110100101111101101100000101;
            sine_reg0   <= 36'sb100010110100110100110111011111001001;
        end
        2797: begin
            cosine_reg0 <= 36'sb110010111001011101010101100010011111;
            sine_reg0   <= 36'sb100010110011100010011001110001011001;
        end
        2798: begin
            cosine_reg0 <= 36'sb110010111100010100110101011110001010;
            sine_reg0   <= 36'sb100010110010010000001110000100001110;
        end
        2799: begin
            cosine_reg0 <= 36'sb110010111111001100011101011101010100;
            sine_reg0   <= 36'sb100010110000111110010100011000011001;
        end
        2800: begin
            cosine_reg0 <= 36'sb110011000010000100001101011110001011;
            sine_reg0   <= 36'sb100010101111101100101100101110101101;
        end
        2801: begin
            cosine_reg0 <= 36'sb110011000100111100000101011110111111;
            sine_reg0   <= 36'sb100010101110011011010111000111111101;
        end
        2802: begin
            cosine_reg0 <= 36'sb110011000111110100000101011101111111;
            sine_reg0   <= 36'sb100010101101001010010011100100111011;
        end
        2803: begin
            cosine_reg0 <= 36'sb110011001010101100001101011001010111;
            sine_reg0   <= 36'sb100010101011111001100010000110011000;
        end
        2804: begin
            cosine_reg0 <= 36'sb110011001101100100011101001111011000;
            sine_reg0   <= 36'sb100010101010101001000010101101000111;
        end
        2805: begin
            cosine_reg0 <= 36'sb110011010000011100110100111110001111;
            sine_reg0   <= 36'sb100010101001011000110101011001111000;
        end
        2806: begin
            cosine_reg0 <= 36'sb110011010011010101010100100100001011;
            sine_reg0   <= 36'sb100010101000001000111010001101011111;
        end
        2807: begin
            cosine_reg0 <= 36'sb110011010110001101111011111111011001;
            sine_reg0   <= 36'sb100010100110111001010001001000101011;
        end
        2808: begin
            cosine_reg0 <= 36'sb110011011001000110101011001110001001;
            sine_reg0   <= 36'sb100010100101101001111010001100001110;
        end
        2809: begin
            cosine_reg0 <= 36'sb110011011011111111100010001110100111;
            sine_reg0   <= 36'sb100010100100011010110101011000111010;
        end
        2810: begin
            cosine_reg0 <= 36'sb110011011110111000100000111111000010;
            sine_reg0   <= 36'sb100010100011001100000010101111011110;
        end
        2811: begin
            cosine_reg0 <= 36'sb110011100001110001100111011101101001;
            sine_reg0   <= 36'sb100010100001111101100010010000101011;
        end
        2812: begin
            cosine_reg0 <= 36'sb110011100100101010110101101000100111;
            sine_reg0   <= 36'sb100010100000101111010011111101010011;
        end
        2813: begin
            cosine_reg0 <= 36'sb110011100111100100001011011110001100;
            sine_reg0   <= 36'sb100010011111100001010111110110000100;
        end
        2814: begin
            cosine_reg0 <= 36'sb110011101010011101101000111100100110;
            sine_reg0   <= 36'sb100010011110010011101101111011110000;
        end
        2815: begin
            cosine_reg0 <= 36'sb110011101101010111001110000010000001;
            sine_reg0   <= 36'sb100010011101000110010110001111000101;
        end
        2816: begin
            cosine_reg0 <= 36'sb110011110000010000111010101100101011;
            sine_reg0   <= 36'sb100010011011111001010000110000110100;
        end
        2817: begin
            cosine_reg0 <= 36'sb110011110011001010101110111010110001;
            sine_reg0   <= 36'sb100010011010101100011101100001101101;
        end
        2818: begin
            cosine_reg0 <= 36'sb110011110110000100101010101010100010;
            sine_reg0   <= 36'sb100010011001011111111100100010011110;
        end
        2819: begin
            cosine_reg0 <= 36'sb110011111000111110101101111010001010;
            sine_reg0   <= 36'sb100010011000010011101101110011110111;
        end
        2820: begin
            cosine_reg0 <= 36'sb110011111011111000111000100111110111;
            sine_reg0   <= 36'sb100010010111000111110001010110100111;
        end
        2821: begin
            cosine_reg0 <= 36'sb110011111110110011001010110001110101;
            sine_reg0   <= 36'sb100010010101111100000111001011011101;
        end
        2822: begin
            cosine_reg0 <= 36'sb110100000001101101100100010110010010;
            sine_reg0   <= 36'sb100010010100110000101111010011000111;
        end
        2823: begin
            cosine_reg0 <= 36'sb110100000100101000000101010011011011;
            sine_reg0   <= 36'sb100010010011100101101001101110010100;
        end
        2824: begin
            cosine_reg0 <= 36'sb110100000111100010101101100111011101;
            sine_reg0   <= 36'sb100010010010011010110110011101110011;
        end
        2825: begin
            cosine_reg0 <= 36'sb110100001010011101011101010000100100;
            sine_reg0   <= 36'sb100010010001010000010101100010010000;
        end
        2826: begin
            cosine_reg0 <= 36'sb110100001101011000010100001100111110;
            sine_reg0   <= 36'sb100010010000000110000110111100011100;
        end
        2827: begin
            cosine_reg0 <= 36'sb110100010000010011010010011010110111;
            sine_reg0   <= 36'sb100010001110111100001010101101000010;
        end
        2828: begin
            cosine_reg0 <= 36'sb110100010011001110010111111000011100;
            sine_reg0   <= 36'sb100010001101110010100000110100110001;
        end
        2829: begin
            cosine_reg0 <= 36'sb110100010110001001100100100011111001;
            sine_reg0   <= 36'sb100010001100101001001001010100010110;
        end
        2830: begin
            cosine_reg0 <= 36'sb110100011001000100111000011011011100;
            sine_reg0   <= 36'sb100010001011100000000100001100011110;
        end
        2831: begin
            cosine_reg0 <= 36'sb110100011100000000010011011101001111;
            sine_reg0   <= 36'sb100010001010010111010001011101110111;
        end
        2832: begin
            cosine_reg0 <= 36'sb110100011110111011110101100111100001;
            sine_reg0   <= 36'sb100010001001001110110001001001001110;
        end
        2833: begin
            cosine_reg0 <= 36'sb110100100001110111011110111000011101;
            sine_reg0   <= 36'sb100010001000000110100011001111001110;
        end
        2834: begin
            cosine_reg0 <= 36'sb110100100100110011001111001110001111;
            sine_reg0   <= 36'sb100010000110111110100111110000100110;
        end
        2835: begin
            cosine_reg0 <= 36'sb110100100111101111000110100111000100;
            sine_reg0   <= 36'sb100010000101110110111110101110000000;
        end
        2836: begin
            cosine_reg0 <= 36'sb110100101010101011000101000001000111;
            sine_reg0   <= 36'sb100010000100101111101000001000001001;
        end
        2837: begin
            cosine_reg0 <= 36'sb110100101101100111001010011010100110;
            sine_reg0   <= 36'sb100010000011101000100011111111101110;
        end
        2838: begin
            cosine_reg0 <= 36'sb110100110000100011010110110001101011;
            sine_reg0   <= 36'sb100010000010100001110010010101011010;
        end
        2839: begin
            cosine_reg0 <= 36'sb110100110011011111101010000100100010;
            sine_reg0   <= 36'sb100010000001011011010011001001111001;
        end
        2840: begin
            cosine_reg0 <= 36'sb110100110110011100000100010001011000;
            sine_reg0   <= 36'sb100010000000010101000110011101110110;
        end
        2841: begin
            cosine_reg0 <= 36'sb110100111001011000100101010110011001;
            sine_reg0   <= 36'sb100001111111001111001100010001111100;
        end
        2842: begin
            cosine_reg0 <= 36'sb110100111100010101001101010001101111;
            sine_reg0   <= 36'sb100001111110001001100100100110110111;
        end
        2843: begin
            cosine_reg0 <= 36'sb110100111111010001111100000001100111;
            sine_reg0   <= 36'sb100001111101000100001111011101010010;
        end
        2844: begin
            cosine_reg0 <= 36'sb110101000010001110110001100100001101;
            sine_reg0   <= 36'sb100001111011111111001100110101110111;
        end
        2845: begin
            cosine_reg0 <= 36'sb110101000101001011101101110111101010;
            sine_reg0   <= 36'sb100001111010111010011100110001010001;
        end
        2846: begin
            cosine_reg0 <= 36'sb110101001000001000110000111010001101;
            sine_reg0   <= 36'sb100001111001110101111111010000001010;
        end
        2847: begin
            cosine_reg0 <= 36'sb110101001011000101111010101001111110;
            sine_reg0   <= 36'sb100001111000110001110100010011001101;
        end
        2848: begin
            cosine_reg0 <= 36'sb110101001110000011001011000101001011;
            sine_reg0   <= 36'sb100001110111101101111011111011000011;
        end
        2849: begin
            cosine_reg0 <= 36'sb110101010001000000100010001001111110;
            sine_reg0   <= 36'sb100001110110101010010110001000010111;
        end
        2850: begin
            cosine_reg0 <= 36'sb110101010011111101111111110110100010;
            sine_reg0   <= 36'sb100001110101100111000010111011110011;
        end
        2851: begin
            cosine_reg0 <= 36'sb110101010110111011100100001001000010;
            sine_reg0   <= 36'sb100001110100100100000010010101111111;
        end
        2852: begin
            cosine_reg0 <= 36'sb110101011001111001001110111111101010;
            sine_reg0   <= 36'sb100001110011100001010100010111100101;
        end
        2853: begin
            cosine_reg0 <= 36'sb110101011100110111000000011000100101;
            sine_reg0   <= 36'sb100001110010011110111001000001001110;
        end
        2854: begin
            cosine_reg0 <= 36'sb110101011111110100111000010001111101;
            sine_reg0   <= 36'sb100001110001011100110000010011100011;
        end
        2855: begin
            cosine_reg0 <= 36'sb110101100010110010110110101001111110;
            sine_reg0   <= 36'sb100001110000011010111010001111001110;
        end
        2856: begin
            cosine_reg0 <= 36'sb110101100101110000111011011110110001;
            sine_reg0   <= 36'sb100001101111011001010110110100110110;
        end
        2857: begin
            cosine_reg0 <= 36'sb110101101000101111000110101110100011;
            sine_reg0   <= 36'sb100001101110011000000110000101000100;
        end
        2858: begin
            cosine_reg0 <= 36'sb110101101011101101011000010111011101;
            sine_reg0   <= 36'sb100001101101010111001000000000100000;
        end
        2859: begin
            cosine_reg0 <= 36'sb110101101110101011110000010111101010;
            sine_reg0   <= 36'sb100001101100010110011100100111110011;
        end
        2860: begin
            cosine_reg0 <= 36'sb110101110001101010001110101101010101;
            sine_reg0   <= 36'sb100001101011010110000011111011100100;
        end
        2861: begin
            cosine_reg0 <= 36'sb110101110100101000110011010110101001;
            sine_reg0   <= 36'sb100001101010010101111101111100011011;
        end
        2862: begin
            cosine_reg0 <= 36'sb110101110111100111011110010001101111;
            sine_reg0   <= 36'sb100001101001010110001010101011000000;
        end
        2863: begin
            cosine_reg0 <= 36'sb110101111010100110001111011100110011;
            sine_reg0   <= 36'sb100001101000010110101010000111111001;
        end
        2864: begin
            cosine_reg0 <= 36'sb110101111101100101000110110101111101;
            sine_reg0   <= 36'sb100001100111010111011100010011101111;
        end
        2865: begin
            cosine_reg0 <= 36'sb110110000000100100000100011011011010;
            sine_reg0   <= 36'sb100001100110011000100001001111000111;
        end
        2866: begin
            cosine_reg0 <= 36'sb110110000011100011001000001011010010;
            sine_reg0   <= 36'sb100001100101011001111000111010101010;
        end
        2867: begin
            cosine_reg0 <= 36'sb110110000110100010010010000011110001;
            sine_reg0   <= 36'sb100001100100011011100011010110111100;
        end
        2868: begin
            cosine_reg0 <= 36'sb110110001001100001100010000011000000;
            sine_reg0   <= 36'sb100001100011011101100000100100100110;
        end
        2869: begin
            cosine_reg0 <= 36'sb110110001100100000111000000111001001;
            sine_reg0   <= 36'sb100001100010011111110000100100001101;
        end
        2870: begin
            cosine_reg0 <= 36'sb110110001111100000010100001110010110;
            sine_reg0   <= 36'sb100001100001100010010011010110011000;
        end
        2871: begin
            cosine_reg0 <= 36'sb110110010010011111110110010110110001;
            sine_reg0   <= 36'sb100001100000100101001000111011101011;
        end
        2872: begin
            cosine_reg0 <= 36'sb110110010101011111011110011110100100;
            sine_reg0   <= 36'sb100001011111101000010001010100101110;
        end
        2873: begin
            cosine_reg0 <= 36'sb110110011000011111001100100011111001;
            sine_reg0   <= 36'sb100001011110101011101100100010000101;
        end
        2874: begin
            cosine_reg0 <= 36'sb110110011011011111000000100100111001;
            sine_reg0   <= 36'sb100001011101101111011010100100010110;
        end
        2875: begin
            cosine_reg0 <= 36'sb110110011110011110111010011111101111;
            sine_reg0   <= 36'sb100001011100110011011011011100000110;
        end
        2876: begin
            cosine_reg0 <= 36'sb110110100001011110111010010010100011;
            sine_reg0   <= 36'sb100001011011110111101111001001111001;
        end
        2877: begin
            cosine_reg0 <= 36'sb110110100100011110111111111011011111;
            sine_reg0   <= 36'sb100001011010111100010101101110010110;
        end
        2878: begin
            cosine_reg0 <= 36'sb110110100111011111001011011000101110;
            sine_reg0   <= 36'sb100001011010000001001111001010000001;
        end
        2879: begin
            cosine_reg0 <= 36'sb110110101010011111011100101000010111;
            sine_reg0   <= 36'sb100001011001000110011011011101011101;
        end
        2880: begin
            cosine_reg0 <= 36'sb110110101101011111110011101000100110;
            sine_reg0   <= 36'sb100001011000001011111010101001001111;
        end
        2881: begin
            cosine_reg0 <= 36'sb110110110000100000010000010111100010;
            sine_reg0   <= 36'sb100001010111010001101100101101111100;
        end
        2882: begin
            cosine_reg0 <= 36'sb110110110011100000110010110011010110;
            sine_reg0   <= 36'sb100001010110010111110001101100000111;
        end
        2883: begin
            cosine_reg0 <= 36'sb110110110110100001011010111010001010;
            sine_reg0   <= 36'sb100001010101011110001001100100010100;
        end
        2884: begin
            cosine_reg0 <= 36'sb110110111001100010001000101010001000;
            sine_reg0   <= 36'sb100001010100100100110100010111000111;
        end
        2885: begin
            cosine_reg0 <= 36'sb110110111100100010111100000001011001;
            sine_reg0   <= 36'sb100001010011101011110010000101000011;
        end
        2886: begin
            cosine_reg0 <= 36'sb110110111111100011110100111110000101;
            sine_reg0   <= 36'sb100001010010110011000010101110101010;
        end
        2887: begin
            cosine_reg0 <= 36'sb110111000010100100110011011110010111;
            sine_reg0   <= 36'sb100001010001111010100110010100100001;
        end
        2888: begin
            cosine_reg0 <= 36'sb110111000101100101110111100000010111;
            sine_reg0   <= 36'sb100001010001000010011100110111001001;
        end
        2889: begin
            cosine_reg0 <= 36'sb110111001000100111000001000010001101;
            sine_reg0   <= 36'sb100001010000001010100110010111000110;
        end
        2890: begin
            cosine_reg0 <= 36'sb110111001011101000010000000010000011;
            sine_reg0   <= 36'sb100001001111010011000010110100111010;
        end
        2891: begin
            cosine_reg0 <= 36'sb110111001110101001100100011110000010;
            sine_reg0   <= 36'sb100001001110011011110010010001000111;
        end
        2892: begin
            cosine_reg0 <= 36'sb110111010001101010111110010100010001;
            sine_reg0   <= 36'sb100001001101100100110100101100010000;
        end
        2893: begin
            cosine_reg0 <= 36'sb110111010100101100011101100010111011;
            sine_reg0   <= 36'sb100001001100101110001010000110110110;
        end
        2894: begin
            cosine_reg0 <= 36'sb110111010111101110000010001000000111;
            sine_reg0   <= 36'sb100001001011110111110010100001011011;
        end
        2895: begin
            cosine_reg0 <= 36'sb110111011010101111101100000001111111;
            sine_reg0   <= 36'sb100001001011000001101101111100100000;
        end
        2896: begin
            cosine_reg0 <= 36'sb110111011101110001011011001110101010;
            sine_reg0   <= 36'sb100001001010001011111100011000100111;
        end
        2897: begin
            cosine_reg0 <= 36'sb110111100000110011001111101100010001;
            sine_reg0   <= 36'sb100001001001010110011101110110010001;
        end
        2898: begin
            cosine_reg0 <= 36'sb110111100011110101001001011000111101;
            sine_reg0   <= 36'sb100001001000100001010010010101111111;
        end
        2899: begin
            cosine_reg0 <= 36'sb110111100110110111001000010010110110;
            sine_reg0   <= 36'sb100001000111101100011001111000010010;
        end
        2900: begin
            cosine_reg0 <= 36'sb110111101001111001001100011000000101;
            sine_reg0   <= 36'sb100001000110110111110100011101101010;
        end
        2901: begin
            cosine_reg0 <= 36'sb110111101100111011010101100110110001;
            sine_reg0   <= 36'sb100001000110000011100010000110101001;
        end
        2902: begin
            cosine_reg0 <= 36'sb110111101111111101100011111101000011;
            sine_reg0   <= 36'sb100001000101001111100010110011101101;
        end
        2903: begin
            cosine_reg0 <= 36'sb110111110010111111110111011001000011;
            sine_reg0   <= 36'sb100001000100011011110110100101010111;
        end
        2904: begin
            cosine_reg0 <= 36'sb110111110110000010001111111000111001;
            sine_reg0   <= 36'sb100001000011101000011101011100001000;
        end
        2905: begin
            cosine_reg0 <= 36'sb110111111001000100101101011010101110;
            sine_reg0   <= 36'sb100001000010110101010111011000011110;
        end
        2906: begin
            cosine_reg0 <= 36'sb110111111100000111001111111100101001;
            sine_reg0   <= 36'sb100001000010000010100100011010111010;
        end
        2907: begin
            cosine_reg0 <= 36'sb110111111111001001110111011100110010;
            sine_reg0   <= 36'sb100001000001010000000100100011111010;
        end
        2908: begin
            cosine_reg0 <= 36'sb111000000010001100100011111001010010;
            sine_reg0   <= 36'sb100001000000011101110111110011111110;
        end
        2909: begin
            cosine_reg0 <= 36'sb111000000101001111010101010000010000;
            sine_reg0   <= 36'sb100000111111101011111110001011100101;
        end
        2910: begin
            cosine_reg0 <= 36'sb111000001000010010001011011111110100;
            sine_reg0   <= 36'sb100000111110111010010111101011001101;
        end
        2911: begin
            cosine_reg0 <= 36'sb111000001011010101000110100110000110;
            sine_reg0   <= 36'sb100000111110001001000100010011010101;
        end
        2912: begin
            cosine_reg0 <= 36'sb111000001110011000000110100001001110;
            sine_reg0   <= 36'sb100000111101011000000100000100011100;
        end
        2913: begin
            cosine_reg0 <= 36'sb111000010001011011001011001111010011;
            sine_reg0   <= 36'sb100000111100100111010110111111000000;
        end
        2914: begin
            cosine_reg0 <= 36'sb111000010100011110010100101110011101;
            sine_reg0   <= 36'sb100000111011110110111101000011011111;
        end
        2915: begin
            cosine_reg0 <= 36'sb111000010111100001100010111100110100;
            sine_reg0   <= 36'sb100000111011000110110110010010010110;
        end
        2916: begin
            cosine_reg0 <= 36'sb111000011010100100110101111000011111;
            sine_reg0   <= 36'sb100000111010010111000010101100000011;
        end
        2917: begin
            cosine_reg0 <= 36'sb111000011101101000001101011111100110;
            sine_reg0   <= 36'sb100000111001100111100010010001000100;
        end
        2918: begin
            cosine_reg0 <= 36'sb111000100000101011101001110000010000;
            sine_reg0   <= 36'sb100000111000111000010101000001110111;
        end
        2919: begin
            cosine_reg0 <= 36'sb111000100011101111001010101000100101;
            sine_reg0   <= 36'sb100000111000001001011010111110111000;
        end
        2920: begin
            cosine_reg0 <= 36'sb111000100110110010110000000110101100;
            sine_reg0   <= 36'sb100000110111011010110100001000100011;
        end
        2921: begin
            cosine_reg0 <= 36'sb111000101001110110011010001000101100;
            sine_reg0   <= 36'sb100000110110101100100000011111010111;
        end
        2922: begin
            cosine_reg0 <= 36'sb111000101100111010001000101100101101;
            sine_reg0   <= 36'sb100000110101111110100000000011101111;
        end
        2923: begin
            cosine_reg0 <= 36'sb111000101111111101111011110000110111;
            sine_reg0   <= 36'sb100000110101010000110010110110001001;
        end
        2924: begin
            cosine_reg0 <= 36'sb111000110011000001110011010011001111;
            sine_reg0   <= 36'sb100000110100100011011000110110111111;
        end
        2925: begin
            cosine_reg0 <= 36'sb111000110110000101101111010001111110;
            sine_reg0   <= 36'sb100000110011110110010010000110101110;
        end
        2926: begin
            cosine_reg0 <= 36'sb111000111001001001101111101011001010;
            sine_reg0   <= 36'sb100000110011001001011110100101110010;
        end
        2927: begin
            cosine_reg0 <= 36'sb111000111100001101110100011100111011;
            sine_reg0   <= 36'sb100000110010011100111110010100100111;
        end
        2928: begin
            cosine_reg0 <= 36'sb111000111111010001111101100101011000;
            sine_reg0   <= 36'sb100000110001110000110001010011101000;
        end
        2929: begin
            cosine_reg0 <= 36'sb111001000010010110001011000010101000;
            sine_reg0   <= 36'sb100000110001000100110111100011010000;
        end
        2930: begin
            cosine_reg0 <= 36'sb111001000101011010011100110010110001;
            sine_reg0   <= 36'sb100000110000011001010001000011111010;
        end
        2931: begin
            cosine_reg0 <= 36'sb111001001000011110110010110011111011;
            sine_reg0   <= 36'sb100000101111101101111101110110000010;
        end
        2932: begin
            cosine_reg0 <= 36'sb111001001011100011001101000100001100;
            sine_reg0   <= 36'sb100000101111000010111101111010000001;
        end
        2933: begin
            cosine_reg0 <= 36'sb111001001110100111101011100001101100;
            sine_reg0   <= 36'sb100000101110011000010001010000010011;
        end
        2934: begin
            cosine_reg0 <= 36'sb111001010001101100001110001010100001;
            sine_reg0   <= 36'sb100000101101101101110111111001010010;
        end
        2935: begin
            cosine_reg0 <= 36'sb111001010100110000110100111100110010;
            sine_reg0   <= 36'sb100000101101000011110001110101011000;
        end
        2936: begin
            cosine_reg0 <= 36'sb111001010111110101011111110110100101;
            sine_reg0   <= 36'sb100000101100011001111111000100111110;
        end
        2937: begin
            cosine_reg0 <= 36'sb111001011010111010001110110110000010;
            sine_reg0   <= 36'sb100000101011110000011111101000100000;
        end
        2938: begin
            cosine_reg0 <= 36'sb111001011101111111000001111001001111;
            sine_reg0   <= 36'sb100000101011000111010011100000010101;
        end
        2939: begin
            cosine_reg0 <= 36'sb111001100001000011111000111110010010;
            sine_reg0   <= 36'sb100000101010011110011010101100111001;
        end
        2940: begin
            cosine_reg0 <= 36'sb111001100100001000110100000011010010;
            sine_reg0   <= 36'sb100000101001110101110101001110100011;
        end
        2941: begin
            cosine_reg0 <= 36'sb111001100111001101110011000110010111;
            sine_reg0   <= 36'sb100000101001001101100011000101101101;
        end
        2942: begin
            cosine_reg0 <= 36'sb111001101010010010110110000101100101;
            sine_reg0   <= 36'sb100000101000100101100100010010110000;
        end
        2943: begin
            cosine_reg0 <= 36'sb111001101101010111111100111111000100;
            sine_reg0   <= 36'sb100000100111111101111000110110000101;
        end
        2944: begin
            cosine_reg0 <= 36'sb111001110000011101000111110000111010;
            sine_reg0   <= 36'sb100000100111010110100000110000000011;
        end
        2945: begin
            cosine_reg0 <= 36'sb111001110011100010010110011001001101;
            sine_reg0   <= 36'sb100000100110101111011100000001000100;
        end
        2946: begin
            cosine_reg0 <= 36'sb111001110110100111101000110110000100;
            sine_reg0   <= 36'sb100000100110001000101010101001011111;
        end
        2947: begin
            cosine_reg0 <= 36'sb111001111001101100111111000101100101;
            sine_reg0   <= 36'sb100000100101100010001100101001101100;
        end
        2948: begin
            cosine_reg0 <= 36'sb111001111100110010011001000101110110;
            sine_reg0   <= 36'sb100000100100111100000010000010000100;
        end
        2949: begin
            cosine_reg0 <= 36'sb111001111111110111110110110100111110;
            sine_reg0   <= 36'sb100000100100010110001010110010111100;
        end
        2950: begin
            cosine_reg0 <= 36'sb111010000010111101011000010001000011;
            sine_reg0   <= 36'sb100000100011110000100110111100101110;
        end
        2951: begin
            cosine_reg0 <= 36'sb111010000110000010111101011000001011;
            sine_reg0   <= 36'sb100000100011001011010110011111110000;
        end
        2952: begin
            cosine_reg0 <= 36'sb111010001001001000100110001000011011;
            sine_reg0   <= 36'sb100000100010100110011001011100011001;
        end
        2953: begin
            cosine_reg0 <= 36'sb111010001100001110010010011111111011;
            sine_reg0   <= 36'sb100000100010000001101111110010111111;
        end
        2954: begin
            cosine_reg0 <= 36'sb111010001111010100000010011100110000;
            sine_reg0   <= 36'sb100000100001011101011001100011111010;
        end
        2955: begin
            cosine_reg0 <= 36'sb111010010010011001110101111101000000;
            sine_reg0   <= 36'sb100000100000111001010110101111100000;
        end
        2956: begin
            cosine_reg0 <= 36'sb111010010101011111101100111110110001;
            sine_reg0   <= 36'sb100000100000010101100111010110000111;
        end
        2957: begin
            cosine_reg0 <= 36'sb111010011000100101100111100000001001;
            sine_reg0   <= 36'sb100000011111110010001011011000000110;
        end
        2958: begin
            cosine_reg0 <= 36'sb111010011011101011100101011111001110;
            sine_reg0   <= 36'sb100000011111001111000010110101110001;
        end
        2959: begin
            cosine_reg0 <= 36'sb111010011110110001100110111010000111;
            sine_reg0   <= 36'sb100000011110101100001101101111011111;
        end
        2960: begin
            cosine_reg0 <= 36'sb111010100001110111101011101110110111;
            sine_reg0   <= 36'sb100000011110001001101100000101100101;
        end
        2961: begin
            cosine_reg0 <= 36'sb111010100100111101110011111011100111;
            sine_reg0   <= 36'sb100000011101100111011101111000011000;
        end
        2962: begin
            cosine_reg0 <= 36'sb111010101000000011111111011110011011;
            sine_reg0   <= 36'sb100000011101000101100011001000001110;
        end
        2963: begin
            cosine_reg0 <= 36'sb111010101011001010001110010101011001;
            sine_reg0   <= 36'sb100000011100100011111011110101011100;
        end
        2964: begin
            cosine_reg0 <= 36'sb111010101110010000100000011110100111;
            sine_reg0   <= 36'sb100000011100000010101000000000010101;
        end
        2965: begin
            cosine_reg0 <= 36'sb111010110001010110110101111000001010;
            sine_reg0   <= 36'sb100000011011100001100111101001010000;
        end
        2966: begin
            cosine_reg0 <= 36'sb111010110100011101001110100000001001;
            sine_reg0   <= 36'sb100000011011000000111010110000100000;
        end
        2967: begin
            cosine_reg0 <= 36'sb111010110111100011101010010100101000;
            sine_reg0   <= 36'sb100000011010100000100001010110011001;
        end
        2968: begin
            cosine_reg0 <= 36'sb111010111010101010001001010011101110;
            sine_reg0   <= 36'sb100000011010000000011011011011001111;
        end
        2969: begin
            cosine_reg0 <= 36'sb111010111101110000101011011011011111;
            sine_reg0   <= 36'sb100000011001100000101000111111010110;
        end
        2970: begin
            cosine_reg0 <= 36'sb111011000000110111010000101010000010;
            sine_reg0   <= 36'sb100000011001000001001010000011000010;
        end
        2971: begin
            cosine_reg0 <= 36'sb111011000011111101111000111101011101;
            sine_reg0   <= 36'sb100000011000100001111110100110100110;
        end
        2972: begin
            cosine_reg0 <= 36'sb111011000111000100100100010011110011;
            sine_reg0   <= 36'sb100000011000000011000110101010010110;
        end
        2973: begin
            cosine_reg0 <= 36'sb111011001010001011010010101011001100;
            sine_reg0   <= 36'sb100000010111100100100010001110100011;
        end
        2974: begin
            cosine_reg0 <= 36'sb111011001101010010000100000001101100;
            sine_reg0   <= 36'sb100000010111000110010001010011100010;
        end
        2975: begin
            cosine_reg0 <= 36'sb111011010000011000111000010101011000;
            sine_reg0   <= 36'sb100000010110101000010011111001100101;
        end
        2976: begin
            cosine_reg0 <= 36'sb111011010011011111101111100100010111;
            sine_reg0   <= 36'sb100000010110001010101010000000111111;
        end
        2977: begin
            cosine_reg0 <= 36'sb111011010110100110101001101100101101;
            sine_reg0   <= 36'sb100000010101101101010011101010000001;
        end
        2978: begin
            cosine_reg0 <= 36'sb111011011001101101100110101100100000;
            sine_reg0   <= 36'sb100000010101010000010000110100111110;
        end
        2979: begin
            cosine_reg0 <= 36'sb111011011100110100100110100001110101;
            sine_reg0   <= 36'sb100000010100110011100001100010000111;
        end
        2980: begin
            cosine_reg0 <= 36'sb111011011111111011101001001010110001;
            sine_reg0   <= 36'sb100000010100010111000101110001101111;
        end
        2981: begin
            cosine_reg0 <= 36'sb111011100011000010101110100101011010;
            sine_reg0   <= 36'sb100000010011111010111101100100000111;
        end
        2982: begin
            cosine_reg0 <= 36'sb111011100110001001110110101111110100;
            sine_reg0   <= 36'sb100000010011011111001000111001100001;
        end
        2983: begin
            cosine_reg0 <= 36'sb111011101001010001000001101000000101;
            sine_reg0   <= 36'sb100000010011000011100111110010001100;
        end
        2984: begin
            cosine_reg0 <= 36'sb111011101100011000001111001100010010;
            sine_reg0   <= 36'sb100000010010101000011010001110011100;
        end
        2985: begin
            cosine_reg0 <= 36'sb111011101111011111011111011010100001;
            sine_reg0   <= 36'sb100000010010001101100000001110011111;
        end
        2986: begin
            cosine_reg0 <= 36'sb111011110010100110110010010000110101;
            sine_reg0   <= 36'sb100000010001110010111001110010100111;
        end
        2987: begin
            cosine_reg0 <= 36'sb111011110101101110000111101101010101;
            sine_reg0   <= 36'sb100000010001011000100110111011000101;
        end
        2988: begin
            cosine_reg0 <= 36'sb111011111000110101011111101110000100;
            sine_reg0   <= 36'sb100000010000111110100111101000001000;
        end
        2989: begin
            cosine_reg0 <= 36'sb111011111011111100111010010001001010;
            sine_reg0   <= 36'sb100000010000100100111011111010000000;
        end
        2990: begin
            cosine_reg0 <= 36'sb111011111111000100010111010100101001;
            sine_reg0   <= 36'sb100000010000001011100011110000111110;
        end
        2991: begin
            cosine_reg0 <= 36'sb111100000010001011110110110110101000;
            sine_reg0   <= 36'sb100000001111110010011111001101010001;
        end
        2992: begin
            cosine_reg0 <= 36'sb111100000101010011011000110101001011;
            sine_reg0   <= 36'sb100000001111011001101110001111001001;
        end
        2993: begin
            cosine_reg0 <= 36'sb111100001000011010111101001110010111;
            sine_reg0   <= 36'sb100000001111000001010000110110110100;
        end
        2994: begin
            cosine_reg0 <= 36'sb111100001011100010100100000000010001;
            sine_reg0   <= 36'sb100000001110101001000111000100100010;
        end
        2995: begin
            cosine_reg0 <= 36'sb111100001110101010001101001000111110;
            sine_reg0   <= 36'sb100000001110010001010000111000100001;
        end
        2996: begin
            cosine_reg0 <= 36'sb111100010001110001111000100110100011;
            sine_reg0   <= 36'sb100000001101111001101110010011000001;
        end
        2997: begin
            cosine_reg0 <= 36'sb111100010100111001100110010111000100;
            sine_reg0   <= 36'sb100000001101100010011111010100010000;
        end
        2998: begin
            cosine_reg0 <= 36'sb111100011000000001010110011000100111;
            sine_reg0   <= 36'sb100000001101001011100011111100011101;
        end
        2999: begin
            cosine_reg0 <= 36'sb111100011011001001001000101001001111;
            sine_reg0   <= 36'sb100000001100110100111100001011110100;
        end
        3000: begin
            cosine_reg0 <= 36'sb111100011110010000111101000111000011;
            sine_reg0   <= 36'sb100000001100011110101000000010100110;
        end
        3001: begin
            cosine_reg0 <= 36'sb111100100001011000110011110000000111;
            sine_reg0   <= 36'sb100000001100001000100111100000111110;
        end
        3002: begin
            cosine_reg0 <= 36'sb111100100100100000101100100010011110;
            sine_reg0   <= 36'sb100000001011110010111010100111001011;
        end
        3003: begin
            cosine_reg0 <= 36'sb111100100111101000100111011100001111;
            sine_reg0   <= 36'sb100000001011011101100001010101011010;
        end
        3004: begin
            cosine_reg0 <= 36'sb111100101010110000100100011011011110;
            sine_reg0   <= 36'sb100000001011001000011011101011111000;
        end
        3005: begin
            cosine_reg0 <= 36'sb111100101101111000100011011110001111;
            sine_reg0   <= 36'sb100000001010110011101001101010110011;
        end
        3006: begin
            cosine_reg0 <= 36'sb111100110001000000100100100010100111;
            sine_reg0   <= 36'sb100000001010011111001011010010010111;
        end
        3007: begin
            cosine_reg0 <= 36'sb111100110100001000100111100110101011;
            sine_reg0   <= 36'sb100000001010001011000000100010110001;
        end
        3008: begin
            cosine_reg0 <= 36'sb111100110111010000101100101000011111;
            sine_reg0   <= 36'sb100000001001110111001001011100001101;
        end
        3009: begin
            cosine_reg0 <= 36'sb111100111010011000110011100110001000;
            sine_reg0   <= 36'sb100000001001100011100101111110110111;
        end
        3010: begin
            cosine_reg0 <= 36'sb111100111101100000111100011101101010;
            sine_reg0   <= 36'sb100000001001010000010110001010111100;
        end
        3011: begin
            cosine_reg0 <= 36'sb111101000000101001000111001101001010;
            sine_reg0   <= 36'sb100000001000111101011010000000100111;
        end
        3012: begin
            cosine_reg0 <= 36'sb111101000011110001010011110010101101;
            sine_reg0   <= 36'sb100000001000101010110001100000000101;
        end
        3013: begin
            cosine_reg0 <= 36'sb111101000110111001100010001100010111;
            sine_reg0   <= 36'sb100000001000011000011100101001011111;
        end
        3014: begin
            cosine_reg0 <= 36'sb111101001010000001110010011000001100;
            sine_reg0   <= 36'sb100000001000000110011011011101000011;
        end
        3015: begin
            cosine_reg0 <= 36'sb111101001101001010000100010100010010;
            sine_reg0   <= 36'sb100000000111110100101101111010111011;
        end
        3016: begin
            cosine_reg0 <= 36'sb111101010000010010010111111110101011;
            sine_reg0   <= 36'sb100000000111100011010100000011010010;
        end
        3017: begin
            cosine_reg0 <= 36'sb111101010011011010101101010101011110;
            sine_reg0   <= 36'sb100000000111010010001101110110010010;
        end
        3018: begin
            cosine_reg0 <= 36'sb111101010110100011000100010110101110;
            sine_reg0   <= 36'sb100000000111000001011011010100000111;
        end
        3019: begin
            cosine_reg0 <= 36'sb111101011001101011011101000000011111;
            sine_reg0   <= 36'sb100000000110110000111100011100111010;
        end
        3020: begin
            cosine_reg0 <= 36'sb111101011100110011110111010000110111;
            sine_reg0   <= 36'sb100000000110100000110001010000110101;
        end
        3021: begin
            cosine_reg0 <= 36'sb111101011111111100010011000101111001;
            sine_reg0   <= 36'sb100000000110010000111001110000000100;
        end
        3022: begin
            cosine_reg0 <= 36'sb111101100011000100110000011101101010;
            sine_reg0   <= 36'sb100000000110000001010101111010101111;
        end
        3023: begin
            cosine_reg0 <= 36'sb111101100110001101001111010110001110;
            sine_reg0   <= 36'sb100000000101110010000101110001000000;
        end
        3024: begin
            cosine_reg0 <= 36'sb111101101001010101101111101101101010;
            sine_reg0   <= 36'sb100000000101100011001001010011000001;
        end
        3025: begin
            cosine_reg0 <= 36'sb111101101100011110010001100010000001;
            sine_reg0   <= 36'sb100000000101010100100000100000111010;
        end
        3026: begin
            cosine_reg0 <= 36'sb111101101111100110110100110001011001;
            sine_reg0   <= 36'sb100000000101000110001011011010110101;
        end
        3027: begin
            cosine_reg0 <= 36'sb111101110010101111011001011001110101;
            sine_reg0   <= 36'sb100000000100111000001010000000111011;
        end
        3028: begin
            cosine_reg0 <= 36'sb111101110101110111111111011001011001;
            sine_reg0   <= 36'sb100000000100101010011100010011010011;
        end
        3029: begin
            cosine_reg0 <= 36'sb111101111001000000100110101110001011;
            sine_reg0   <= 36'sb100000000100011101000010010010001000;
        end
        3030: begin
            cosine_reg0 <= 36'sb111101111100001001001111010110001110;
            sine_reg0   <= 36'sb100000000100001111111011111101100000;
        end
        3031: begin
            cosine_reg0 <= 36'sb111101111111010001111001001111100110;
            sine_reg0   <= 36'sb100000000100000011001001010101100101;
        end
        3032: begin
            cosine_reg0 <= 36'sb111110000010011010100100011000011000;
            sine_reg0   <= 36'sb100000000011110110101010011010011101;
        end
        3033: begin
            cosine_reg0 <= 36'sb111110000101100011010000101110101000;
            sine_reg0   <= 36'sb100000000011101010011111001100010001;
        end
        3034: begin
            cosine_reg0 <= 36'sb111110001000101011111110010000011010;
            sine_reg0   <= 36'sb100000000011011110100111101011001001;
        end
        3035: begin
            cosine_reg0 <= 36'sb111110001011110100101100111011110010;
            sine_reg0   <= 36'sb100000000011010011000011110111001010;
        end
        3036: begin
            cosine_reg0 <= 36'sb111110001110111101011100101110110101;
            sine_reg0   <= 36'sb100000000011000111110011110000011110;
        end
        3037: begin
            cosine_reg0 <= 36'sb111110010010000110001101100111100110;
            sine_reg0   <= 36'sb100000000010111100110111010111001001;
        end
        3038: begin
            cosine_reg0 <= 36'sb111110010101001110111111100100001011;
            sine_reg0   <= 36'sb100000000010110010001110101011010101;
        end
        3039: begin
            cosine_reg0 <= 36'sb111110011000010111110010100010100110;
            sine_reg0   <= 36'sb100000000010100111111001101101000101;
        end
        3040: begin
            cosine_reg0 <= 36'sb111110011011100000100110100000111100;
            sine_reg0   <= 36'sb100000000010011101111000011100100011;
        end
        3041: begin
            cosine_reg0 <= 36'sb111110011110101001011011011101010001;
            sine_reg0   <= 36'sb100000000010010100001010111001110010;
        end
        3042: begin
            cosine_reg0 <= 36'sb111110100001110010010001010101101010;
            sine_reg0   <= 36'sb100000000010001010110001000100111010;
        end
        3043: begin
            cosine_reg0 <= 36'sb111110100100111011001000001000001010;
            sine_reg0   <= 36'sb100000000010000001101010111110000000;
        end
        3044: begin
            cosine_reg0 <= 36'sb111110101000000011111111110010110110;
            sine_reg0   <= 36'sb100000000001111000111000100101001010;
        end
        3045: begin
            cosine_reg0 <= 36'sb111110101011001100111000010011110001;
            sine_reg0   <= 36'sb100000000001110000011001111010011101;
        end
        3046: begin
            cosine_reg0 <= 36'sb111110101110010101110001101001000000;
            sine_reg0   <= 36'sb100000000001101000001110111101111111;
        end
        3047: begin
            cosine_reg0 <= 36'sb111110110001011110101011110000100111;
            sine_reg0   <= 36'sb100000000001100000010111101111110100;
        end
        3048: begin
            cosine_reg0 <= 36'sb111110110100100111100110101000101010;
            sine_reg0   <= 36'sb100000000001011000110100010000000001;
        end
        3049: begin
            cosine_reg0 <= 36'sb111110110111110000100010001111001100;
            sine_reg0   <= 36'sb100000000001010001100100011110101100;
        end
        3050: begin
            cosine_reg0 <= 36'sb111110111010111001011110100010010011;
            sine_reg0   <= 36'sb100000000001001010101000011011111000;
        end
        3051: begin
            cosine_reg0 <= 36'sb111110111110000010011011100000000010;
            sine_reg0   <= 36'sb100000000001000100000000000111101001;
        end
        3052: begin
            cosine_reg0 <= 36'sb111111000001001011011001000110011100;
            sine_reg0   <= 36'sb100000000000111101101011100010000101;
        end
        3053: begin
            cosine_reg0 <= 36'sb111111000100010100010111010011100111;
            sine_reg0   <= 36'sb100000000000110111101010101011001110;
        end
        3054: begin
            cosine_reg0 <= 36'sb111111000111011101010110000101100110;
            sine_reg0   <= 36'sb100000000000110001111101100011001000;
        end
        3055: begin
            cosine_reg0 <= 36'sb111111001010100110010101011010011101;
            sine_reg0   <= 36'sb100000000000101100100100001001111000;
        end
        3056: begin
            cosine_reg0 <= 36'sb111111001101101111010101010000010001;
            sine_reg0   <= 36'sb100000000000100111011110011111100000;
        end
        3057: begin
            cosine_reg0 <= 36'sb111111010000111000010101100101000100;
            sine_reg0   <= 36'sb100000000000100010101100100100000011;
        end
        3058: begin
            cosine_reg0 <= 36'sb111111010100000001010110010110111100;
            sine_reg0   <= 36'sb100000000000011110001110010111100101;
        end
        3059: begin
            cosine_reg0 <= 36'sb111111010111001010010111100011111100;
            sine_reg0   <= 36'sb100000000000011010000011111010001000;
        end
        3060: begin
            cosine_reg0 <= 36'sb111111011010010011011001001010001000;
            sine_reg0   <= 36'sb100000000000010110001101001011101110;
        end
        3061: begin
            cosine_reg0 <= 36'sb111111011101011100011011000111100101;
            sine_reg0   <= 36'sb100000000000010010101010001100011011;
        end
        3062: begin
            cosine_reg0 <= 36'sb111111100000100101011101011010010101;
            sine_reg0   <= 36'sb100000000000001111011010111100010000;
        end
        3063: begin
            cosine_reg0 <= 36'sb111111100011101110100000000000011110;
            sine_reg0   <= 36'sb100000000000001100011111011011001111;
        end
        3064: begin
            cosine_reg0 <= 36'sb111111100110110111100010111000000011;
            sine_reg0   <= 36'sb100000000000001001110111101001011010;
        end
        3065: begin
            cosine_reg0 <= 36'sb111111101010000000100101111111001000;
            sine_reg0   <= 36'sb100000000000000111100011100110110011;
        end
        3066: begin
            cosine_reg0 <= 36'sb111111101101001001101001010011110010;
            sine_reg0   <= 36'sb100000000000000101100011010011011011;
        end
        3067: begin
            cosine_reg0 <= 36'sb111111110000010010101100110100000011;
            sine_reg0   <= 36'sb100000000000000011110110101111010100;
        end
        3068: begin
            cosine_reg0 <= 36'sb111111110011011011110000011110000001;
            sine_reg0   <= 36'sb100000000000000010011101111010011101;
        end
        3069: begin
            cosine_reg0 <= 36'sb111111110110100100110100001111101111;
            sine_reg0   <= 36'sb100000000000000001011000110100111001;
        end
        3070: begin
            cosine_reg0 <= 36'sb111111111001101101111000000111010000;
            sine_reg0   <= 36'sb100000000000000000100111011110101000;
        end
        3071: begin
            cosine_reg0 <= 36'sb111111111100110110111100000010101010;
            sine_reg0   <= 36'sb100000000000000000001001110111101011;
        end
        3072: begin
            cosine_reg0 <= 36'sb0;
            sine_reg0   <= 36'sb100000000000000000000000000000000001;
        end
        3073: begin
            cosine_reg0 <= 36'sb11001001000011111101010110;
            sine_reg0   <= 36'sb100000000000000000001001110111101011;
        end
        3074: begin
            cosine_reg0 <= 36'sb110010010000111111000110000;
            sine_reg0   <= 36'sb100000000000000000100111011110101000;
        end
        3075: begin
            cosine_reg0 <= 36'sb1001011011001011110000010001;
            sine_reg0   <= 36'sb100000000000000001011000110100111001;
        end
        3076: begin
            cosine_reg0 <= 36'sb1100100100001111100001111111;
            sine_reg0   <= 36'sb100000000000000010011101111010011101;
        end
        3077: begin
            cosine_reg0 <= 36'sb1111101101010011001011111101;
            sine_reg0   <= 36'sb100000000000000011110110101111010100;
        end
        3078: begin
            cosine_reg0 <= 36'sb10010110110010110101100001110;
            sine_reg0   <= 36'sb100000000000000101100011010011011011;
        end
        3079: begin
            cosine_reg0 <= 36'sb10101111111011010000000111000;
            sine_reg0   <= 36'sb100000000000000111100011100110110011;
        end
        3080: begin
            cosine_reg0 <= 36'sb11001001000011101000111111101;
            sine_reg0   <= 36'sb100000000000001001110111101001011010;
        end
        3081: begin
            cosine_reg0 <= 36'sb11100010001011111111111100010;
            sine_reg0   <= 36'sb100000000000001100011111011011001111;
        end
        3082: begin
            cosine_reg0 <= 36'sb11111011010100010100101101011;
            sine_reg0   <= 36'sb100000000000001111011010111100010000;
        end
        3083: begin
            cosine_reg0 <= 36'sb100010100011100100111000011011;
            sine_reg0   <= 36'sb100000000000010010101010001100011011;
        end
        3084: begin
            cosine_reg0 <= 36'sb100101101100100110110101111000;
            sine_reg0   <= 36'sb100000000000010110001101001011101110;
        end
        3085: begin
            cosine_reg0 <= 36'sb101000110101101000011100000100;
            sine_reg0   <= 36'sb100000000000011010000011111010001000;
        end
        3086: begin
            cosine_reg0 <= 36'sb101011111110101001101001000100;
            sine_reg0   <= 36'sb100000000000011110001110010111100101;
        end
        3087: begin
            cosine_reg0 <= 36'sb101111000111101010011010111100;
            sine_reg0   <= 36'sb100000000000100010101100100100000011;
        end
        3088: begin
            cosine_reg0 <= 36'sb110010010000101010101111101111;
            sine_reg0   <= 36'sb100000000000100111011110011111100000;
        end
        3089: begin
            cosine_reg0 <= 36'sb110101011001101010100101100011;
            sine_reg0   <= 36'sb100000000000101100100100001001111000;
        end
        3090: begin
            cosine_reg0 <= 36'sb111000100010101001111010011010;
            sine_reg0   <= 36'sb100000000000110001111101100011001000;
        end
        3091: begin
            cosine_reg0 <= 36'sb111011101011101000101100011001;
            sine_reg0   <= 36'sb100000000000110111101010101011001110;
        end
        3092: begin
            cosine_reg0 <= 36'sb111110110100100110111001100100;
            sine_reg0   <= 36'sb100000000000111101101011100010000101;
        end
        3093: begin
            cosine_reg0 <= 36'sb1000001111101100100011111111110;
            sine_reg0   <= 36'sb100000000001000100000000000111101001;
        end
        3094: begin
            cosine_reg0 <= 36'sb1000101000110100001011101101101;
            sine_reg0   <= 36'sb100000000001001010101000011011111000;
        end
        3095: begin
            cosine_reg0 <= 36'sb1001000001111011101110000110100;
            sine_reg0   <= 36'sb100000000001010001100100011110101100;
        end
        3096: begin
            cosine_reg0 <= 36'sb1001011011000011001010111010110;
            sine_reg0   <= 36'sb100000000001011000110100010000000001;
        end
        3097: begin
            cosine_reg0 <= 36'sb1001110100001010100001111011001;
            sine_reg0   <= 36'sb100000000001100000010111101111110100;
        end
        3098: begin
            cosine_reg0 <= 36'sb1010001101010001110010111000000;
            sine_reg0   <= 36'sb100000000001101000001110111101111111;
        end
        3099: begin
            cosine_reg0 <= 36'sb1010100110011000111101100001111;
            sine_reg0   <= 36'sb100000000001110000011001111010011101;
        end
        3100: begin
            cosine_reg0 <= 36'sb1010111111100000000001101001010;
            sine_reg0   <= 36'sb100000000001111000111000100101001010;
        end
        3101: begin
            cosine_reg0 <= 36'sb1011011000100110111110111110110;
            sine_reg0   <= 36'sb100000000010000001101010111110000000;
        end
        3102: begin
            cosine_reg0 <= 36'sb1011110001101101110101010010110;
            sine_reg0   <= 36'sb100000000010001010110001000100111010;
        end
        3103: begin
            cosine_reg0 <= 36'sb1100001010110100100100010101111;
            sine_reg0   <= 36'sb100000000010010100001010111001110010;
        end
        3104: begin
            cosine_reg0 <= 36'sb1100100011111011001011111000100;
            sine_reg0   <= 36'sb100000000010011101111000011100100011;
        end
        3105: begin
            cosine_reg0 <= 36'sb1100111101000001101011101011010;
            sine_reg0   <= 36'sb100000000010100111111001101101000101;
        end
        3106: begin
            cosine_reg0 <= 36'sb1101010110001000000011011110101;
            sine_reg0   <= 36'sb100000000010110010001110101011010101;
        end
        3107: begin
            cosine_reg0 <= 36'sb1101101111001110010011000011010;
            sine_reg0   <= 36'sb100000000010111100110111010111001001;
        end
        3108: begin
            cosine_reg0 <= 36'sb1110001000010100011010001001011;
            sine_reg0   <= 36'sb100000000011000111110011110000011110;
        end
        3109: begin
            cosine_reg0 <= 36'sb1110100001011010011000100001110;
            sine_reg0   <= 36'sb100000000011010011000011110111001010;
        end
        3110: begin
            cosine_reg0 <= 36'sb1110111010100000001101111100110;
            sine_reg0   <= 36'sb100000000011011110100111101011001001;
        end
        3111: begin
            cosine_reg0 <= 36'sb1111010011100101111010001011000;
            sine_reg0   <= 36'sb100000000011101010011111001100010001;
        end
        3112: begin
            cosine_reg0 <= 36'sb1111101100101011011100111101000;
            sine_reg0   <= 36'sb100000000011110110101010011010011101;
        end
        3113: begin
            cosine_reg0 <= 36'sb10000000101110000110110000011010;
            sine_reg0   <= 36'sb100000000100000011001001010101100101;
        end
        3114: begin
            cosine_reg0 <= 36'sb10000011110110110000101001110010;
            sine_reg0   <= 36'sb100000000100001111111011111101100000;
        end
        3115: begin
            cosine_reg0 <= 36'sb10000110111111011001010001110101;
            sine_reg0   <= 36'sb100000000100011101000010010010001000;
        end
        3116: begin
            cosine_reg0 <= 36'sb10001010001000000000100110100111;
            sine_reg0   <= 36'sb100000000100101010011100010011010011;
        end
        3117: begin
            cosine_reg0 <= 36'sb10001101010000100110100110001011;
            sine_reg0   <= 36'sb100000000100111000001010000000111011;
        end
        3118: begin
            cosine_reg0 <= 36'sb10010000011001001011001110100111;
            sine_reg0   <= 36'sb100000000101000110001011011010110101;
        end
        3119: begin
            cosine_reg0 <= 36'sb10010011100001101110011101111111;
            sine_reg0   <= 36'sb100000000101010100100000100000111010;
        end
        3120: begin
            cosine_reg0 <= 36'sb10010110101010010000010010010110;
            sine_reg0   <= 36'sb100000000101100011001001010011000001;
        end
        3121: begin
            cosine_reg0 <= 36'sb10011001110010110000101001110010;
            sine_reg0   <= 36'sb100000000101110010000101110001000000;
        end
        3122: begin
            cosine_reg0 <= 36'sb10011100111011001111100010010110;
            sine_reg0   <= 36'sb100000000110000001010101111010101111;
        end
        3123: begin
            cosine_reg0 <= 36'sb10100000000011101100111010000111;
            sine_reg0   <= 36'sb100000000110010000111001110000000100;
        end
        3124: begin
            cosine_reg0 <= 36'sb10100011001100001000101111001001;
            sine_reg0   <= 36'sb100000000110100000110001010000110101;
        end
        3125: begin
            cosine_reg0 <= 36'sb10100110010100100010111111100001;
            sine_reg0   <= 36'sb100000000110110000111100011100111010;
        end
        3126: begin
            cosine_reg0 <= 36'sb10101001011100111011101001010010;
            sine_reg0   <= 36'sb100000000111000001011011010100000111;
        end
        3127: begin
            cosine_reg0 <= 36'sb10101100100101010010101010100010;
            sine_reg0   <= 36'sb100000000111010010001101110110010010;
        end
        3128: begin
            cosine_reg0 <= 36'sb10101111101101101000000001010101;
            sine_reg0   <= 36'sb100000000111100011010100000011010010;
        end
        3129: begin
            cosine_reg0 <= 36'sb10110010110101111011101011101110;
            sine_reg0   <= 36'sb100000000111110100101101111010111011;
        end
        3130: begin
            cosine_reg0 <= 36'sb10110101111110001101100111110100;
            sine_reg0   <= 36'sb100000001000000110011011011101000011;
        end
        3131: begin
            cosine_reg0 <= 36'sb10111001000110011101110011101001;
            sine_reg0   <= 36'sb100000001000011000011100101001011111;
        end
        3132: begin
            cosine_reg0 <= 36'sb10111100001110101100001101010011;
            sine_reg0   <= 36'sb100000001000101010110001100000000101;
        end
        3133: begin
            cosine_reg0 <= 36'sb10111111010110111000110010110110;
            sine_reg0   <= 36'sb100000001000111101011010000000100111;
        end
        3134: begin
            cosine_reg0 <= 36'sb11000010011111000011100010010110;
            sine_reg0   <= 36'sb100000001001010000010110001010111100;
        end
        3135: begin
            cosine_reg0 <= 36'sb11000101100111001100011001111000;
            sine_reg0   <= 36'sb100000001001100011100101111110110111;
        end
        3136: begin
            cosine_reg0 <= 36'sb11001000101111010011010111100001;
            sine_reg0   <= 36'sb100000001001110111001001011100001101;
        end
        3137: begin
            cosine_reg0 <= 36'sb11001011110111011000011001010101;
            sine_reg0   <= 36'sb100000001010001011000000100010110001;
        end
        3138: begin
            cosine_reg0 <= 36'sb11001110111111011011011101011001;
            sine_reg0   <= 36'sb100000001010011111001011010010010111;
        end
        3139: begin
            cosine_reg0 <= 36'sb11010010000111011100100001110001;
            sine_reg0   <= 36'sb100000001010110011101001101010110011;
        end
        3140: begin
            cosine_reg0 <= 36'sb11010101001111011011100100100010;
            sine_reg0   <= 36'sb100000001011001000011011101011111000;
        end
        3141: begin
            cosine_reg0 <= 36'sb11011000010111011000100011110001;
            sine_reg0   <= 36'sb100000001011011101100001010101011010;
        end
        3142: begin
            cosine_reg0 <= 36'sb11011011011111010011011101100010;
            sine_reg0   <= 36'sb100000001011110010111010100111001011;
        end
        3143: begin
            cosine_reg0 <= 36'sb11011110100111001100001111111001;
            sine_reg0   <= 36'sb100000001100001000100111100000111110;
        end
        3144: begin
            cosine_reg0 <= 36'sb11100001101111000010111000111101;
            sine_reg0   <= 36'sb100000001100011110101000000010100110;
        end
        3145: begin
            cosine_reg0 <= 36'sb11100100110110110111010110110001;
            sine_reg0   <= 36'sb100000001100110100111100001011110100;
        end
        3146: begin
            cosine_reg0 <= 36'sb11100111111110101001100111011001;
            sine_reg0   <= 36'sb100000001101001011100011111100011101;
        end
        3147: begin
            cosine_reg0 <= 36'sb11101011000110011001101000111100;
            sine_reg0   <= 36'sb100000001101100010011111010100010000;
        end
        3148: begin
            cosine_reg0 <= 36'sb11101110001110000111011001011101;
            sine_reg0   <= 36'sb100000001101111001101110010011000001;
        end
        3149: begin
            cosine_reg0 <= 36'sb11110001010101110010110111000010;
            sine_reg0   <= 36'sb100000001110010001010000111000100001;
        end
        3150: begin
            cosine_reg0 <= 36'sb11110100011101011011111111101111;
            sine_reg0   <= 36'sb100000001110101001000111000100100010;
        end
        3151: begin
            cosine_reg0 <= 36'sb11110111100101000010110001101001;
            sine_reg0   <= 36'sb100000001111000001010000110110110100;
        end
        3152: begin
            cosine_reg0 <= 36'sb11111010101100100111001010110101;
            sine_reg0   <= 36'sb100000001111011001101110001111001001;
        end
        3153: begin
            cosine_reg0 <= 36'sb11111101110100001001001001011000;
            sine_reg0   <= 36'sb100000001111110010011111001101010001;
        end
        3154: begin
            cosine_reg0 <= 36'sb100000000111011101000101011010111;
            sine_reg0   <= 36'sb100000010000001011100011110000111110;
        end
        3155: begin
            cosine_reg0 <= 36'sb100000100000011000101101110110110;
            sine_reg0   <= 36'sb100000010000100100111011111010000000;
        end
        3156: begin
            cosine_reg0 <= 36'sb100000111001010100000010001111100;
            sine_reg0   <= 36'sb100000010000111110100111101000001000;
        end
        3157: begin
            cosine_reg0 <= 36'sb100001010010001111000010010101011;
            sine_reg0   <= 36'sb100000010001011000100110111011000101;
        end
        3158: begin
            cosine_reg0 <= 36'sb100001101011001001101101111001011;
            sine_reg0   <= 36'sb100000010001110010111001110010100111;
        end
        3159: begin
            cosine_reg0 <= 36'sb100010000100000100000100101011111;
            sine_reg0   <= 36'sb100000010010001101100000001110011111;
        end
        3160: begin
            cosine_reg0 <= 36'sb100010011100111110000110011101110;
            sine_reg0   <= 36'sb100000010010101000011010001110011100;
        end
        3161: begin
            cosine_reg0 <= 36'sb100010110101110111110010111111011;
            sine_reg0   <= 36'sb100000010011000011100111110010001100;
        end
        3162: begin
            cosine_reg0 <= 36'sb100011001110110001001010000001100;
            sine_reg0   <= 36'sb100000010011011111001000111001100001;
        end
        3163: begin
            cosine_reg0 <= 36'sb100011100111101010001011010100110;
            sine_reg0   <= 36'sb100000010011111010111101100100000111;
        end
        3164: begin
            cosine_reg0 <= 36'sb100100000000100010110110101001111;
            sine_reg0   <= 36'sb100000010100010111000101110001101111;
        end
        3165: begin
            cosine_reg0 <= 36'sb100100011001011011001011110001011;
            sine_reg0   <= 36'sb100000010100110011100001100010000111;
        end
        3166: begin
            cosine_reg0 <= 36'sb100100110010010011001010011100000;
            sine_reg0   <= 36'sb100000010101010000010000110100111110;
        end
        3167: begin
            cosine_reg0 <= 36'sb100101001011001010110010011010011;
            sine_reg0   <= 36'sb100000010101101101010011101010000001;
        end
        3168: begin
            cosine_reg0 <= 36'sb100101100100000010000011011101001;
            sine_reg0   <= 36'sb100000010110001010101010000000111111;
        end
        3169: begin
            cosine_reg0 <= 36'sb100101111100111000111101010101000;
            sine_reg0   <= 36'sb100000010110101000010011111001100101;
        end
        3170: begin
            cosine_reg0 <= 36'sb100110010101101111011111110010100;
            sine_reg0   <= 36'sb100000010111000110010001010011100010;
        end
        3171: begin
            cosine_reg0 <= 36'sb100110101110100101101010100110100;
            sine_reg0   <= 36'sb100000010111100100100010001110100011;
        end
        3172: begin
            cosine_reg0 <= 36'sb100111000111011011011101100001101;
            sine_reg0   <= 36'sb100000011000000011000110101010010110;
        end
        3173: begin
            cosine_reg0 <= 36'sb100111100000010000111000010100011;
            sine_reg0   <= 36'sb100000011000100001111110100110100110;
        end
        3174: begin
            cosine_reg0 <= 36'sb100111111001000101111010101111110;
            sine_reg0   <= 36'sb100000011001000001001010000011000010;
        end
        3175: begin
            cosine_reg0 <= 36'sb101000010001111010100100100100001;
            sine_reg0   <= 36'sb100000011001100000101000111111010110;
        end
        3176: begin
            cosine_reg0 <= 36'sb101000101010101110110101100010010;
            sine_reg0   <= 36'sb100000011010000000011011011011001111;
        end
        3177: begin
            cosine_reg0 <= 36'sb101001000011100010101101011011000;
            sine_reg0   <= 36'sb100000011010100000100001010110011001;
        end
        3178: begin
            cosine_reg0 <= 36'sb101001011100010110001011111110111;
            sine_reg0   <= 36'sb100000011011000000111010110000100000;
        end
        3179: begin
            cosine_reg0 <= 36'sb101001110101001001010000111110110;
            sine_reg0   <= 36'sb100000011011100001100111101001010000;
        end
        3180: begin
            cosine_reg0 <= 36'sb101010001101111011111100001011001;
            sine_reg0   <= 36'sb100000011100000010101000000000010101;
        end
        3181: begin
            cosine_reg0 <= 36'sb101010100110101110001101010100111;
            sine_reg0   <= 36'sb100000011100100011111011110101011100;
        end
        3182: begin
            cosine_reg0 <= 36'sb101010111111100000000100001100101;
            sine_reg0   <= 36'sb100000011101000101100011001000001110;
        end
        3183: begin
            cosine_reg0 <= 36'sb101011011000010001100000100011001;
            sine_reg0   <= 36'sb100000011101100111011101111000011000;
        end
        3184: begin
            cosine_reg0 <= 36'sb101011110001000010100010001001001;
            sine_reg0   <= 36'sb100000011110001001101100000101100101;
        end
        3185: begin
            cosine_reg0 <= 36'sb101100001001110011001000101111001;
            sine_reg0   <= 36'sb100000011110101100001101101111011111;
        end
        3186: begin
            cosine_reg0 <= 36'sb101100100010100011010100000110010;
            sine_reg0   <= 36'sb100000011111001111000010110101110001;
        end
        3187: begin
            cosine_reg0 <= 36'sb101100111011010011000011111110111;
            sine_reg0   <= 36'sb100000011111110010001011011000000110;
        end
        3188: begin
            cosine_reg0 <= 36'sb101101010100000010011000001001111;
            sine_reg0   <= 36'sb100000100000010101100111010110000111;
        end
        3189: begin
            cosine_reg0 <= 36'sb101101101100110001010000011000000;
            sine_reg0   <= 36'sb100000100000111001010110101111100000;
        end
        3190: begin
            cosine_reg0 <= 36'sb101110000101011111101100011010000;
            sine_reg0   <= 36'sb100000100001011101011001100011111010;
        end
        3191: begin
            cosine_reg0 <= 36'sb101110011110001101101100000000101;
            sine_reg0   <= 36'sb100000100010000001101111110010111111;
        end
        3192: begin
            cosine_reg0 <= 36'sb101110110110111011001110111100101;
            sine_reg0   <= 36'sb100000100010100110011001011100011001;
        end
        3193: begin
            cosine_reg0 <= 36'sb101111001111101000010100111110101;
            sine_reg0   <= 36'sb100000100011001011010110011111110000;
        end
        3194: begin
            cosine_reg0 <= 36'sb101111101000010100111101110111101;
            sine_reg0   <= 36'sb100000100011110000100110111100101110;
        end
        3195: begin
            cosine_reg0 <= 36'sb110000000001000001001001011000010;
            sine_reg0   <= 36'sb100000100100010110001010110010111100;
        end
        3196: begin
            cosine_reg0 <= 36'sb110000011001101100110111010001010;
            sine_reg0   <= 36'sb100000100100111100000010000010000100;
        end
        3197: begin
            cosine_reg0 <= 36'sb110000110010011000000111010011011;
            sine_reg0   <= 36'sb100000100101100010001100101001101100;
        end
        3198: begin
            cosine_reg0 <= 36'sb110001001011000010111001001111100;
            sine_reg0   <= 36'sb100000100110001000101010101001011111;
        end
        3199: begin
            cosine_reg0 <= 36'sb110001100011101101001100110110011;
            sine_reg0   <= 36'sb100000100110101111011100000001000100;
        end
        3200: begin
            cosine_reg0 <= 36'sb110001111100010111000001111000110;
            sine_reg0   <= 36'sb100000100111010110100000110000000011;
        end
        3201: begin
            cosine_reg0 <= 36'sb110010010101000000011000000111100;
            sine_reg0   <= 36'sb100000100111111101111000110110000101;
        end
        3202: begin
            cosine_reg0 <= 36'sb110010101101101001001111010011011;
            sine_reg0   <= 36'sb100000101000100101100100010010110000;
        end
        3203: begin
            cosine_reg0 <= 36'sb110011000110010001100111001101001;
            sine_reg0   <= 36'sb100000101001001101100011000101101101;
        end
        3204: begin
            cosine_reg0 <= 36'sb110011011110111001011111100101110;
            sine_reg0   <= 36'sb100000101001110101110101001110100011;
        end
        3205: begin
            cosine_reg0 <= 36'sb110011110111100000111000001101110;
            sine_reg0   <= 36'sb100000101010011110011010101100111001;
        end
        3206: begin
            cosine_reg0 <= 36'sb110100010000000111110000110110001;
            sine_reg0   <= 36'sb100000101011000111010011100000010101;
        end
        3207: begin
            cosine_reg0 <= 36'sb110100101000101110001001001111110;
            sine_reg0   <= 36'sb100000101011110000011111101000100000;
        end
        3208: begin
            cosine_reg0 <= 36'sb110101000001010100000001001011011;
            sine_reg0   <= 36'sb100000101100011001111111000100111110;
        end
        3209: begin
            cosine_reg0 <= 36'sb110101011001111001011000011001110;
            sine_reg0   <= 36'sb100000101101000011110001110101011000;
        end
        3210: begin
            cosine_reg0 <= 36'sb110101110010011110001110101011111;
            sine_reg0   <= 36'sb100000101101101101110111111001010010;
        end
        3211: begin
            cosine_reg0 <= 36'sb110110001011000010100011110010100;
            sine_reg0   <= 36'sb100000101110011000010001010000010011;
        end
        3212: begin
            cosine_reg0 <= 36'sb110110100011100110010111011110100;
            sine_reg0   <= 36'sb100000101111000010111101111010000001;
        end
        3213: begin
            cosine_reg0 <= 36'sb110110111100001001101001100000101;
            sine_reg0   <= 36'sb100000101111101101111101110110000010;
        end
        3214: begin
            cosine_reg0 <= 36'sb110111010100101100011001101001111;
            sine_reg0   <= 36'sb100000110000011001010001000011111010;
        end
        3215: begin
            cosine_reg0 <= 36'sb110111101101001110100111101011000;
            sine_reg0   <= 36'sb100000110001000100110111100011010000;
        end
        3216: begin
            cosine_reg0 <= 36'sb111000000101110000010011010101000;
            sine_reg0   <= 36'sb100000110001110000110001010011101000;
        end
        3217: begin
            cosine_reg0 <= 36'sb111000011110010001011100011000101;
            sine_reg0   <= 36'sb100000110010011100111110010100100111;
        end
        3218: begin
            cosine_reg0 <= 36'sb111000110110110010000010100110110;
            sine_reg0   <= 36'sb100000110011001001011110100101110010;
        end
        3219: begin
            cosine_reg0 <= 36'sb111001001111010010000101110000010;
            sine_reg0   <= 36'sb100000110011110110010010000110101110;
        end
        3220: begin
            cosine_reg0 <= 36'sb111001100111110001100101100110001;
            sine_reg0   <= 36'sb100000110100100011011000110110111111;
        end
        3221: begin
            cosine_reg0 <= 36'sb111010000000010000100001111001001;
            sine_reg0   <= 36'sb100000110101010000110010110110001001;
        end
        3222: begin
            cosine_reg0 <= 36'sb111010011000101110111010011010011;
            sine_reg0   <= 36'sb100000110101111110100000000011101111;
        end
        3223: begin
            cosine_reg0 <= 36'sb111010110001001100101110111010100;
            sine_reg0   <= 36'sb100000110110101100100000011111010111;
        end
        3224: begin
            cosine_reg0 <= 36'sb111011001001101001111111001010100;
            sine_reg0   <= 36'sb100000110111011010110100001000100011;
        end
        3225: begin
            cosine_reg0 <= 36'sb111011100010000110101010111011011;
            sine_reg0   <= 36'sb100000111000001001011010111110111000;
        end
        3226: begin
            cosine_reg0 <= 36'sb111011111010100010110001111110000;
            sine_reg0   <= 36'sb100000111000111000010101000001110111;
        end
        3227: begin
            cosine_reg0 <= 36'sb111100010010111110010100000011010;
            sine_reg0   <= 36'sb100000111001100111100010010001000100;
        end
        3228: begin
            cosine_reg0 <= 36'sb111100101011011001010000111100001;
            sine_reg0   <= 36'sb100000111010010111000010101100000011;
        end
        3229: begin
            cosine_reg0 <= 36'sb111101000011110011101000011001100;
            sine_reg0   <= 36'sb100000111011000110110110010010010110;
        end
        3230: begin
            cosine_reg0 <= 36'sb111101011100001101011010001100011;
            sine_reg0   <= 36'sb100000111011110110111101000011011111;
        end
        3231: begin
            cosine_reg0 <= 36'sb111101110100100110100110000101101;
            sine_reg0   <= 36'sb100000111100100111010110111111000000;
        end
        3232: begin
            cosine_reg0 <= 36'sb111110001100111111001011110110010;
            sine_reg0   <= 36'sb100000111101011000000100000100011100;
        end
        3233: begin
            cosine_reg0 <= 36'sb111110100101010111001011001111010;
            sine_reg0   <= 36'sb100000111110001001000100010011010101;
        end
        3234: begin
            cosine_reg0 <= 36'sb111110111101101110100100000001100;
            sine_reg0   <= 36'sb100000111110111010010111101011001101;
        end
        3235: begin
            cosine_reg0 <= 36'sb111111010110000101010101111110000;
            sine_reg0   <= 36'sb100000111111101011111110001011100101;
        end
        3236: begin
            cosine_reg0 <= 36'sb111111101110011011100000110101110;
            sine_reg0   <= 36'sb100001000000011101110111110011111110;
        end
        3237: begin
            cosine_reg0 <= 36'sb1000000000110110001000100011001110;
            sine_reg0   <= 36'sb100001000001010000000100100011111010;
        end
        3238: begin
            cosine_reg0 <= 36'sb1000000011111000110000000011010111;
            sine_reg0   <= 36'sb100001000010000010100100011010111010;
        end
        3239: begin
            cosine_reg0 <= 36'sb1000000110111011010010100101010010;
            sine_reg0   <= 36'sb100001000010110101010111011000011110;
        end
        3240: begin
            cosine_reg0 <= 36'sb1000001001111101110000000111000111;
            sine_reg0   <= 36'sb100001000011101000011101011100001000;
        end
        3241: begin
            cosine_reg0 <= 36'sb1000001101000000001000100110111101;
            sine_reg0   <= 36'sb100001000100011011110110100101010111;
        end
        3242: begin
            cosine_reg0 <= 36'sb1000010000000010011100000010111101;
            sine_reg0   <= 36'sb100001000101001111100010110011101101;
        end
        3243: begin
            cosine_reg0 <= 36'sb1000010011000100101010011001001111;
            sine_reg0   <= 36'sb100001000110000011100010000110101001;
        end
        3244: begin
            cosine_reg0 <= 36'sb1000010110000110110011100111111011;
            sine_reg0   <= 36'sb100001000110110111110100011101101010;
        end
        3245: begin
            cosine_reg0 <= 36'sb1000011001001000110111101101001010;
            sine_reg0   <= 36'sb100001000111101100011001111000010010;
        end
        3246: begin
            cosine_reg0 <= 36'sb1000011100001010110110100111000011;
            sine_reg0   <= 36'sb100001001000100001010010010101111111;
        end
        3247: begin
            cosine_reg0 <= 36'sb1000011111001100110000010011101111;
            sine_reg0   <= 36'sb100001001001010110011101110110010001;
        end
        3248: begin
            cosine_reg0 <= 36'sb1000100010001110100100110001010110;
            sine_reg0   <= 36'sb100001001010001011111100011000100111;
        end
        3249: begin
            cosine_reg0 <= 36'sb1000100101010000010011111110000001;
            sine_reg0   <= 36'sb100001001011000001101101111100100000;
        end
        3250: begin
            cosine_reg0 <= 36'sb1000101000010001111101110111111001;
            sine_reg0   <= 36'sb100001001011110111110010100001011011;
        end
        3251: begin
            cosine_reg0 <= 36'sb1000101011010011100010011101000101;
            sine_reg0   <= 36'sb100001001100101110001010000110110110;
        end
        3252: begin
            cosine_reg0 <= 36'sb1000101110010101000001101011101111;
            sine_reg0   <= 36'sb100001001101100100110100101100010000;
        end
        3253: begin
            cosine_reg0 <= 36'sb1000110001010110011011100001111110;
            sine_reg0   <= 36'sb100001001110011011110010010001000111;
        end
        3254: begin
            cosine_reg0 <= 36'sb1000110100010111101111111101111101;
            sine_reg0   <= 36'sb100001001111010011000010110100111010;
        end
        3255: begin
            cosine_reg0 <= 36'sb1000110111011000111110111101110011;
            sine_reg0   <= 36'sb100001010000001010100110010111000110;
        end
        3256: begin
            cosine_reg0 <= 36'sb1000111010011010001000011111101001;
            sine_reg0   <= 36'sb100001010001000010011100110111001001;
        end
        3257: begin
            cosine_reg0 <= 36'sb1000111101011011001100100001101001;
            sine_reg0   <= 36'sb100001010001111010100110010100100001;
        end
        3258: begin
            cosine_reg0 <= 36'sb1001000000011100001011000001111011;
            sine_reg0   <= 36'sb100001010010110011000010101110101010;
        end
        3259: begin
            cosine_reg0 <= 36'sb1001000011011101000011111110100111;
            sine_reg0   <= 36'sb100001010011101011110010000101000011;
        end
        3260: begin
            cosine_reg0 <= 36'sb1001000110011101110111010101111000;
            sine_reg0   <= 36'sb100001010100100100110100010111000111;
        end
        3261: begin
            cosine_reg0 <= 36'sb1001001001011110100101000101110110;
            sine_reg0   <= 36'sb100001010101011110001001100100010100;
        end
        3262: begin
            cosine_reg0 <= 36'sb1001001100011111001101001100101010;
            sine_reg0   <= 36'sb100001010110010111110001101100000111;
        end
        3263: begin
            cosine_reg0 <= 36'sb1001001111011111101111101000011110;
            sine_reg0   <= 36'sb100001010111010001101100101101111100;
        end
        3264: begin
            cosine_reg0 <= 36'sb1001010010100000001100010111011010;
            sine_reg0   <= 36'sb100001011000001011111010101001001111;
        end
        3265: begin
            cosine_reg0 <= 36'sb1001010101100000100011010111101001;
            sine_reg0   <= 36'sb100001011001000110011011011101011101;
        end
        3266: begin
            cosine_reg0 <= 36'sb1001011000100000110100100111010010;
            sine_reg0   <= 36'sb100001011010000001001111001010000001;
        end
        3267: begin
            cosine_reg0 <= 36'sb1001011011100001000000000100100001;
            sine_reg0   <= 36'sb100001011010111100010101101110010110;
        end
        3268: begin
            cosine_reg0 <= 36'sb1001011110100001000101101101011101;
            sine_reg0   <= 36'sb100001011011110111101111001001111001;
        end
        3269: begin
            cosine_reg0 <= 36'sb1001100001100001000101100000010001;
            sine_reg0   <= 36'sb100001011100110011011011011100000110;
        end
        3270: begin
            cosine_reg0 <= 36'sb1001100100100000111111011011000111;
            sine_reg0   <= 36'sb100001011101101111011010100100010110;
        end
        3271: begin
            cosine_reg0 <= 36'sb1001100111100000110011011100000111;
            sine_reg0   <= 36'sb100001011110101011101100100010000101;
        end
        3272: begin
            cosine_reg0 <= 36'sb1001101010100000100001100001011100;
            sine_reg0   <= 36'sb100001011111101000010001010100101110;
        end
        3273: begin
            cosine_reg0 <= 36'sb1001101101100000001001101001001111;
            sine_reg0   <= 36'sb100001100000100101001000111011101011;
        end
        3274: begin
            cosine_reg0 <= 36'sb1001110000011111101011110001101010;
            sine_reg0   <= 36'sb100001100001100010010011010110011000;
        end
        3275: begin
            cosine_reg0 <= 36'sb1001110011011111000111111000110111;
            sine_reg0   <= 36'sb100001100010011111110000100100001101;
        end
        3276: begin
            cosine_reg0 <= 36'sb1001110110011110011101111101000000;
            sine_reg0   <= 36'sb100001100011011101100000100100100110;
        end
        3277: begin
            cosine_reg0 <= 36'sb1001111001011101101101111100001111;
            sine_reg0   <= 36'sb100001100100011011100011010110111100;
        end
        3278: begin
            cosine_reg0 <= 36'sb1001111100011100110111110100101110;
            sine_reg0   <= 36'sb100001100101011001111000111010101010;
        end
        3279: begin
            cosine_reg0 <= 36'sb1001111111011011111011100100100110;
            sine_reg0   <= 36'sb100001100110011000100001001111000111;
        end
        3280: begin
            cosine_reg0 <= 36'sb1010000010011010111001001010000011;
            sine_reg0   <= 36'sb100001100111010111011100010011101111;
        end
        3281: begin
            cosine_reg0 <= 36'sb1010000101011001110000100011001101;
            sine_reg0   <= 36'sb100001101000010110101010000111111001;
        end
        3282: begin
            cosine_reg0 <= 36'sb1010001000011000100001101110010001;
            sine_reg0   <= 36'sb100001101001010110001010101011000000;
        end
        3283: begin
            cosine_reg0 <= 36'sb1010001011010111001100101001010111;
            sine_reg0   <= 36'sb100001101010010101111101111100011011;
        end
        3284: begin
            cosine_reg0 <= 36'sb1010001110010101110001010010101011;
            sine_reg0   <= 36'sb100001101011010110000011111011100100;
        end
        3285: begin
            cosine_reg0 <= 36'sb1010010001010100001111101000010110;
            sine_reg0   <= 36'sb100001101100010110011100100111110011;
        end
        3286: begin
            cosine_reg0 <= 36'sb1010010100010010100111101000100011;
            sine_reg0   <= 36'sb100001101101010111001000000000100000;
        end
        3287: begin
            cosine_reg0 <= 36'sb1010010111010000111001010001011101;
            sine_reg0   <= 36'sb100001101110011000000110000101000100;
        end
        3288: begin
            cosine_reg0 <= 36'sb1010011010001111000100100001001111;
            sine_reg0   <= 36'sb100001101111011001010110110100110110;
        end
        3289: begin
            cosine_reg0 <= 36'sb1010011101001101001001010110000010;
            sine_reg0   <= 36'sb100001110000011010111010001111001110;
        end
        3290: begin
            cosine_reg0 <= 36'sb1010100000001011000111101110000011;
            sine_reg0   <= 36'sb100001110001011100110000010011100011;
        end
        3291: begin
            cosine_reg0 <= 36'sb1010100011001000111111100111011011;
            sine_reg0   <= 36'sb100001110010011110111001000001001110;
        end
        3292: begin
            cosine_reg0 <= 36'sb1010100110000110110001000000010110;
            sine_reg0   <= 36'sb100001110011100001010100010111100101;
        end
        3293: begin
            cosine_reg0 <= 36'sb1010101001000100011011110110111110;
            sine_reg0   <= 36'sb100001110100100100000010010101111111;
        end
        3294: begin
            cosine_reg0 <= 36'sb1010101100000010000000001001011110;
            sine_reg0   <= 36'sb100001110101100111000010111011110011;
        end
        3295: begin
            cosine_reg0 <= 36'sb1010101110111111011101110110000010;
            sine_reg0   <= 36'sb100001110110101010010110001000010111;
        end
        3296: begin
            cosine_reg0 <= 36'sb1010110001111100110100111010110101;
            sine_reg0   <= 36'sb100001110111101101111011111011000011;
        end
        3297: begin
            cosine_reg0 <= 36'sb1010110100111010000101010110000010;
            sine_reg0   <= 36'sb100001111000110001110100010011001101;
        end
        3298: begin
            cosine_reg0 <= 36'sb1010110111110111001111000101110011;
            sine_reg0   <= 36'sb100001111001110101111111010000001010;
        end
        3299: begin
            cosine_reg0 <= 36'sb1010111010110100010010001000010110;
            sine_reg0   <= 36'sb100001111010111010011100110001010001;
        end
        3300: begin
            cosine_reg0 <= 36'sb1010111101110001001110011011110011;
            sine_reg0   <= 36'sb100001111011111111001100110101110111;
        end
        3301: begin
            cosine_reg0 <= 36'sb1011000000101110000011111110011001;
            sine_reg0   <= 36'sb100001111101000100001111011101010010;
        end
        3302: begin
            cosine_reg0 <= 36'sb1011000011101010110010101110010001;
            sine_reg0   <= 36'sb100001111110001001100100100110110111;
        end
        3303: begin
            cosine_reg0 <= 36'sb1011000110100111011010101001100111;
            sine_reg0   <= 36'sb100001111111001111001100010001111100;
        end
        3304: begin
            cosine_reg0 <= 36'sb1011001001100011111011101110101000;
            sine_reg0   <= 36'sb100010000000010101000110011101110110;
        end
        3305: begin
            cosine_reg0 <= 36'sb1011001100100000010101111011011110;
            sine_reg0   <= 36'sb100010000001011011010011001001111001;
        end
        3306: begin
            cosine_reg0 <= 36'sb1011001111011100101001001110010101;
            sine_reg0   <= 36'sb100010000010100001110010010101011010;
        end
        3307: begin
            cosine_reg0 <= 36'sb1011010010011000110101100101011010;
            sine_reg0   <= 36'sb100010000011101000100011111111101110;
        end
        3308: begin
            cosine_reg0 <= 36'sb1011010101010100111010111110111001;
            sine_reg0   <= 36'sb100010000100101111101000001000001001;
        end
        3309: begin
            cosine_reg0 <= 36'sb1011011000010000111001011000111100;
            sine_reg0   <= 36'sb100010000101110110111110101110000000;
        end
        3310: begin
            cosine_reg0 <= 36'sb1011011011001100110000110001110001;
            sine_reg0   <= 36'sb100010000110111110100111110000100110;
        end
        3311: begin
            cosine_reg0 <= 36'sb1011011110001000100001000111100011;
            sine_reg0   <= 36'sb100010001000000110100011001111001110;
        end
        3312: begin
            cosine_reg0 <= 36'sb1011100001000100001010011000011111;
            sine_reg0   <= 36'sb100010001001001110110001001001001110;
        end
        3313: begin
            cosine_reg0 <= 36'sb1011100011111111101100100010110001;
            sine_reg0   <= 36'sb100010001010010111010001011101110111;
        end
        3314: begin
            cosine_reg0 <= 36'sb1011100110111011000111100100100100;
            sine_reg0   <= 36'sb100010001011100000000100001100011110;
        end
        3315: begin
            cosine_reg0 <= 36'sb1011101001110110011011011100000111;
            sine_reg0   <= 36'sb100010001100101001001001010100010110;
        end
        3316: begin
            cosine_reg0 <= 36'sb1011101100110001101000000111100100;
            sine_reg0   <= 36'sb100010001101110010100000110100110001;
        end
        3317: begin
            cosine_reg0 <= 36'sb1011101111101100101101100101001001;
            sine_reg0   <= 36'sb100010001110111100001010101101000010;
        end
        3318: begin
            cosine_reg0 <= 36'sb1011110010100111101011110011000010;
            sine_reg0   <= 36'sb100010010000000110000110111100011100;
        end
        3319: begin
            cosine_reg0 <= 36'sb1011110101100010100010101111011100;
            sine_reg0   <= 36'sb100010010001010000010101100010010000;
        end
        3320: begin
            cosine_reg0 <= 36'sb1011111000011101010010011000100011;
            sine_reg0   <= 36'sb100010010010011010110110011101110011;
        end
        3321: begin
            cosine_reg0 <= 36'sb1011111011010111111010101100100101;
            sine_reg0   <= 36'sb100010010011100101101001101110010100;
        end
        3322: begin
            cosine_reg0 <= 36'sb1011111110010010011011101001101110;
            sine_reg0   <= 36'sb100010010100110000101111010011000111;
        end
        3323: begin
            cosine_reg0 <= 36'sb1100000001001100110101001110001011;
            sine_reg0   <= 36'sb100010010101111100000111001011011101;
        end
        3324: begin
            cosine_reg0 <= 36'sb1100000100000111000111011000001001;
            sine_reg0   <= 36'sb100010010111000111110001010110100111;
        end
        3325: begin
            cosine_reg0 <= 36'sb1100000111000001010010000101110110;
            sine_reg0   <= 36'sb100010011000010011101101110011110111;
        end
        3326: begin
            cosine_reg0 <= 36'sb1100001001111011010101010101011110;
            sine_reg0   <= 36'sb100010011001011111111100100010011110;
        end
        3327: begin
            cosine_reg0 <= 36'sb1100001100110101010001000101001111;
            sine_reg0   <= 36'sb100010011010101100011101100001101101;
        end
        3328: begin
            cosine_reg0 <= 36'sb1100001111101111000101010011010101;
            sine_reg0   <= 36'sb100010011011111001010000110000110100;
        end
        3329: begin
            cosine_reg0 <= 36'sb1100010010101000110001111101111111;
            sine_reg0   <= 36'sb100010011101000110010110001111000101;
        end
        3330: begin
            cosine_reg0 <= 36'sb1100010101100010010111000011011010;
            sine_reg0   <= 36'sb100010011110010011101101111011110000;
        end
        3331: begin
            cosine_reg0 <= 36'sb1100011000011011110100100001110100;
            sine_reg0   <= 36'sb100010011111100001010111110110000100;
        end
        3332: begin
            cosine_reg0 <= 36'sb1100011011010101001010010111011001;
            sine_reg0   <= 36'sb100010100000101111010011111101010011;
        end
        3333: begin
            cosine_reg0 <= 36'sb1100011110001110011000100010010111;
            sine_reg0   <= 36'sb100010100001111101100010010000101011;
        end
        3334: begin
            cosine_reg0 <= 36'sb1100100001000111011111000000111110;
            sine_reg0   <= 36'sb100010100011001100000010101111011110;
        end
        3335: begin
            cosine_reg0 <= 36'sb1100100100000000011101110001011001;
            sine_reg0   <= 36'sb100010100100011010110101011000111010;
        end
        3336: begin
            cosine_reg0 <= 36'sb1100100110111001010100110001110111;
            sine_reg0   <= 36'sb100010100101101001111010001100001110;
        end
        3337: begin
            cosine_reg0 <= 36'sb1100101001110010000100000000100111;
            sine_reg0   <= 36'sb100010100110111001010001001000101011;
        end
        3338: begin
            cosine_reg0 <= 36'sb1100101100101010101011011011110101;
            sine_reg0   <= 36'sb100010101000001000111010001101011111;
        end
        3339: begin
            cosine_reg0 <= 36'sb1100101111100011001011000001110001;
            sine_reg0   <= 36'sb100010101001011000110101011001111000;
        end
        3340: begin
            cosine_reg0 <= 36'sb1100110010011011100010110000101000;
            sine_reg0   <= 36'sb100010101010101001000010101101000111;
        end
        3341: begin
            cosine_reg0 <= 36'sb1100110101010011110010100110101001;
            sine_reg0   <= 36'sb100010101011111001100010000110011000;
        end
        3342: begin
            cosine_reg0 <= 36'sb1100111000001011111010100010000001;
            sine_reg0   <= 36'sb100010101101001010010011100100111011;
        end
        3343: begin
            cosine_reg0 <= 36'sb1100111011000011111010100001000001;
            sine_reg0   <= 36'sb100010101110011011010111000111111101;
        end
        3344: begin
            cosine_reg0 <= 36'sb1100111101111011110010100001110101;
            sine_reg0   <= 36'sb100010101111101100101100101110101101;
        end
        3345: begin
            cosine_reg0 <= 36'sb1101000000110011100010100010101100;
            sine_reg0   <= 36'sb100010110000111110010100011000011001;
        end
        3346: begin
            cosine_reg0 <= 36'sb1101000011101011001010100001110110;
            sine_reg0   <= 36'sb100010110010010000001110000100001110;
        end
        3347: begin
            cosine_reg0 <= 36'sb1101000110100010101010011101100001;
            sine_reg0   <= 36'sb100010110011100010011001110001011001;
        end
        3348: begin
            cosine_reg0 <= 36'sb1101001001011010000010010011111011;
            sine_reg0   <= 36'sb100010110100110100110111011111001001;
        end
        3349: begin
            cosine_reg0 <= 36'sb1101001100010001010010000011010100;
            sine_reg0   <= 36'sb100010110110000111100111001100101001;
        end
        3350: begin
            cosine_reg0 <= 36'sb1101001111001000011001101001111011;
            sine_reg0   <= 36'sb100010110111011010101000111001000111;
        end
        3351: begin
            cosine_reg0 <= 36'sb1101010001111111011001000101111110;
            sine_reg0   <= 36'sb100010111000101101111100100011110001;
        end
        3352: begin
            cosine_reg0 <= 36'sb1101010100110110010000010101101101;
            sine_reg0   <= 36'sb100010111010000001100010001011110001;
        end
        3353: begin
            cosine_reg0 <= 36'sb1101010111101100111111010111010111;
            sine_reg0   <= 36'sb100010111011010101011001110000010110;
        end
        3354: begin
            cosine_reg0 <= 36'sb1101011010100011100110001001001011;
            sine_reg0   <= 36'sb100010111100101001100011010000101010;
        end
        3355: begin
            cosine_reg0 <= 36'sb1101011101011010000100101001011001;
            sine_reg0   <= 36'sb100010111101111101111110101011111011;
        end
        3356: begin
            cosine_reg0 <= 36'sb1101100000010000011010110110001111;
            sine_reg0   <= 36'sb100010111111010010101100000001010100;
        end
        3357: begin
            cosine_reg0 <= 36'sb1101100011000110101000101101111111;
            sine_reg0   <= 36'sb100011000000100111101011010000000001;
        end
        3358: begin
            cosine_reg0 <= 36'sb1101100101111100101110001110110110;
            sine_reg0   <= 36'sb100011000001111100111100010111001101;
        end
        3359: begin
            cosine_reg0 <= 36'sb1101101000110010101011010111000101;
            sine_reg0   <= 36'sb100011000011010010011111010110000100;
        end
        3360: begin
            cosine_reg0 <= 36'sb1101101011101000100000000100111100;
            sine_reg0   <= 36'sb100011000100101000010100001011110010;
        end
        3361: begin
            cosine_reg0 <= 36'sb1101101110011110001100010110101010;
            sine_reg0   <= 36'sb100011000101111110011010110111100000;
        end
        3362: begin
            cosine_reg0 <= 36'sb1101110001010011110000001010011111;
            sine_reg0   <= 36'sb100011000111010100110011011000011010;
        end
        3363: begin
            cosine_reg0 <= 36'sb1101110100001001001011011110101100;
            sine_reg0   <= 36'sb100011001000101011011101101101101100;
        end
        3364: begin
            cosine_reg0 <= 36'sb1101110110111110011110010001100000;
            sine_reg0   <= 36'sb100011001010000010011001110110011110;
        end
        3365: begin
            cosine_reg0 <= 36'sb1101111001110011101000100001001100;
            sine_reg0   <= 36'sb100011001011011001100111110001111100;
        end
        3366: begin
            cosine_reg0 <= 36'sb1101111100101000101010001100000000;
            sine_reg0   <= 36'sb100011001100110001000111011111010000;
        end
        3367: begin
            cosine_reg0 <= 36'sb1101111111011101100011010000001011;
            sine_reg0   <= 36'sb100011001110001000111000111101100100;
        end
        3368: begin
            cosine_reg0 <= 36'sb1110000010010010010011101100000000;
            sine_reg0   <= 36'sb100011001111100000111100001100000010;
        end
        3369: begin
            cosine_reg0 <= 36'sb1110000101000110111011011101101101;
            sine_reg0   <= 36'sb100011010000111001010001001001110011;
        end
        3370: begin
            cosine_reg0 <= 36'sb1110000111111011011010100011100100;
            sine_reg0   <= 36'sb100011010010010001110111110110000001;
        end
        3371: begin
            cosine_reg0 <= 36'sb1110001010101111110000111011110110;
            sine_reg0   <= 36'sb100011010011101010110000001111110101;
        end
        3372: begin
            cosine_reg0 <= 36'sb1110001101100011111110100100110010;
            sine_reg0   <= 36'sb100011010101000011111010010110011001;
        end
        3373: begin
            cosine_reg0 <= 36'sb1110010000011000000011011100101011;
            sine_reg0   <= 36'sb100011010110011101010110001000110101;
        end
        3374: begin
            cosine_reg0 <= 36'sb1110010011001011111111100001110000;
            sine_reg0   <= 36'sb100011010111110111000011100110010010;
        end
        3375: begin
            cosine_reg0 <= 36'sb1110010101111111110010110010010100;
            sine_reg0   <= 36'sb100011011001010001000010101101111010;
        end
        3376: begin
            cosine_reg0 <= 36'sb1110011000110011011101001100100110;
            sine_reg0   <= 36'sb100011011010101011010011011110110100;
        end
        3377: begin
            cosine_reg0 <= 36'sb1110011011100110111110101110111000;
            sine_reg0   <= 36'sb100011011100000101110101111000001001;
        end
        3378: begin
            cosine_reg0 <= 36'sb1110011110011010010111010111011100;
            sine_reg0   <= 36'sb100011011101100000101001111001000000;
        end
        3379: begin
            cosine_reg0 <= 36'sb1110100001001101100111000100100010;
            sine_reg0   <= 36'sb100011011110111011101111100000100011;
        end
        3380: begin
            cosine_reg0 <= 36'sb1110100100000000101101110100011101;
            sine_reg0   <= 36'sb100011100000010111000110101101111000;
        end
        3381: begin
            cosine_reg0 <= 36'sb1110100110110011101011100101011101;
            sine_reg0   <= 36'sb100011100001110010101111100000001000;
        end
        3382: begin
            cosine_reg0 <= 36'sb1110101001100110100000010101110101;
            sine_reg0   <= 36'sb100011100011001110101001110110011001;
        end
        3383: begin
            cosine_reg0 <= 36'sb1110101100011001001100000011110101;
            sine_reg0   <= 36'sb100011100100101010110101101111110100;
        end
        3384: begin
            cosine_reg0 <= 36'sb1110101111001011101110101101110000;
            sine_reg0   <= 36'sb100011100110000111010011001011011111;
        end
        3385: begin
            cosine_reg0 <= 36'sb1110110001111110001000010001111000;
            sine_reg0   <= 36'sb100011100111100100000010001000100001;
        end
        3386: begin
            cosine_reg0 <= 36'sb1110110100110000011000101110011111;
            sine_reg0   <= 36'sb100011101001000001000010100110000001;
        end
        3387: begin
            cosine_reg0 <= 36'sb1110110111100010100000000001110110;
            sine_reg0   <= 36'sb100011101010011110010100100011000110;
        end
        3388: begin
            cosine_reg0 <= 36'sb1110111010010100011110001010010000;
            sine_reg0   <= 36'sb100011101011111011110111111110110110;
        end
        3389: begin
            cosine_reg0 <= 36'sb1110111101000110010011000101111111;
            sine_reg0   <= 36'sb100011101101011001101100111000010111;
        end
        3390: begin
            cosine_reg0 <= 36'sb1110111111110111111110110011010101;
            sine_reg0   <= 36'sb100011101110110111110011001110110000;
        end
        3391: begin
            cosine_reg0 <= 36'sb1111000010101001100001010000100100;
            sine_reg0   <= 36'sb100011110000010110001011000001000111;
        end
        3392: begin
            cosine_reg0 <= 36'sb1111000101011010111010011100000000;
            sine_reg0   <= 36'sb100011110001110100110100001110100001;
        end
        3393: begin
            cosine_reg0 <= 36'sb1111001000001100001010010011111011;
            sine_reg0   <= 36'sb100011110011010011101110110110000011;
        end
        3394: begin
            cosine_reg0 <= 36'sb1111001010111101010000110110100111;
            sine_reg0   <= 36'sb100011110100110010111010110110110100;
        end
        3395: begin
            cosine_reg0 <= 36'sb1111001101101110001110000010010111;
            sine_reg0   <= 36'sb100011110110010010011000001111111001;
        end
        3396: begin
            cosine_reg0 <= 36'sb1111010000011111000001110101011111;
            sine_reg0   <= 36'sb100011110111110010000111000000010111;
        end
        3397: begin
            cosine_reg0 <= 36'sb1111010011001111101100001110010000;
            sine_reg0   <= 36'sb100011111001010010000111000111010010;
        end
        3398: begin
            cosine_reg0 <= 36'sb1111010110000000001101001010111110;
            sine_reg0   <= 36'sb100011111010110010011000100011101111;
        end
        3399: begin
            cosine_reg0 <= 36'sb1111011000110000100100101001111100;
            sine_reg0   <= 36'sb100011111100010010111011010100110100;
        end
        3400: begin
            cosine_reg0 <= 36'sb1111011011100000110010101001011101;
            sine_reg0   <= 36'sb100011111101110011101111011001100100;
        end
        3401: begin
            cosine_reg0 <= 36'sb1111011110010000110111000111110101;
            sine_reg0   <= 36'sb100011111111010100110100110001000100;
        end
        3402: begin
            cosine_reg0 <= 36'sb1111100001000000110010000011011000;
            sine_reg0   <= 36'sb100100000000110110001011011010011000;
        end
        3403: begin
            cosine_reg0 <= 36'sb1111100011110000100011011010010111;
            sine_reg0   <= 36'sb100100000010010111110011010100100100;
        end
        3404: begin
            cosine_reg0 <= 36'sb1111100110100000001011001011000111;
            sine_reg0   <= 36'sb100100000011111001101100011110101100;
        end
        3405: begin
            cosine_reg0 <= 36'sb1111101001001111101001010011111101;
            sine_reg0   <= 36'sb100100000101011011110110110111110011;
        end
        3406: begin
            cosine_reg0 <= 36'sb1111101011111110111101110011001010;
            sine_reg0   <= 36'sb100100000110111110010010011110111101;
        end
        3407: begin
            cosine_reg0 <= 36'sb1111101110101110001000100111000100;
            sine_reg0   <= 36'sb100100001000100000111111010011001100;
        end
        3408: begin
            cosine_reg0 <= 36'sb1111110001011101001001101101111111;
            sine_reg0   <= 36'sb100100001010000011111101010011100101;
        end
        3409: begin
            cosine_reg0 <= 36'sb1111110100001100000001000110001101;
            sine_reg0   <= 36'sb100100001011100111001100011111001010;
        end
        3410: begin
            cosine_reg0 <= 36'sb1111110110111010101110101110000100;
            sine_reg0   <= 36'sb100100001101001010101100110100111110;
        end
        3411: begin
            cosine_reg0 <= 36'sb1111111001101001010010100011111000;
            sine_reg0   <= 36'sb100100001110101110011110010100000011;
        end
        3412: begin
            cosine_reg0 <= 36'sb1111111100010111101100100101111100;
            sine_reg0   <= 36'sb100100010000010010100000111011011100;
        end
        3413: begin
            cosine_reg0 <= 36'sb1111111111000101111100110010100110;
            sine_reg0   <= 36'sb100100010001110110110100101010001011;
        end
        3414: begin
            cosine_reg0 <= 36'sb10000000001110100000011001000001010;
            sine_reg0   <= 36'sb100100010011011011011001011111010011;
        end
        3415: begin
            cosine_reg0 <= 36'sb10000000100100001111111100100111101;
            sine_reg0   <= 36'sb100100010101000000001111011001110101;
        end
        3416: begin
            cosine_reg0 <= 36'sb10000000111001111110010000111010011;
            sine_reg0   <= 36'sb100100010110100101010110011000110011;
        end
        3417: begin
            cosine_reg0 <= 36'sb10000001001111101011010101101100000;
            sine_reg0   <= 36'sb100100011000001010101110011011001111;
        end
        3418: begin
            cosine_reg0 <= 36'sb10000001100101010111001010101111011;
            sine_reg0   <= 36'sb100100011001110000010111100000001011;
        end
        3419: begin
            cosine_reg0 <= 36'sb10000001111011000001101111110110111;
            sine_reg0   <= 36'sb100100011011010110010001100110100110;
        end
        3420: begin
            cosine_reg0 <= 36'sb10000010010000101011000100110101011;
            sine_reg0   <= 36'sb100100011100111100011100101101100100;
        end
        3421: begin
            cosine_reg0 <= 36'sb10000010100110010011001001011101011;
            sine_reg0   <= 36'sb100100011110100010111000110100000100;
        end
        3422: begin
            cosine_reg0 <= 36'sb10000010111011111001111101100001100;
            sine_reg0   <= 36'sb100100100000001001100101111001000111;
        end
        3423: begin
            cosine_reg0 <= 36'sb10000011010001011111100000110100100;
            sine_reg0   <= 36'sb100100100001110000100011111011101110;
        end
        3424: begin
            cosine_reg0 <= 36'sb10000011100111000011110011001001000;
            sine_reg0   <= 36'sb100100100011010111110010111010111011;
        end
        3425: begin
            cosine_reg0 <= 36'sb10000011111100100110110100010001110;
            sine_reg0   <= 36'sb100100100100111111010010110101101011;
        end
        3426: begin
            cosine_reg0 <= 36'sb10000100010010001000100100000001100;
            sine_reg0   <= 36'sb100100100110100111000011101011000001;
        end
        3427: begin
            cosine_reg0 <= 36'sb10000100100111101001000010001010111;
            sine_reg0   <= 36'sb100100101000001111000101011001111100;
        end
        3428: begin
            cosine_reg0 <= 36'sb10000100111101001000001110100000101;
            sine_reg0   <= 36'sb100100101001110111011000000001011100;
        end
        3429: begin
            cosine_reg0 <= 36'sb10000101010010100110001000110101101;
            sine_reg0   <= 36'sb100100101011011111111011100000100001;
        end
        3430: begin
            cosine_reg0 <= 36'sb10000101101000000010110000111100011;
            sine_reg0   <= 36'sb100100101101001000101111110110001001;
        end
        3431: begin
            cosine_reg0 <= 36'sb10000101111101011110000110100111111;
            sine_reg0   <= 36'sb100100101110110001110101000001010101;
        end
        3432: begin
            cosine_reg0 <= 36'sb10000110010010111000001001101010111;
            sine_reg0   <= 36'sb100100110000011011001011000001000100;
        end
        3433: begin
            cosine_reg0 <= 36'sb10000110101000010000111001111000000;
            sine_reg0   <= 36'sb100100110010000100110001110100010100;
        end
        3434: begin
            cosine_reg0 <= 36'sb10000110111101101000010111000010010;
            sine_reg0   <= 36'sb100100110011101110101001011010000100;
        end
        3435: begin
            cosine_reg0 <= 36'sb10000111010010111110100000111100011;
            sine_reg0   <= 36'sb100100110101011000110001110001010100;
        end
        3436: begin
            cosine_reg0 <= 36'sb10000111101000010011010111011001010;
            sine_reg0   <= 36'sb100100110111000011001010111001000001;
        end
        3437: begin
            cosine_reg0 <= 36'sb10000111111101100110111010001011101;
            sine_reg0   <= 36'sb100100111000101101110100110000001010;
        end
        3438: begin
            cosine_reg0 <= 36'sb10001000010010111001001001000110100;
            sine_reg0   <= 36'sb100100111010011000101111010101101110;
        end
        3439: begin
            cosine_reg0 <= 36'sb10001000101000001010000011111100100;
            sine_reg0   <= 36'sb100100111100000011111010101000101010;
        end
        3440: begin
            cosine_reg0 <= 36'sb10001000111101011001101010100000110;
            sine_reg0   <= 36'sb100100111101101111010110100111111100;
        end
        3441: begin
            cosine_reg0 <= 36'sb10001001010010100111111100100110001;
            sine_reg0   <= 36'sb100100111111011011000011010010100010;
        end
        3442: begin
            cosine_reg0 <= 36'sb10001001100111110100111001111111011;
            sine_reg0   <= 36'sb100101000001000111000000100111011001;
        end
        3443: begin
            cosine_reg0 <= 36'sb10001001111101000000100010011111100;
            sine_reg0   <= 36'sb100101000010110011001110100101011111;
        end
        3444: begin
            cosine_reg0 <= 36'sb10001010010010001010110101111001100;
            sine_reg0   <= 36'sb100101000100011111101101001011110010;
        end
        3445: begin
            cosine_reg0 <= 36'sb10001010100111010011110100000000010;
            sine_reg0   <= 36'sb100101000110001100011100011001001110;
        end
        3446: begin
            cosine_reg0 <= 36'sb10001010111100011011011100100110110;
            sine_reg0   <= 36'sb100101000111111001011100001100101111;
        end
        3447: begin
            cosine_reg0 <= 36'sb10001011010001100001101111100000000;
            sine_reg0   <= 36'sb100101001001100110101100100101010100;
        end
        3448: begin
            cosine_reg0 <= 36'sb10001011100110100110101100011110111;
            sine_reg0   <= 36'sb100101001011010100001101100001111000;
        end
        3449: begin
            cosine_reg0 <= 36'sb10001011111011101010010011010110100;
            sine_reg0   <= 36'sb100101001101000001111111000001011001;
        end
        3450: begin
            cosine_reg0 <= 36'sb10001100010000101100100011111001110;
            sine_reg0   <= 36'sb100101001110110000000001000010110001;
        end
        3451: begin
            cosine_reg0 <= 36'sb10001100100101101101011101111011110;
            sine_reg0   <= 36'sb100101010000011110010011100100111110;
        end
        3452: begin
            cosine_reg0 <= 36'sb10001100111010101101000001001111100;
            sine_reg0   <= 36'sb100101010010001100110110100110111011;
        end
        3453: begin
            cosine_reg0 <= 36'sb10001101001111101011001101101000001;
            sine_reg0   <= 36'sb100101010011111011101010000111100100;
        end
        3454: begin
            cosine_reg0 <= 36'sb10001101100100101000000010111000100;
            sine_reg0   <= 36'sb100101010101101010101110000101110110;
        end
        3455: begin
            cosine_reg0 <= 36'sb10001101111001100011100000110100000;
            sine_reg0   <= 36'sb100101010111011010000010100000101010;
        end
        3456: begin
            cosine_reg0 <= 36'sb10001110001110011101100111001101011;
            sine_reg0   <= 36'sb100101011001001001100111010110111101;
        end
        3457: begin
            cosine_reg0 <= 36'sb10001110100011010110010101111000000;
            sine_reg0   <= 36'sb100101011010111001011100100111101010;
        end
        3458: begin
            cosine_reg0 <= 36'sb10001110111000001101101100100110111;
            sine_reg0   <= 36'sb100101011100101001100010010001101100;
        end
        3459: begin
            cosine_reg0 <= 36'sb10001111001101000011101011001101000;
            sine_reg0   <= 36'sb100101011110011001111000010011111101;
        end
        3460: begin
            cosine_reg0 <= 36'sb10001111100001111000010001011101111;
            sine_reg0   <= 36'sb100101100000001010011110101101011001;
        end
        3461: begin
            cosine_reg0 <= 36'sb10001111110110101011011111001100010;
            sine_reg0   <= 36'sb100101100001111011010101011100111010;
        end
        3462: begin
            cosine_reg0 <= 36'sb10010000001011011101010100001011101;
            sine_reg0   <= 36'sb100101100011101100011100100001011001;
        end
        3463: begin
            cosine_reg0 <= 36'sb10010000100000001101110000001111000;
            sine_reg0   <= 36'sb100101100101011101110011111001110011;
        end
        3464: begin
            cosine_reg0 <= 36'sb10010000110100111100110011001001100;
            sine_reg0   <= 36'sb100101100111001111011011100101000000;
        end
        3465: begin
            cosine_reg0 <= 36'sb10010001001001101010011100101110101;
            sine_reg0   <= 36'sb100101101001000001010011100001111011;
        end
        3466: begin
            cosine_reg0 <= 36'sb10010001011110010110101100110001010;
            sine_reg0   <= 36'sb100101101010110011011011101111011101;
        end
        3467: begin
            cosine_reg0 <= 36'sb10010001110011000001100011000100111;
            sine_reg0   <= 36'sb100101101100100101110100001100011111;
        end
        3468: begin
            cosine_reg0 <= 36'sb10010010000111101010111111011100110;
            sine_reg0   <= 36'sb100101101110011000011100110111111100;
        end
        3469: begin
            cosine_reg0 <= 36'sb10010010011100010011000001101011111;
            sine_reg0   <= 36'sb100101110000001011010101110000101101;
        end
        3470: begin
            cosine_reg0 <= 36'sb10010010110000111001101001100101110;
            sine_reg0   <= 36'sb100101110001111110011110110101101011;
        end
        3471: begin
            cosine_reg0 <= 36'sb10010011000101011110110110111101101;
            sine_reg0   <= 36'sb100101110011110001111000000101101110;
        end
        3472: begin
            cosine_reg0 <= 36'sb10010011011010000010101001100110111;
            sine_reg0   <= 36'sb100101110101100101100001011111101111;
        end
        3473: begin
            cosine_reg0 <= 36'sb10010011101110100101000001010100101;
            sine_reg0   <= 36'sb100101110111011001011011000010101000;
        end
        3474: begin
            cosine_reg0 <= 36'sb10010100000011000101111101111010011;
            sine_reg0   <= 36'sb100101111001001101100100101101010001;
        end
        3475: begin
            cosine_reg0 <= 36'sb10010100010111100101011111001011011;
            sine_reg0   <= 36'sb100101111011000001111110011110100001;
        end
        3476: begin
            cosine_reg0 <= 36'sb10010100101100000011100100111011000;
            sine_reg0   <= 36'sb100101111100110110101000010101010010;
        end
        3477: begin
            cosine_reg0 <= 36'sb10010101000000100000001110111100101;
            sine_reg0   <= 36'sb100101111110101011100010010000011011;
        end
        3478: begin
            cosine_reg0 <= 36'sb10010101010100111011011101000011110;
            sine_reg0   <= 36'sb100110000000100000101100001110110100;
        end
        3479: begin
            cosine_reg0 <= 36'sb10010101101001010101001111000011101;
            sine_reg0   <= 36'sb100110000010010110000110001111010110;
        end
        3480: begin
            cosine_reg0 <= 36'sb10010101111101101101100100101111110;
            sine_reg0   <= 36'sb100110000100001011110000010000110110;
        end
        3481: begin
            cosine_reg0 <= 36'sb10010110010010000100011101111011100;
            sine_reg0   <= 36'sb100110000110000001101010010010001110;
        end
        3482: begin
            cosine_reg0 <= 36'sb10010110100110011001111010011010011;
            sine_reg0   <= 36'sb100110000111110111110100010010010100;
        end
        3483: begin
            cosine_reg0 <= 36'sb10010110111010101101111001111111110;
            sine_reg0   <= 36'sb100110001001101110001110001111111111;
        end
        3484: begin
            cosine_reg0 <= 36'sb10010111001111000000011100011111010;
            sine_reg0   <= 36'sb100110001011100100111000001010000110;
        end
        3485: begin
            cosine_reg0 <= 36'sb10010111100011010001100001101100001;
            sine_reg0   <= 36'sb100110001101011011110001111111100001;
        end
        3486: begin
            cosine_reg0 <= 36'sb10010111110111100001001001011010000;
            sine_reg0   <= 36'sb100110001111010010111011101111000101;
        end
        3487: begin
            cosine_reg0 <= 36'sb10011000001011101111010011011100100;
            sine_reg0   <= 36'sb100110010001001010010101010111101001;
        end
        3488: begin
            cosine_reg0 <= 36'sb10011000011111111011111111100111000;
            sine_reg0   <= 36'sb100110010011000001111110111000000100;
        end
        3489: begin
            cosine_reg0 <= 36'sb10011000110100000111001101101101000;
            sine_reg0   <= 36'sb100110010100111001111000001111001100;
        end
        3490: begin
            cosine_reg0 <= 36'sb10011001001000010000111101100010010;
            sine_reg0   <= 36'sb100110010110110010000001011011110110;
        end
        3491: begin
            cosine_reg0 <= 36'sb10011001011100011001001110111010001;
            sine_reg0   <= 36'sb100110011000101010011010011100111001;
        end
        3492: begin
            cosine_reg0 <= 36'sb10011001110000100000000001101000011;
            sine_reg0   <= 36'sb100110011010100011000011010001001011;
        end
        3493: begin
            cosine_reg0 <= 36'sb10011010000100100101010101100000011;
            sine_reg0   <= 36'sb100110011100011011111011110111100000;
        end
        3494: begin
            cosine_reg0 <= 36'sb10011010011000101001001010010110000;
            sine_reg0   <= 36'sb100110011110010101000100001110101111;
        end
        3495: begin
            cosine_reg0 <= 36'sb10011010101100101011011111111100101;
            sine_reg0   <= 36'sb100110100000001110011100010101101101;
        end
        3496: begin
            cosine_reg0 <= 36'sb10011011000000101100010110001000001;
            sine_reg0   <= 36'sb100110100010001000000100001011001111;
        end
        3497: begin
            cosine_reg0 <= 36'sb10011011010100101011101100101100000;
            sine_reg0   <= 36'sb100110100100000001111011101110001001;
        end
        3498: begin
            cosine_reg0 <= 36'sb10011011101000101001100011011100000;
            sine_reg0   <= 36'sb100110100101111100000010111101010001;
        end
        3499: begin
            cosine_reg0 <= 36'sb10011011111100100101111010001011110;
            sine_reg0   <= 36'sb100110100111110110011001110111011100;
        end
        3500: begin
            cosine_reg0 <= 36'sb10011100010000100000110000101110111;
            sine_reg0   <= 36'sb100110101001110001000000011011011101;
        end
        3501: begin
            cosine_reg0 <= 36'sb10011100100100011010000110111001011;
            sine_reg0   <= 36'sb100110101011101011110110101000001010;
        end
        3502: begin
            cosine_reg0 <= 36'sb10011100111000010001111100011110101;
            sine_reg0   <= 36'sb100110101101100110111100011100010110;
        end
        3503: begin
            cosine_reg0 <= 36'sb10011101001100001000010001010010101;
            sine_reg0   <= 36'sb100110101111100010010001110110110101;
        end
        3504: begin
            cosine_reg0 <= 36'sb10011101011111111101000101001000111;
            sine_reg0   <= 36'sb100110110001011101110110110110011100;
        end
        3505: begin
            cosine_reg0 <= 36'sb10011101110011110000010111110101100;
            sine_reg0   <= 36'sb100110110011011001101011011001111110;
        end
        3506: begin
            cosine_reg0 <= 36'sb10011110000111100010001001001100000;
            sine_reg0   <= 36'sb100110110101010101101111100000001111;
        end
        3507: begin
            cosine_reg0 <= 36'sb10011110011011010010011001000000010;
            sine_reg0   <= 36'sb100110110111010010000011001000000011;
        end
        3508: begin
            cosine_reg0 <= 36'sb10011110101111000001000111000110001;
            sine_reg0   <= 36'sb100110111001001110100110010000001100;
        end
        3509: begin
            cosine_reg0 <= 36'sb10011111000010101110010011010001011;
            sine_reg0   <= 36'sb100110111011001011011000110111011101;
        end
        3510: begin
            cosine_reg0 <= 36'sb10011111010110011001111101010101111;
            sine_reg0   <= 36'sb100110111101001000011010111100101011;
        end
        3511: begin
            cosine_reg0 <= 36'sb10011111101010000100000101000111100;
            sine_reg0   <= 36'sb100110111111000101101100011110100111;
        end
        3512: begin
            cosine_reg0 <= 36'sb10011111111101101100101010011010001;
            sine_reg0   <= 36'sb100111000001000011001101011100000101;
        end
        3513: begin
            cosine_reg0 <= 36'sb10100000010001010011101101000001101;
            sine_reg0   <= 36'sb100111000011000000111101110011110111;
        end
        3514: begin
            cosine_reg0 <= 36'sb10100000100100111001001100110001111;
            sine_reg0   <= 36'sb100111000100111110111101100100101111;
        end
        3515: begin
            cosine_reg0 <= 36'sb10100000111000011101001001011110110;
            sine_reg0   <= 36'sb100111000110111101001100101101011111;
        end
        3516: begin
            cosine_reg0 <= 36'sb10100001001011111111100010111100011;
            sine_reg0   <= 36'sb100111001000111011101011001100111011;
        end
        3517: begin
            cosine_reg0 <= 36'sb10100001011111100000011000111110100;
            sine_reg0   <= 36'sb100111001010111010011001000001110100;
        end
        3518: begin
            cosine_reg0 <= 36'sb10100001110010111111101011011001010;
            sine_reg0   <= 36'sb100111001100111001010110001010111011;
        end
        3519: begin
            cosine_reg0 <= 36'sb10100010000110011101011010000000100;
            sine_reg0   <= 36'sb100111001110111000100010100111000010;
        end
        3520: begin
            cosine_reg0 <= 36'sb10100010011001111001100100101000010;
            sine_reg0   <= 36'sb100111010000110111111110010100111100;
        end
        3521: begin
            cosine_reg0 <= 36'sb10100010101101010100001011000100100;
            sine_reg0   <= 36'sb100111010010110111101001010011011000;
        end
        3522: begin
            cosine_reg0 <= 36'sb10100011000000101101001101001001010;
            sine_reg0   <= 36'sb100111010100110111100011100001001001;
        end
        3523: begin
            cosine_reg0 <= 36'sb10100011010100000100101010101010101;
            sine_reg0   <= 36'sb100111010110110111101100111101000000;
        end
        3524: begin
            cosine_reg0 <= 36'sb10100011100111011010100011011100101;
            sine_reg0   <= 36'sb100111011000111000000101100101101101;
        end
        3525: begin
            cosine_reg0 <= 36'sb10100011111010101110110111010011011;
            sine_reg0   <= 36'sb100111011010111000101101011010000010;
        end
        3526: begin
            cosine_reg0 <= 36'sb10100100001110000001100110000011000;
            sine_reg0   <= 36'sb100111011100111001100100011000101111;
        end
        3527: begin
            cosine_reg0 <= 36'sb10100100100001010010101111011111011;
            sine_reg0   <= 36'sb100111011110111010101010100000100100;
        end
        3528: begin
            cosine_reg0 <= 36'sb10100100110100100010010011011100110;
            sine_reg0   <= 36'sb100111100000111011111111110000010010;
        end
        3529: begin
            cosine_reg0 <= 36'sb10100101000111110000010001101111011;
            sine_reg0   <= 36'sb100111100010111101100100000110101010;
        end
        3530: begin
            cosine_reg0 <= 36'sb10100101011010111100101010001011001;
            sine_reg0   <= 36'sb100111100100111111010111100010011010;
        end
        3531: begin
            cosine_reg0 <= 36'sb10100101101110000111011100100100011;
            sine_reg0   <= 36'sb100111100111000001011010000010010100;
        end
        3532: begin
            cosine_reg0 <= 36'sb10100110000001010000101000101111010;
            sine_reg0   <= 36'sb100111101001000011101011100101000110;
        end
        3533: begin
            cosine_reg0 <= 36'sb10100110010100011000001110100000000;
            sine_reg0   <= 36'sb100111101011000110001100001001100010;
        end
        3534: begin
            cosine_reg0 <= 36'sb10100110100111011110001101101010110;
            sine_reg0   <= 36'sb100111101101001000111011101110010101;
        end
        3535: begin
            cosine_reg0 <= 36'sb10100110111010100010100110000011101;
            sine_reg0   <= 36'sb100111101111001011111010010010010000;
        end
        3536: begin
            cosine_reg0 <= 36'sb10100111001101100101010111011111000;
            sine_reg0   <= 36'sb100111110001001111000111110100000001;
        end
        3537: begin
            cosine_reg0 <= 36'sb10100111100000100110100001110001001;
            sine_reg0   <= 36'sb100111110011010010100100010010011000;
        end
        3538: begin
            cosine_reg0 <= 36'sb10100111110011100110000100101110011;
            sine_reg0   <= 36'sb100111110101010110001111101100000011;
        end
        3539: begin
            cosine_reg0 <= 36'sb10101000000110100100000000001010110;
            sine_reg0   <= 36'sb100111110111011010001001111111110010;
        end
        3540: begin
            cosine_reg0 <= 36'sb10101000011001100000010011111010110;
            sine_reg0   <= 36'sb100111111001011110010011001100010011;
        end
        3541: begin
            cosine_reg0 <= 36'sb10101000101100011010111111110010101;
            sine_reg0   <= 36'sb100111111011100010101011010000010101;
        end
        3542: begin
            cosine_reg0 <= 36'sb10101000111111010100000011100110110;
            sine_reg0   <= 36'sb100111111101100111010010001010100101;
        end
        3543: begin
            cosine_reg0 <= 36'sb10101001010010001011011111001011011;
            sine_reg0   <= 36'sb100111111111101100000111111001110011;
        end
        3544: begin
            cosine_reg0 <= 36'sb10101001100101000001010010010101000;
            sine_reg0   <= 36'sb101000000001110001001100011100101011;
        end
        3545: begin
            cosine_reg0 <= 36'sb10101001110111110101011100111000000;
            sine_reg0   <= 36'sb101000000011110110011111110001111100;
        end
        3546: begin
            cosine_reg0 <= 36'sb10101010001010100111111110101000101;
            sine_reg0   <= 36'sb101000000101111100000001111000010101;
        end
        3547: begin
            cosine_reg0 <= 36'sb10101010011101011000110111011011011;
            sine_reg0   <= 36'sb101000001000000001110010101110100001;
        end
        3548: begin
            cosine_reg0 <= 36'sb10101010110000001000000111000100101;
            sine_reg0   <= 36'sb101000001010000111110010010011010000;
        end
        3549: begin
            cosine_reg0 <= 36'sb10101011000010110101101101011000111;
            sine_reg0   <= 36'sb101000001100001110000000100101001110;
        end
        3550: begin
            cosine_reg0 <= 36'sb10101011010101100001101010001100101;
            sine_reg0   <= 36'sb101000001110010100011101100011001000;
        end
        3551: begin
            cosine_reg0 <= 36'sb10101011101000001011111101010100010;
            sine_reg0   <= 36'sb101000010000011011001001001011101100;
        end
        3552: begin
            cosine_reg0 <= 36'sb10101011111010110100100110100100011;
            sine_reg0   <= 36'sb101000010010100010000011011101100110;
        end
        3553: begin
            cosine_reg0 <= 36'sb10101100001101011011100101110001010;
            sine_reg0   <= 36'sb101000010100101001001100010111100100;
        end
        3554: begin
            cosine_reg0 <= 36'sb10101100100000000000111010101111101;
            sine_reg0   <= 36'sb101000010110110000100011111000010001;
        end
        3555: begin
            cosine_reg0 <= 36'sb10101100110010100100100101010100000;
            sine_reg0   <= 36'sb101000011000111000001001111110011011;
        end
        3556: begin
            cosine_reg0 <= 36'sb10101101000101000110100101010010111;
            sine_reg0   <= 36'sb101000011010111111111110101000101101;
        end
        3557: begin
            cosine_reg0 <= 36'sb10101101010111100110111010100000110;
            sine_reg0   <= 36'sb101000011101001000000001110101110100;
        end
        3558: begin
            cosine_reg0 <= 36'sb10101101101010000101100100110010011;
            sine_reg0   <= 36'sb101000011111010000010011100100011101;
        end
        3559: begin
            cosine_reg0 <= 36'sb10101101111100100010100011111100010;
            sine_reg0   <= 36'sb101000100001011000110011110011010010;
        end
        3560: begin
            cosine_reg0 <= 36'sb10101110001110111101110111110011001;
            sine_reg0   <= 36'sb101000100011100001100010100001000000;
        end
        3561: begin
            cosine_reg0 <= 36'sb10101110100001010111100000001011011;
            sine_reg0   <= 36'sb101000100101101010011111101100010010;
        end
        3562: begin
            cosine_reg0 <= 36'sb10101110110011101111011100111001111;
            sine_reg0   <= 36'sb101000100111110011101011010011110101;
        end
        3563: begin
            cosine_reg0 <= 36'sb10101111000110000101101101110011001;
            sine_reg0   <= 36'sb101000101001111101000101010110010010;
        end
        3564: begin
            cosine_reg0 <= 36'sb10101111011000011010010010101100000;
            sine_reg0   <= 36'sb101000101100000110101101110010010111;
        end
        3565: begin
            cosine_reg0 <= 36'sb10101111101010101101001011011001001;
            sine_reg0   <= 36'sb101000101110010000100100100110101100;
        end
        3566: begin
            cosine_reg0 <= 36'sb10101111111100111110010111101111001;
            sine_reg0   <= 36'sb101000110000011010101001110001111111;
        end
        3567: begin
            cosine_reg0 <= 36'sb10110000001111001101110111100010110;
            sine_reg0   <= 36'sb101000110010100100111101010010111001;
        end
        3568: begin
            cosine_reg0 <= 36'sb10110000100001011011101010101000111;
            sine_reg0   <= 36'sb101000110100101111011111001000000101;
        end
        3569: begin
            cosine_reg0 <= 36'sb10110000110011100111110000110110001;
            sine_reg0   <= 36'sb101000110110111010001111010000001101;
        end
        3570: begin
            cosine_reg0 <= 36'sb10110001000101110010001001111111010;
            sine_reg0   <= 36'sb101000111001000101001101101001111101;
        end
        3571: begin
            cosine_reg0 <= 36'sb10110001010111111010110101111001010;
            sine_reg0   <= 36'sb101000111011010000011010010011111110;
        end
        3572: begin
            cosine_reg0 <= 36'sb10110001101010000001110100011000110;
            sine_reg0   <= 36'sb101000111101011011110101001100111011;
        end
        3573: begin
            cosine_reg0 <= 36'sb10110001111100000111000101010010110;
            sine_reg0   <= 36'sb101000111111100111011110010011011101;
        end
        3574: begin
            cosine_reg0 <= 36'sb10110010001110001010101000011011111;
            sine_reg0   <= 36'sb101001000001110011010101100110001110;
        end
        3575: begin
            cosine_reg0 <= 36'sb10110010100000001100011101101001001;
            sine_reg0   <= 36'sb101001000011111111011011000011111001;
        end
        3576: begin
            cosine_reg0 <= 36'sb10110010110010001100100100101111011;
            sine_reg0   <= 36'sb101001000110001011101110101011000110;
        end
        3577: begin
            cosine_reg0 <= 36'sb10110011000100001010111101100011101;
            sine_reg0   <= 36'sb101001001000011000010000011010011111;
        end
        3578: begin
            cosine_reg0 <= 36'sb10110011010110000111100111111010100;
            sine_reg0   <= 36'sb101001001010100101000000010000101110;
        end
        3579: begin
            cosine_reg0 <= 36'sb10110011101000000010100011101001001;
            sine_reg0   <= 36'sb101001001100110001111110001100011011;
        end
        3580: begin
            cosine_reg0 <= 36'sb10110011111001111011110000100100100;
            sine_reg0   <= 36'sb101001001110111111001010001100010000;
        end
        3581: begin
            cosine_reg0 <= 36'sb10110100001011110011001110100001011;
            sine_reg0   <= 36'sb101001010001001100100100001110110110;
        end
        3582: begin
            cosine_reg0 <= 36'sb10110100011101101000111101010101000;
            sine_reg0   <= 36'sb101001010011011010001100010010110101;
        end
        3583: begin
            cosine_reg0 <= 36'sb10110100101111011100111100110100001;
            sine_reg0   <= 36'sb101001010101101000000010010110110110;
        end
        3584: begin
            cosine_reg0 <= 36'sb10110101000001001111001100110011111;
            sine_reg0   <= 36'sb101001010111110110000110011001100001;
        end
        3585: begin
            cosine_reg0 <= 36'sb10110101010010111111101101001001010;
            sine_reg0   <= 36'sb101001011010000100011000011001011111;
        end
        3586: begin
            cosine_reg0 <= 36'sb10110101100100101110011101101001011;
            sine_reg0   <= 36'sb101001011100010010111000010101011000;
        end
        3587: begin
            cosine_reg0 <= 36'sb10110101110110011011011110001001010;
            sine_reg0   <= 36'sb101001011110100001100110001011110101;
        end
        3588: begin
            cosine_reg0 <= 36'sb10110110001000000110101110011110000;
            sine_reg0   <= 36'sb101001100000110000100001111011011100;
        end
        3589: begin
            cosine_reg0 <= 36'sb10110110011001110000001110011100101;
            sine_reg0   <= 36'sb101001100010111111101011100010110111;
        end
        3590: begin
            cosine_reg0 <= 36'sb10110110101011010111111101111010010;
            sine_reg0   <= 36'sb101001100101001111000011000000101100;
        end
        3591: begin
            cosine_reg0 <= 36'sb10110110111100111101111100101100001;
            sine_reg0   <= 36'sb101001100111011110101000010011100011;
        end
        3592: begin
            cosine_reg0 <= 36'sb10110111001110100010001010100111010;
            sine_reg0   <= 36'sb101001101001101110011011011010000101;
        end
        3593: begin
            cosine_reg0 <= 36'sb10110111100000000100100111100000111;
            sine_reg0   <= 36'sb101001101011111110011100010010110111;
        end
        3594: begin
            cosine_reg0 <= 36'sb10110111110001100101010011001110010;
            sine_reg0   <= 36'sb101001101110001110101010111100100001;
        end
        3595: begin
            cosine_reg0 <= 36'sb10111000000011000100001101100100011;
            sine_reg0   <= 36'sb101001110000011111000111010101101010;
        end
        3596: begin
            cosine_reg0 <= 36'sb10111000010100100001010110011000101;
            sine_reg0   <= 36'sb101001110010101111110001011100111010;
        end
        3597: begin
            cosine_reg0 <= 36'sb10111000100101111100101101100000010;
            sine_reg0   <= 36'sb101001110101000000101001010000110110;
        end
        3598: begin
            cosine_reg0 <= 36'sb10111000110111010110010010110000011;
            sine_reg0   <= 36'sb101001110111010001101110110000000110;
        end
        3599: begin
            cosine_reg0 <= 36'sb10111001001000101110000101111110011;
            sine_reg0   <= 36'sb101001111001100011000001111001001111;
        end
        3600: begin
            cosine_reg0 <= 36'sb10111001011010000100000110111111011;
            sine_reg0   <= 36'sb101001111011110100100010101010111001;
        end
        3601: begin
            cosine_reg0 <= 36'sb10111001101011011000010101101000111;
            sine_reg0   <= 36'sb101001111110000110010001000011101010;
        end
        3602: begin
            cosine_reg0 <= 36'sb10111001111100101010110001110000001;
            sine_reg0   <= 36'sb101010000000011000001101000010000111;
        end
        3603: begin
            cosine_reg0 <= 36'sb10111010001101111011011011001010100;
            sine_reg0   <= 36'sb101010000010101010010110100100110111;
        end
        3604: begin
            cosine_reg0 <= 36'sb10111010011111001010010001101101001;
            sine_reg0   <= 36'sb101010000100111100101101101010100000;
        end
        3605: begin
            cosine_reg0 <= 36'sb10111010110000010111010101001101110;
            sine_reg0   <= 36'sb101010000111001111010010010001100111;
        end
        3606: begin
            cosine_reg0 <= 36'sb10111011000001100010100101100001011;
            sine_reg0   <= 36'sb101010001001100010000100011000110001;
        end
        3607: begin
            cosine_reg0 <= 36'sb10111011010010101100000010011101110;
            sine_reg0   <= 36'sb101010001011110101000011111110100101;
        end
        3608: begin
            cosine_reg0 <= 36'sb10111011100011110011101011111000000;
            sine_reg0   <= 36'sb101010001110001000010001000001100111;
        end
        3609: begin
            cosine_reg0 <= 36'sb10111011110100111001100001100101110;
            sine_reg0   <= 36'sb101010010000011011101011100000011110;
        end
        3610: begin
            cosine_reg0 <= 36'sb10111100000101111101100011011100011;
            sine_reg0   <= 36'sb101010010010101111010011011001101101;
        end
        3611: begin
            cosine_reg0 <= 36'sb10111100010110111111110001010001100;
            sine_reg0   <= 36'sb101010010101000011001000101011111010;
        end
        3612: begin
            cosine_reg0 <= 36'sb10111100101000000000001010111010011;
            sine_reg0   <= 36'sb101010010111010111001011010101101001;
        end
        3613: begin
            cosine_reg0 <= 36'sb10111100111000111110110000001100101;
            sine_reg0   <= 36'sb101010011001101011011011010101100000;
        end
        3614: begin
            cosine_reg0 <= 36'sb10111101001001111011100000111101111;
            sine_reg0   <= 36'sb101010011011111111111000101010000011;
        end
        3615: begin
            cosine_reg0 <= 36'sb10111101011010110110011101000011100;
            sine_reg0   <= 36'sb101010011110010100100011010001110110;
        end
        3616: begin
            cosine_reg0 <= 36'sb10111101101011101111100100010011010;
            sine_reg0   <= 36'sb101010100000101001011011001011011101;
        end
        3617: begin
            cosine_reg0 <= 36'sb10111101111100100110110110100010100;
            sine_reg0   <= 36'sb101010100010111110100000010101011110;
        end
        3618: begin
            cosine_reg0 <= 36'sb10111110001101011100010011100111000;
            sine_reg0   <= 36'sb101010100101010011110010101110011011;
        end
        3619: begin
            cosine_reg0 <= 36'sb10111110011110001111111011010110010;
            sine_reg0   <= 36'sb101010100111101001010010010100111001;
        end
        3620: begin
            cosine_reg0 <= 36'sb10111110101111000001101101100110000;
            sine_reg0   <= 36'sb101010101001111110111111000111011011;
        end
        3621: begin
            cosine_reg0 <= 36'sb10111110111111110001101010001011111;
            sine_reg0   <= 36'sb101010101100010100111001000100100101;
        end
        3622: begin
            cosine_reg0 <= 36'sb10111111010000011111110000111101011;
            sine_reg0   <= 36'sb101010101110101011000000001010111011;
        end
        3623: begin
            cosine_reg0 <= 36'sb10111111100001001100000001110000100;
            sine_reg0   <= 36'sb101010110001000001010100011001000000;
        end
        3624: begin
            cosine_reg0 <= 36'sb10111111110001110110011100011010101;
            sine_reg0   <= 36'sb101010110011010111110101101101011000;
        end
        3625: begin
            cosine_reg0 <= 36'sb11000000000010011111000000110001101;
            sine_reg0   <= 36'sb101010110101101110100100000110100101;
        end
        3626: begin
            cosine_reg0 <= 36'sb11000000010011000101101110101011011;
            sine_reg0   <= 36'sb101010111000000101011111100011001010;
        end
        3627: begin
            cosine_reg0 <= 36'sb11000000100011101010100101111101011;
            sine_reg0   <= 36'sb101010111010011100101000000001101011;
        end
        3628: begin
            cosine_reg0 <= 36'sb11000000110100001101100110011101101;
            sine_reg0   <= 36'sb101010111100110011111101100000101010;
        end
        3629: begin
            cosine_reg0 <= 36'sb11000001000100101110110000000001110;
            sine_reg0   <= 36'sb101010111111001011011111111110101010;
        end
        3630: begin
            cosine_reg0 <= 36'sb11000001010101001110000010011111101;
            sine_reg0   <= 36'sb101011000001100011001111011010001101;
        end
        3631: begin
            cosine_reg0 <= 36'sb11000001100101101011011101101101000;
            sine_reg0   <= 36'sb101011000011111011001011110001110111;
        end
        3632: begin
            cosine_reg0 <= 36'sb11000001110110000111000001011111111;
            sine_reg0   <= 36'sb101011000110010011010101000100001000;
        end
        3633: begin
            cosine_reg0 <= 36'sb11000010000110100000101101101110000;
            sine_reg0   <= 36'sb101011001000101011101011001111100011;
        end
        3634: begin
            cosine_reg0 <= 36'sb11000010010110111000100010001101011;
            sine_reg0   <= 36'sb101011001011000100001110010010101010;
        end
        3635: begin
            cosine_reg0 <= 36'sb11000010100111001110011110110011110;
            sine_reg0   <= 36'sb101011001101011100111110001100000000;
        end
        3636: begin
            cosine_reg0 <= 36'sb11000010110111100010100011010111010;
            sine_reg0   <= 36'sb101011001111110101111010111010000110;
        end
        3637: begin
            cosine_reg0 <= 36'sb11000011000111110100101111101101100;
            sine_reg0   <= 36'sb101011010010001111000100011011011101;
        end
        3638: begin
            cosine_reg0 <= 36'sb11000011011000000101000011101100110;
            sine_reg0   <= 36'sb101011010100101000011010101110100111;
        end
        3639: begin
            cosine_reg0 <= 36'sb11000011101000010011011111001010110;
            sine_reg0   <= 36'sb101011010111000001111101110010000101;
        end
        3640: begin
            cosine_reg0 <= 36'sb11000011111000100000000001111101110;
            sine_reg0   <= 36'sb101011011001011011101101100100011010;
        end
        3641: begin
            cosine_reg0 <= 36'sb11000100001000101010101011111011100;
            sine_reg0   <= 36'sb101011011011110101101010000100000101;
        end
        3642: begin
            cosine_reg0 <= 36'sb11000100011000110011011100111010001;
            sine_reg0   <= 36'sb101011011110001111110011001111101000;
        end
        3643: begin
            cosine_reg0 <= 36'sb11000100101000111010010100101111110;
            sine_reg0   <= 36'sb101011100000101010001001000101100101;
        end
        3644: begin
            cosine_reg0 <= 36'sb11000100111000111111010011010010011;
            sine_reg0   <= 36'sb101011100011000100101011100100011011;
        end
        3645: begin
            cosine_reg0 <= 36'sb11000101001001000010011000011000000;
            sine_reg0   <= 36'sb101011100101011111011010101010101011;
        end
        3646: begin
            cosine_reg0 <= 36'sb11000101011001000011100011110110111;
            sine_reg0   <= 36'sb101011100111111010010110010110110110;
        end
        3647: begin
            cosine_reg0 <= 36'sb11000101101001000010110101100101000;
            sine_reg0   <= 36'sb101011101010010101011110100111011100;
        end
        3648: begin
            cosine_reg0 <= 36'sb11000101111001000000001101011000100;
            sine_reg0   <= 36'sb101011101100110000110011011010111110;
        end
        3649: begin
            cosine_reg0 <= 36'sb11000110001000111011101011000111110;
            sine_reg0   <= 36'sb101011101111001100010100101111111100;
        end
        3650: begin
            cosine_reg0 <= 36'sb11000110011000110101001110101000101;
            sine_reg0   <= 36'sb101011110001101000000010100100110110;
        end
        3651: begin
            cosine_reg0 <= 36'sb11000110101000101100110111110001100;
            sine_reg0   <= 36'sb101011110100000011111100111000001100;
        end
        3652: begin
            cosine_reg0 <= 36'sb11000110111000100010100110011000101;
            sine_reg0   <= 36'sb101011110110100000000011101000011101;
        end
        3653: begin
            cosine_reg0 <= 36'sb11000111001000010110011010010100001;
            sine_reg0   <= 36'sb101011111000111100010110110100001010;
        end
        3654: begin
            cosine_reg0 <= 36'sb11000111011000001000010011011010001;
            sine_reg0   <= 36'sb101011111011011000110110011001110001;
        end
        3655: begin
            cosine_reg0 <= 36'sb11000111100111111000010001100001001;
            sine_reg0   <= 36'sb101011111101110101100010010111110011;
        end
        3656: begin
            cosine_reg0 <= 36'sb11000111110111100110010100011111011;
            sine_reg0   <= 36'sb101100000000010010011010101100101111;
        end
        3657: begin
            cosine_reg0 <= 36'sb11001000000111010010011100001011001;
            sine_reg0   <= 36'sb101100000010101111011111010111000100;
        end
        3658: begin
            cosine_reg0 <= 36'sb11001000010110111100101000011010101;
            sine_reg0   <= 36'sb101100000101001100110000010101010001;
        end
        3659: begin
            cosine_reg0 <= 36'sb11001000100110100100111001000100011;
            sine_reg0   <= 36'sb101100000111101010001101100101110101;
        end
        3660: begin
            cosine_reg0 <= 36'sb11001000110110001011001101111110100;
            sine_reg0   <= 36'sb101100001010000111110111000111001111;
        end
        3661: begin
            cosine_reg0 <= 36'sb11001001000101101111100110111111101;
            sine_reg0   <= 36'sb101100001100100101101100110111111110;
        end
        3662: begin
            cosine_reg0 <= 36'sb11001001010101010010000011111110001;
            sine_reg0   <= 36'sb101100001111000011101110110110100000;
        end
        3663: begin
            cosine_reg0 <= 36'sb11001001100100110010100100110000010;
            sine_reg0   <= 36'sb101100010001100001111101000001010100;
        end
        3664: begin
            cosine_reg0 <= 36'sb11001001110100010001001001001100100;
            sine_reg0   <= 36'sb101100010100000000010111010110111001;
        end
        3665: begin
            cosine_reg0 <= 36'sb11001010000011101101110001001001011;
            sine_reg0   <= 36'sb101100010110011110111101110101101011;
        end
        3666: begin
            cosine_reg0 <= 36'sb11001010010011001000011100011101010;
            sine_reg0   <= 36'sb101100011000111101110000011100001011;
        end
        3667: begin
            cosine_reg0 <= 36'sb11001010100010100001001010111110110;
            sine_reg0   <= 36'sb101100011011011100101111001000110101;
        end
        3668: begin
            cosine_reg0 <= 36'sb11001010110001110111111100100100011;
            sine_reg0   <= 36'sb101100011101111011111001111010001001;
        end
        3669: begin
            cosine_reg0 <= 36'sb11001011000001001100110001000100100;
            sine_reg0   <= 36'sb101100100000011011010000101110100010;
        end
        3670: begin
            cosine_reg0 <= 36'sb11001011010000011111101000010101111;
            sine_reg0   <= 36'sb101100100010111010110011100100100000;
        end
        3671: begin
            cosine_reg0 <= 36'sb11001011011111110000100010001110111;
            sine_reg0   <= 36'sb101100100101011010100010011010100000;
        end
        3672: begin
            cosine_reg0 <= 36'sb11001011101110111111011110100110001;
            sine_reg0   <= 36'sb101100100111111010011101001110111111;
        end
        3673: begin
            cosine_reg0 <= 36'sb11001011111110001100011101010010011;
            sine_reg0   <= 36'sb101100101010011010100100000000011011;
        end
        3674: begin
            cosine_reg0 <= 36'sb11001100001101010111011110001010001;
            sine_reg0   <= 36'sb101100101100111010110110101101010000;
        end
        3675: begin
            cosine_reg0 <= 36'sb11001100011100100000100001000100000;
            sine_reg0   <= 36'sb101100101111011011010101010011111101;
        end
        3676: begin
            cosine_reg0 <= 36'sb11001100101011100111100101110110101;
            sine_reg0   <= 36'sb101100110001111011111111110010111101;
        end
        3677: begin
            cosine_reg0 <= 36'sb11001100111010101100101100011000111;
            sine_reg0   <= 36'sb101100110100011100110110001000101111;
        end
        3678: begin
            cosine_reg0 <= 36'sb11001101001001101111110100100001010;
            sine_reg0   <= 36'sb101100110110111101111000010011101110;
        end
        3679: begin
            cosine_reg0 <= 36'sb11001101011000110000111110000110100;
            sine_reg0   <= 36'sb101100111001011111000110010010011000;
        end
        3680: begin
            cosine_reg0 <= 36'sb11001101100111110000001000111111100;
            sine_reg0   <= 36'sb101100111100000000100000000011001000;
        end
        3681: begin
            cosine_reg0 <= 36'sb11001101110110101101010101000010111;
            sine_reg0   <= 36'sb101100111110100010000101100100011100;
        end
        3682: begin
            cosine_reg0 <= 36'sb11001110000101101000100010000111011;
            sine_reg0   <= 36'sb101101000001000011110110110100110000;
        end
        3683: begin
            cosine_reg0 <= 36'sb11001110010100100001110000000011111;
            sine_reg0   <= 36'sb101101000011100101110011110010011111;
        end
        3684: begin
            cosine_reg0 <= 36'sb11001110100011011000111110101111010;
            sine_reg0   <= 36'sb101101000110000111111100011100000110;
        end
        3685: begin
            cosine_reg0 <= 36'sb11001110110010001110001110000000001;
            sine_reg0   <= 36'sb101101001000101010010000110000000010;
        end
        3686: begin
            cosine_reg0 <= 36'sb11001111000001000001011101101101100;
            sine_reg0   <= 36'sb101101001011001100110000101100101101;
        end
        3687: begin
            cosine_reg0 <= 36'sb11001111001111110010101101101110010;
            sine_reg0   <= 36'sb101101001101101111011100010000100100;
        end
        3688: begin
            cosine_reg0 <= 36'sb11001111011110100001111101111001010;
            sine_reg0   <= 36'sb101101010000010010010011011010000010;
        end
        3689: begin
            cosine_reg0 <= 36'sb11001111101101001111001110000101010;
            sine_reg0   <= 36'sb101101010010110101010110000111100011;
        end
        3690: begin
            cosine_reg0 <= 36'sb11001111111011111010011110001001100;
            sine_reg0   <= 36'sb101101010101011000100100010111100010;
        end
        3691: begin
            cosine_reg0 <= 36'sb11010000001010100011101101111100101;
            sine_reg0   <= 36'sb101101010111111011111110001000011011;
        end
        3692: begin
            cosine_reg0 <= 36'sb11010000011001001010111101010101110;
            sine_reg0   <= 36'sb101101011010011111100011011000101000;
        end
        3693: begin
            cosine_reg0 <= 36'sb11010000100111110000001100001011111;
            sine_reg0   <= 36'sb101101011101000011010100000110100101;
        end
        3694: begin
            cosine_reg0 <= 36'sb11010000110110010011011010010101111;
            sine_reg0   <= 36'sb101101011111100111010000010000101101;
        end
        3695: begin
            cosine_reg0 <= 36'sb11010001000100110100100111101011000;
            sine_reg0   <= 36'sb101101100010001011010111110101011011;
        end
        3696: begin
            cosine_reg0 <= 36'sb11010001010011010011110100000010001;
            sine_reg0   <= 36'sb101101100100101111101010110011001001;
        end
        3697: begin
            cosine_reg0 <= 36'sb11010001100001110000111111010010010;
            sine_reg0   <= 36'sb101101100111010100001001001000010011;
        end
        3698: begin
            cosine_reg0 <= 36'sb11010001110000001100001001010010101;
            sine_reg0   <= 36'sb101101101001111000110010110011010010;
        end
        3699: begin
            cosine_reg0 <= 36'sb11010001111110100101010001111010011;
            sine_reg0   <= 36'sb101101101100011101100111110010100001;
        end
        3700: begin
            cosine_reg0 <= 36'sb11010010001100111100011001000000100;
            sine_reg0   <= 36'sb101101101111000010101000000100011010;
        end
        3701: begin
            cosine_reg0 <= 36'sb11010010011011010001011110011100001;
            sine_reg0   <= 36'sb101101110001100111110011100111011001;
        end
        3702: begin
            cosine_reg0 <= 36'sb11010010101001100100100010000100011;
            sine_reg0   <= 36'sb101101110100001101001010011001110110;
        end
        3703: begin
            cosine_reg0 <= 36'sb11010010110111110101100011110000101;
            sine_reg0   <= 36'sb101101110110110010101100011010001011;
        end
        3704: begin
            cosine_reg0 <= 36'sb11010011000110000100100011011000000;
            sine_reg0   <= 36'sb101101111001011000011001100110110100;
        end
        3705: begin
            cosine_reg0 <= 36'sb11010011010100010001100000110001101;
            sine_reg0   <= 36'sb101101111011111110010001111110001000;
        end
        3706: begin
            cosine_reg0 <= 36'sb11010011100010011100011011110100111;
            sine_reg0   <= 36'sb101101111110100100010101011110100011;
        end
        3707: begin
            cosine_reg0 <= 36'sb11010011110000100101010100011000110;
            sine_reg0   <= 36'sb101110000001001010100100000110011110;
        end
        3708: begin
            cosine_reg0 <= 36'sb11010011111110101100001010010100111;
            sine_reg0   <= 36'sb101110000011110000111101110100010001;
        end
        3709: begin
            cosine_reg0 <= 36'sb11010100001100110000111101100000011;
            sine_reg0   <= 36'sb101110000110010111100010100110011000;
        end
        3710: begin
            cosine_reg0 <= 36'sb11010100011010110011101101110010100;
            sine_reg0   <= 36'sb101110001000111110010010011011001001;
        end
        3711: begin
            cosine_reg0 <= 36'sb11010100101000110100011011000010110;
            sine_reg0   <= 36'sb101110001011100101001101010001000000;
        end
        3712: begin
            cosine_reg0 <= 36'sb11010100110110110011000101001000011;
            sine_reg0   <= 36'sb101110001110001100010011000110010101;
        end
        3713: begin
            cosine_reg0 <= 36'sb11010101000100101111101011111010110;
            sine_reg0   <= 36'sb101110010000110011100011111001100000;
        end
        3714: begin
            cosine_reg0 <= 36'sb11010101010010101010001111010001010;
            sine_reg0   <= 36'sb101110010011011010111111101000111100;
        end
        3715: begin
            cosine_reg0 <= 36'sb11010101100000100010101111000011100;
            sine_reg0   <= 36'sb101110010110000010100110010010111111;
        end
        3716: begin
            cosine_reg0 <= 36'sb11010101101110011001001011001000101;
            sine_reg0   <= 36'sb101110011000101010010111110110000100;
        end
        3717: begin
            cosine_reg0 <= 36'sb11010101111100001101100011011000010;
            sine_reg0   <= 36'sb101110011011010010010100010000100010;
        end
        3718: begin
            cosine_reg0 <= 36'sb11010110001001111111110111101001111;
            sine_reg0   <= 36'sb101110011101111010011011100000110010;
        end
        3719: begin
            cosine_reg0 <= 36'sb11010110010111110000000111110100111;
            sine_reg0   <= 36'sb101110100000100010101101100101001100;
        end
        3720: begin
            cosine_reg0 <= 36'sb11010110100101011110010011110001000;
            sine_reg0   <= 36'sb101110100011001011001010011100001001;
        end
        3721: begin
            cosine_reg0 <= 36'sb11010110110011001010011011010101100;
            sine_reg0   <= 36'sb101110100101110011110010000100000000;
        end
        3722: begin
            cosine_reg0 <= 36'sb11010111000000110100011110011010001;
            sine_reg0   <= 36'sb101110101000011100100100011011001010;
        end
        3723: begin
            cosine_reg0 <= 36'sb11010111001110011100011100110110010;
            sine_reg0   <= 36'sb101110101011000101100001011111111110;
        end
        3724: begin
            cosine_reg0 <= 36'sb11010111011100000010010110100001110;
            sine_reg0   <= 36'sb101110101101101110101001010000110100;
        end
        3725: begin
            cosine_reg0 <= 36'sb11010111101001100110001011010100001;
            sine_reg0   <= 36'sb101110110000010111111011101100000100;
        end
        3726: begin
            cosine_reg0 <= 36'sb11010111110111000111111011000100111;
            sine_reg0   <= 36'sb101110110011000001011000110000000101;
        end
        3727: begin
            cosine_reg0 <= 36'sb11011000000100100111100101101011110;
            sine_reg0   <= 36'sb101110110101101011000000011011001111;
        end
        3728: begin
            cosine_reg0 <= 36'sb11011000010010000101001011000000100;
            sine_reg0   <= 36'sb101110111000010100110010101011111010;
        end
        3729: begin
            cosine_reg0 <= 36'sb11011000011111100000101010111010110;
            sine_reg0   <= 36'sb101110111010111110101111100000011100;
        end
        3730: begin
            cosine_reg0 <= 36'sb11011000101100111010000101010010010;
            sine_reg0   <= 36'sb101110111101101000110110110111001100;
        end
        3731: begin
            cosine_reg0 <= 36'sb11011000111010010001011001111110110;
            sine_reg0   <= 36'sb101111000000010011001000101110100011;
        end
        3732: begin
            cosine_reg0 <= 36'sb11011001000111100110101000110111111;
            sine_reg0   <= 36'sb101111000010111101100101000100110110;
        end
        3733: begin
            cosine_reg0 <= 36'sb11011001010100111001110001110101100;
            sine_reg0   <= 36'sb101111000101101000001011111000011101;
        end
        3734: begin
            cosine_reg0 <= 36'sb11011001100010001010110100101111100;
            sine_reg0   <= 36'sb101111001000010010111101000111101110;
        end
        3735: begin
            cosine_reg0 <= 36'sb11011001101111011001110001011101100;
            sine_reg0   <= 36'sb101111001010111101111000110001000000;
        end
        3736: begin
            cosine_reg0 <= 36'sb11011001111100100110100111110111100;
            sine_reg0   <= 36'sb101111001101101000111110110010101001;
        end
        3737: begin
            cosine_reg0 <= 36'sb11011010001001110001010111110101011;
            sine_reg0   <= 36'sb101111010000010100001111001011000001;
        end
        3738: begin
            cosine_reg0 <= 36'sb11011010010110111010000001001110111;
            sine_reg0   <= 36'sb101111010010111111101001111000011101;
        end
        3739: begin
            cosine_reg0 <= 36'sb11011010100100000000100011111011111;
            sine_reg0   <= 36'sb101111010101101011001110111001010011;
        end
        3740: begin
            cosine_reg0 <= 36'sb11011010110001000100111111110100100;
            sine_reg0   <= 36'sb101111011000010110111110001011111011;
        end
        3741: begin
            cosine_reg0 <= 36'sb11011010111110000111010100110000100;
            sine_reg0   <= 36'sb101111011011000010110111101110101001;
        end
        3742: begin
            cosine_reg0 <= 36'sb11011011001011000111100010100111111;
            sine_reg0   <= 36'sb101111011101101110111011011111110100;
        end
        3743: begin
            cosine_reg0 <= 36'sb11011011011000000101101001010010101;
            sine_reg0   <= 36'sb101111100000011011001001011101110010;
        end
        3744: begin
            cosine_reg0 <= 36'sb11011011100101000001101000101000101;
            sine_reg0   <= 36'sb101111100011000111100001100110111000;
        end
        3745: begin
            cosine_reg0 <= 36'sb11011011110001111011100000100010010;
            sine_reg0   <= 36'sb101111100101110100000011111001011100;
        end
        3746: begin
            cosine_reg0 <= 36'sb11011011111110110011010000110111001;
            sine_reg0   <= 36'sb101111101000100000110000010011110100;
        end
        3747: begin
            cosine_reg0 <= 36'sb11011100001011101000111001011111100;
            sine_reg0   <= 36'sb101111101011001101100110110100010101;
        end
        3748: begin
            cosine_reg0 <= 36'sb11011100011000011100011010010011100;
            sine_reg0   <= 36'sb101111101101111010100111011001010101;
        end
        3749: begin
            cosine_reg0 <= 36'sb11011100100101001101110011001011010;
            sine_reg0   <= 36'sb101111110000100111110010000001001001;
        end
        3750: begin
            cosine_reg0 <= 36'sb11011100110001111101000011111110101;
            sine_reg0   <= 36'sb101111110011010101000110101010000101;
        end
        3751: begin
            cosine_reg0 <= 36'sb11011100111110101010001100100110001;
            sine_reg0   <= 36'sb101111110110000010100101010010100000;
        end
        3752: begin
            cosine_reg0 <= 36'sb11011101001011010101001100111001101;
            sine_reg0   <= 36'sb101111111000110000001101111000101101;
        end
        3753: begin
            cosine_reg0 <= 36'sb11011101010111111110000100110001011;
            sine_reg0   <= 36'sb101111111011011110000000011011000011;
        end
        3754: begin
            cosine_reg0 <= 36'sb11011101100100100100110100000101101;
            sine_reg0   <= 36'sb101111111110001011111100110111110110;
        end
        3755: begin
            cosine_reg0 <= 36'sb11011101110001001001011010101110101;
            sine_reg0   <= 36'sb110000000000111010000011001101011010;
        end
        3756: begin
            cosine_reg0 <= 36'sb11011101111101101011111000100100100;
            sine_reg0   <= 36'sb110000000011101000010011011010000100;
        end
        3757: begin
            cosine_reg0 <= 36'sb11011110001010001100001101011111101;
            sine_reg0   <= 36'sb110000000110010110101101011100001000;
        end
        3758: begin
            cosine_reg0 <= 36'sb11011110010110101010011001011000010;
            sine_reg0   <= 36'sb110000001001000101010001010001111100;
        end
        3759: begin
            cosine_reg0 <= 36'sb11011110100011000110011100000110110;
            sine_reg0   <= 36'sb110000001011110011111110111001110011;
        end
        3760: begin
            cosine_reg0 <= 36'sb11011110101111100000010101100011011;
            sine_reg0   <= 36'sb110000001110100010110110010010000001;
        end
        3761: begin
            cosine_reg0 <= 36'sb11011110111011111000000101100110100;
            sine_reg0   <= 36'sb110000010001010001110111011000111100;
        end
        3762: begin
            cosine_reg0 <= 36'sb11011111001000001101101100001000011;
            sine_reg0   <= 36'sb110000010100000001000010001100110110;
        end
        3763: begin
            cosine_reg0 <= 36'sb11011111010100100001001001000001101;
            sine_reg0   <= 36'sb110000010110110000010110101100000011;
        end
        3764: begin
            cosine_reg0 <= 36'sb11011111100000110010011100001010100;
            sine_reg0   <= 36'sb110000011001011111110100110100111001;
        end
        3765: begin
            cosine_reg0 <= 36'sb11011111101101000001100101011011100;
            sine_reg0   <= 36'sb110000011100001111011100100101101001;
        end
        3766: begin
            cosine_reg0 <= 36'sb11011111111001001110100100101101000;
            sine_reg0   <= 36'sb110000011110111111001101111100101000;
        end
        3767: begin
            cosine_reg0 <= 36'sb11100000000101011001011001110111100;
            sine_reg0   <= 36'sb110000100001101111001000111000001011;
        end
        3768: begin
            cosine_reg0 <= 36'sb11100000010001100010000100110011100;
            sine_reg0   <= 36'sb110000100100011111001101010110100011;
        end
        3769: begin
            cosine_reg0 <= 36'sb11100000011101101000100101011001100;
            sine_reg0   <= 36'sb110000100111001111011011010110000100;
        end
        3770: begin
            cosine_reg0 <= 36'sb11100000101001101100111011100010001;
            sine_reg0   <= 36'sb110000101001111111110010110101000010;
        end
        3771: begin
            cosine_reg0 <= 36'sb11100000110101101111000111000101110;
            sine_reg0   <= 36'sb110000101100110000010011110001110000;
        end
        3772: begin
            cosine_reg0 <= 36'sb11100001000001101111000111111101001;
            sine_reg0   <= 36'sb110000101111100000111110001010100001;
        end
        3773: begin
            cosine_reg0 <= 36'sb11100001001101101100111110000000111;
            sine_reg0   <= 36'sb110000110010010001110001111101101001;
        end
        3774: begin
            cosine_reg0 <= 36'sb11100001011001101000101001001001100;
            sine_reg0   <= 36'sb110000110101000010101111001001011001;
        end
        3775: begin
            cosine_reg0 <= 36'sb11100001100101100010001001001111101;
            sine_reg0   <= 36'sb110000110111110011110101101100000101;
        end
        3776: begin
            cosine_reg0 <= 36'sb11100001110001011001011110001011111;
            sine_reg0   <= 36'sb110000111010100101000101100100000000;
        end
        3777: begin
            cosine_reg0 <= 36'sb11100001111101001110100111110111001;
            sine_reg0   <= 36'sb110000111101010110011110101111011100;
        end
        3778: begin
            cosine_reg0 <= 36'sb11100010001001000001100110001010000;
            sine_reg0   <= 36'sb110001000000001000000001001100101011;
        end
        3779: begin
            cosine_reg0 <= 36'sb11100010010100110010011000111101001;
            sine_reg0   <= 36'sb110001000010111001101100111010000001;
        end
        3780: begin
            cosine_reg0 <= 36'sb11100010100000100001000000001001010;
            sine_reg0   <= 36'sb110001000101101011100001110101110000;
        end
        3781: begin
            cosine_reg0 <= 36'sb11100010101100001101011011100111010;
            sine_reg0   <= 36'sb110001001000011101011111111110001010;
        end
        3782: begin
            cosine_reg0 <= 36'sb11100010110111110111101011001111111;
            sine_reg0   <= 36'sb110001001011001111100111010001100001;
        end
        3783: begin
            cosine_reg0 <= 36'sb11100011000011011111101110111011111;
            sine_reg0   <= 36'sb110001001110000001110111101110001000;
        end
        3784: begin
            cosine_reg0 <= 36'sb11100011001111000101100110100100001;
            sine_reg0   <= 36'sb110001010000110100010001010010010000;
        end
        3785: begin
            cosine_reg0 <= 36'sb11100011011010101001010010000001100;
            sine_reg0   <= 36'sb110001010011100110110011111100001011;
        end
        3786: begin
            cosine_reg0 <= 36'sb11100011100110001010110001001100111;
            sine_reg0   <= 36'sb110001010110011001011111101010001011;
        end
        3787: begin
            cosine_reg0 <= 36'sb11100011110001101010000011111111000;
            sine_reg0   <= 36'sb110001011001001100010100011010100011;
        end
        3788: begin
            cosine_reg0 <= 36'sb11100011111101000111001010010001000;
            sine_reg0   <= 36'sb110001011011111111010010001011100011;
        end
        3789: begin
            cosine_reg0 <= 36'sb11100100001000100010000011111011101;
            sine_reg0   <= 36'sb110001011110110010011000111011011110;
        end
        3790: begin
            cosine_reg0 <= 36'sb11100100010011111010110000111000000;
            sine_reg0   <= 36'sb110001100001100101101000101000100100;
        end
        3791: begin
            cosine_reg0 <= 36'sb11100100011111010001010000111110111;
            sine_reg0   <= 36'sb110001100100011001000001010001001000;
        end
        3792: begin
            cosine_reg0 <= 36'sb11100100101010100101100100001001100;
            sine_reg0   <= 36'sb110001100111001100100010110011011010;
        end
        3793: begin
            cosine_reg0 <= 36'sb11100100110101110111101010010000110;
            sine_reg0   <= 36'sb110001101010000000001101001101101100;
        end
        3794: begin
            cosine_reg0 <= 36'sb11100101000001000111100011001101110;
            sine_reg0   <= 36'sb110001101100110100000000011110010000;
        end
        3795: begin
            cosine_reg0 <= 36'sb11100101001100010101001110111001011;
            sine_reg0   <= 36'sb110001101111100111111100100011010101;
        end
        3796: begin
            cosine_reg0 <= 36'sb11100101010111100000101101001100111;
            sine_reg0   <= 36'sb110001110010011100000001011011001110;
        end
        3797: begin
            cosine_reg0 <= 36'sb11100101100010101001111110000001011;
            sine_reg0   <= 36'sb110001110101010000001111000100001010;
        end
        3798: begin
            cosine_reg0 <= 36'sb11100101101101110001000001001111111;
            sine_reg0   <= 36'sb110001111000000100100101011100011100;
        end
        3799: begin
            cosine_reg0 <= 36'sb11100101111000110101110110110001101;
            sine_reg0   <= 36'sb110001111010111001000100100010010011;
        end
        3800: begin
            cosine_reg0 <= 36'sb11100110000011111000011110011111110;
            sine_reg0   <= 36'sb110001111101101101101100010100000000;
        end
        3801: begin
            cosine_reg0 <= 36'sb11100110001110111000111000010011100;
            sine_reg0   <= 36'sb110010000000100010011100101111110101;
        end
        3802: begin
            cosine_reg0 <= 36'sb11100110011001110111000100000110000;
            sine_reg0   <= 36'sb110010000011010111010101110100000000;
        end
        3803: begin
            cosine_reg0 <= 36'sb11100110100100110011000001110000100;
            sine_reg0   <= 36'sb110010000110001100010111011110110100;
        end
        3804: begin
            cosine_reg0 <= 36'sb11100110101111101100110001001100010;
            sine_reg0   <= 36'sb110010001001000001100001101110100000;
        end
        3805: begin
            cosine_reg0 <= 36'sb11100110111010100100010010010010100;
            sine_reg0   <= 36'sb110010001011110110110100100001010100;
        end
        3806: begin
            cosine_reg0 <= 36'sb11100111000101011001100100111100110;
            sine_reg0   <= 36'sb110010001110101100001111110101100001;
        end
        3807: begin
            cosine_reg0 <= 36'sb11100111010000001100101001000100000;
            sine_reg0   <= 36'sb110010010001100001110011101001010110;
        end
        3808: begin
            cosine_reg0 <= 36'sb11100111011010111101011110100001110;
            sine_reg0   <= 36'sb110010010100010111011111111011000100;
        end
        3809: begin
            cosine_reg0 <= 36'sb11100111100101101100000101001111100;
            sine_reg0   <= 36'sb110010010111001101010100101000111011;
        end
        3810: begin
            cosine_reg0 <= 36'sb11100111110000011000011101000110011;
            sine_reg0   <= 36'sb110010011010000011010001110001001010;
        end
        3811: begin
            cosine_reg0 <= 36'sb11100111111011000010100101111111111;
            sine_reg0   <= 36'sb110010011100111001010111010010000001;
        end
        3812: begin
            cosine_reg0 <= 36'sb11101000000101101010011111110101100;
            sine_reg0   <= 36'sb110010011111101111100101001001110001;
        end
        3813: begin
            cosine_reg0 <= 36'sb11101000010000010000001010100000101;
            sine_reg0   <= 36'sb110010100010100101111011010110100111;
        end
        3814: begin
            cosine_reg0 <= 36'sb11101000011010110011100101111010110;
            sine_reg0   <= 36'sb110010100101011100011001110110110101;
        end
        3815: begin
            cosine_reg0 <= 36'sb11101000100101010100110001111101010;
            sine_reg0   <= 36'sb110010101000010011000000101000101001;
        end
        3816: begin
            cosine_reg0 <= 36'sb11101000101111110011101110100001111;
            sine_reg0   <= 36'sb110010101011001001101111101010010011;
        end
        3817: begin
            cosine_reg0 <= 36'sb11101000111010010000011011100001111;
            sine_reg0   <= 36'sb110010101110000000100110111010000010;
        end
        3818: begin
            cosine_reg0 <= 36'sb11101001000100101010111000110111001;
            sine_reg0   <= 36'sb110010110000110111100110010110000101;
        end
        3819: begin
            cosine_reg0 <= 36'sb11101001001111000011000110011010111;
            sine_reg0   <= 36'sb110010110011101110101101111100101100;
        end
        3820: begin
            cosine_reg0 <= 36'sb11101001011001011001000100000110111;
            sine_reg0   <= 36'sb110010110110100101111101101100000101;
        end
        3821: begin
            cosine_reg0 <= 36'sb11101001100011101100110001110100111;
            sine_reg0   <= 36'sb110010111001011101010101100010011111;
        end
        3822: begin
            cosine_reg0 <= 36'sb11101001101101111110001111011110010;
            sine_reg0   <= 36'sb110010111100010100110101011110001010;
        end
        3823: begin
            cosine_reg0 <= 36'sb11101001111000001101011100111100111;
            sine_reg0   <= 36'sb110010111111001100011101011101010100;
        end
        3824: begin
            cosine_reg0 <= 36'sb11101010000010011010011010001010011;
            sine_reg0   <= 36'sb110011000010000100001101011110001011;
        end
        3825: begin
            cosine_reg0 <= 36'sb11101010001100100101000111000000011;
            sine_reg0   <= 36'sb110011000100111100000101011110111111;
        end
        3826: begin
            cosine_reg0 <= 36'sb11101010010110101101100011011000101;
            sine_reg0   <= 36'sb110011000111110100000101011101111111;
        end
        3827: begin
            cosine_reg0 <= 36'sb11101010100000110011101111001101000;
            sine_reg0   <= 36'sb110011001010101100001101011001010111;
        end
        3828: begin
            cosine_reg0 <= 36'sb11101010101010110111101010010111001;
            sine_reg0   <= 36'sb110011001101100100011101001111011000;
        end
        3829: begin
            cosine_reg0 <= 36'sb11101010110100111001010100110001000;
            sine_reg0   <= 36'sb110011010000011100110100111110001111;
        end
        3830: begin
            cosine_reg0 <= 36'sb11101010111110111000101110010100001;
            sine_reg0   <= 36'sb110011010011010101010100100100001011;
        end
        3831: begin
            cosine_reg0 <= 36'sb11101011001000110101110110111010101;
            sine_reg0   <= 36'sb110011010110001101111011111111011001;
        end
        3832: begin
            cosine_reg0 <= 36'sb11101011010010110000101110011110010;
            sine_reg0   <= 36'sb110011011001000110101011001110001001;
        end
        3833: begin
            cosine_reg0 <= 36'sb11101011011100101001010100111000110;
            sine_reg0   <= 36'sb110011011011111111100010001110100111;
        end
        3834: begin
            cosine_reg0 <= 36'sb11101011100110011111101010000100010;
            sine_reg0   <= 36'sb110011011110111000100000111111000010;
        end
        3835: begin
            cosine_reg0 <= 36'sb11101011110000010011101101111010101;
            sine_reg0   <= 36'sb110011100001110001100111011101101001;
        end
        3836: begin
            cosine_reg0 <= 36'sb11101011111010000101100000010101101;
            sine_reg0   <= 36'sb110011100100101010110101101000100111;
        end
        3837: begin
            cosine_reg0 <= 36'sb11101100000011110101000001001111100;
            sine_reg0   <= 36'sb110011100111100100001011011110001100;
        end
        3838: begin
            cosine_reg0 <= 36'sb11101100001101100010010000100010000;
            sine_reg0   <= 36'sb110011101010011101101000111100100110;
        end
        3839: begin
            cosine_reg0 <= 36'sb11101100010111001101001110000111011;
            sine_reg0   <= 36'sb110011101101010111001110000010000001;
        end
        3840: begin
            cosine_reg0 <= 36'sb11101100100000110101111001111001100;
            sine_reg0   <= 36'sb110011110000010000111010101100101011;
        end
        3841: begin
            cosine_reg0 <= 36'sb11101100101010011100010011110010011;
            sine_reg0   <= 36'sb110011110011001010101110111010110001;
        end
        3842: begin
            cosine_reg0 <= 36'sb11101100110100000000011011101100010;
            sine_reg0   <= 36'sb110011110110000100101010101010100010;
        end
        3843: begin
            cosine_reg0 <= 36'sb11101100111101100010010001100001001;
            sine_reg0   <= 36'sb110011111000111110101101111010001010;
        end
        3844: begin
            cosine_reg0 <= 36'sb11101101000111000001110101001011001;
            sine_reg0   <= 36'sb110011111011111000111000100111110111;
        end
        3845: begin
            cosine_reg0 <= 36'sb11101101010000011111000110100100011;
            sine_reg0   <= 36'sb110011111110110011001010110001110101;
        end
        3846: begin
            cosine_reg0 <= 36'sb11101101011001111010000101100111001;
            sine_reg0   <= 36'sb110100000001101101100100010110010010;
        end
        3847: begin
            cosine_reg0 <= 36'sb11101101100011010010110010001101100;
            sine_reg0   <= 36'sb110100000100101000000101010011011011;
        end
        3848: begin
            cosine_reg0 <= 36'sb11101101101100101001001100010001101;
            sine_reg0   <= 36'sb110100000111100010101101100111011101;
        end
        3849: begin
            cosine_reg0 <= 36'sb11101101110101111101010011101110000;
            sine_reg0   <= 36'sb110100001010011101011101010000100100;
        end
        3850: begin
            cosine_reg0 <= 36'sb11101101111111001111001000011100100;
            sine_reg0   <= 36'sb110100001101011000010100001100111110;
        end
        3851: begin
            cosine_reg0 <= 36'sb11101110001000011110101010010111110;
            sine_reg0   <= 36'sb110100010000010011010010011010110111;
        end
        3852: begin
            cosine_reg0 <= 36'sb11101110010001101011111001011001111;
            sine_reg0   <= 36'sb110100010011001110010111111000011100;
        end
        3853: begin
            cosine_reg0 <= 36'sb11101110011010110110110101011101010;
            sine_reg0   <= 36'sb110100010110001001100100100011111001;
        end
        3854: begin
            cosine_reg0 <= 36'sb11101110100011111111011110011100010;
            sine_reg0   <= 36'sb110100011001000100111000011011011100;
        end
        3855: begin
            cosine_reg0 <= 36'sb11101110101101000101110100010001001;
            sine_reg0   <= 36'sb110100011100000000010011011101001111;
        end
        3856: begin
            cosine_reg0 <= 36'sb11101110110110001001110110110110010;
            sine_reg0   <= 36'sb110100011110111011110101100111100001;
        end
        3857: begin
            cosine_reg0 <= 36'sb11101110111111001011100110000110010;
            sine_reg0   <= 36'sb110100100001110111011110111000011101;
        end
        3858: begin
            cosine_reg0 <= 36'sb11101111001000001011000001111011010;
            sine_reg0   <= 36'sb110100100100110011001111001110001111;
        end
        3859: begin
            cosine_reg0 <= 36'sb11101111010001001000001010010000000;
            sine_reg0   <= 36'sb110100100111101111000110100111000100;
        end
        3860: begin
            cosine_reg0 <= 36'sb11101111011010000010111110111110111;
            sine_reg0   <= 36'sb110100101010101011000101000001000111;
        end
        3861: begin
            cosine_reg0 <= 36'sb11101111100010111011100000000010010;
            sine_reg0   <= 36'sb110100101101100111001010011010100110;
        end
        3862: begin
            cosine_reg0 <= 36'sb11101111101011110001101101010100110;
            sine_reg0   <= 36'sb110100110000100011010110110001101011;
        end
        3863: begin
            cosine_reg0 <= 36'sb11101111110100100101100110110000111;
            sine_reg0   <= 36'sb110100110011011111101010000100100010;
        end
        3864: begin
            cosine_reg0 <= 36'sb11101111111101010111001100010001010;
            sine_reg0   <= 36'sb110100110110011100000100010001011000;
        end
        3865: begin
            cosine_reg0 <= 36'sb11110000000110000110011101110000100;
            sine_reg0   <= 36'sb110100111001011000100101010110011001;
        end
        3866: begin
            cosine_reg0 <= 36'sb11110000001110110011011011001001001;
            sine_reg0   <= 36'sb110100111100010101001101010001101111;
        end
        3867: begin
            cosine_reg0 <= 36'sb11110000010111011110000100010101110;
            sine_reg0   <= 36'sb110100111111010001111100000001100111;
        end
        3868: begin
            cosine_reg0 <= 36'sb11110000100000000110011001010001001;
            sine_reg0   <= 36'sb110101000010001110110001100100001101;
        end
        3869: begin
            cosine_reg0 <= 36'sb11110000101000101100011001110101111;
            sine_reg0   <= 36'sb110101000101001011101101110111101010;
        end
        3870: begin
            cosine_reg0 <= 36'sb11110000110001010000000101111110110;
            sine_reg0   <= 36'sb110101001000001000110000111010001101;
        end
        3871: begin
            cosine_reg0 <= 36'sb11110000111001110001011101100110011;
            sine_reg0   <= 36'sb110101001011000101111010101001111110;
        end
        3872: begin
            cosine_reg0 <= 36'sb11110001000010010000100000100111101;
            sine_reg0   <= 36'sb110101001110000011001011000101001011;
        end
        3873: begin
            cosine_reg0 <= 36'sb11110001001010101101001110111101001;
            sine_reg0   <= 36'sb110101010001000000100010001001111110;
        end
        3874: begin
            cosine_reg0 <= 36'sb11110001010011000111101000100001101;
            sine_reg0   <= 36'sb110101010011111101111111110110100010;
        end
        3875: begin
            cosine_reg0 <= 36'sb11110001011011011111101101010000001;
            sine_reg0   <= 36'sb110101010110111011100100001001000010;
        end
        3876: begin
            cosine_reg0 <= 36'sb11110001100011110101011101000011011;
            sine_reg0   <= 36'sb110101011001111001001110111111101010;
        end
        3877: begin
            cosine_reg0 <= 36'sb11110001101100001000110111110110010;
            sine_reg0   <= 36'sb110101011100110111000000011000100101;
        end
        3878: begin
            cosine_reg0 <= 36'sb11110001110100011001111101100011101;
            sine_reg0   <= 36'sb110101011111110100111000010001111101;
        end
        3879: begin
            cosine_reg0 <= 36'sb11110001111100101000101110000110010;
            sine_reg0   <= 36'sb110101100010110010110110101001111110;
        end
        3880: begin
            cosine_reg0 <= 36'sb11110010000100110101001001011001010;
            sine_reg0   <= 36'sb110101100101110000111011011110110001;
        end
        3881: begin
            cosine_reg0 <= 36'sb11110010001100111111001111010111100;
            sine_reg0   <= 36'sb110101101000101111000110101110100011;
        end
        3882: begin
            cosine_reg0 <= 36'sb11110010010101000110111111111100000;
            sine_reg0   <= 36'sb110101101011101101011000010111011101;
        end
        3883: begin
            cosine_reg0 <= 36'sb11110010011101001100011011000001101;
            sine_reg0   <= 36'sb110101101110101011110000010111101010;
        end
        3884: begin
            cosine_reg0 <= 36'sb11110010100101001111100000100011100;
            sine_reg0   <= 36'sb110101110001101010001110101101010101;
        end
        3885: begin
            cosine_reg0 <= 36'sb11110010101101010000010000011100101;
            sine_reg0   <= 36'sb110101110100101000110011010110101001;
        end
        3886: begin
            cosine_reg0 <= 36'sb11110010110101001110101010101000000;
            sine_reg0   <= 36'sb110101110111100111011110010001101111;
        end
        3887: begin
            cosine_reg0 <= 36'sb11110010111101001010101111000000111;
            sine_reg0   <= 36'sb110101111010100110001111011100110011;
        end
        3888: begin
            cosine_reg0 <= 36'sb11110011000101000100011101100010001;
            sine_reg0   <= 36'sb110101111101100101000110110101111101;
        end
        3889: begin
            cosine_reg0 <= 36'sb11110011001100111011110110000111001;
            sine_reg0   <= 36'sb110110000000100100000100011011011010;
        end
        3890: begin
            cosine_reg0 <= 36'sb11110011010100110000111000101010110;
            sine_reg0   <= 36'sb110110000011100011001000001011010010;
        end
        3891: begin
            cosine_reg0 <= 36'sb11110011011100100011100101001000100;
            sine_reg0   <= 36'sb110110000110100010010010000011110001;
        end
        3892: begin
            cosine_reg0 <= 36'sb11110011100100010011111011011011010;
            sine_reg0   <= 36'sb110110001001100001100010000011000000;
        end
        3893: begin
            cosine_reg0 <= 36'sb11110011101100000001111011011110011;
            sine_reg0   <= 36'sb110110001100100000111000000111001001;
        end
        3894: begin
            cosine_reg0 <= 36'sb11110011110011101101100101001101000;
            sine_reg0   <= 36'sb110110001111100000010100001110010110;
        end
        3895: begin
            cosine_reg0 <= 36'sb11110011111011010110111000100010101;
            sine_reg0   <= 36'sb110110010010011111110110010110110001;
        end
        3896: begin
            cosine_reg0 <= 36'sb11110100000010111101110101011010010;
            sine_reg0   <= 36'sb110110010101011111011110011110100100;
        end
        3897: begin
            cosine_reg0 <= 36'sb11110100001010100010011011101111011;
            sine_reg0   <= 36'sb110110011000011111001100100011111001;
        end
        3898: begin
            cosine_reg0 <= 36'sb11110100010010000100101011011101010;
            sine_reg0   <= 36'sb110110011011011111000000100100111001;
        end
        3899: begin
            cosine_reg0 <= 36'sb11110100011001100100100100011111010;
            sine_reg0   <= 36'sb110110011110011110111010011111101111;
        end
        3900: begin
            cosine_reg0 <= 36'sb11110100100001000010000110110000111;
            sine_reg0   <= 36'sb110110100001011110111010010010100011;
        end
        3901: begin
            cosine_reg0 <= 36'sb11110100101000011101010010001101010;
            sine_reg0   <= 36'sb110110100100011110111111111011011111;
        end
        3902: begin
            cosine_reg0 <= 36'sb11110100101111110110000110101111111;
            sine_reg0   <= 36'sb110110100111011111001011011000101110;
        end
        3903: begin
            cosine_reg0 <= 36'sb11110100110111001100100100010100011;
            sine_reg0   <= 36'sb110110101010011111011100101000010111;
        end
        3904: begin
            cosine_reg0 <= 36'sb11110100111110100000101010110110001;
            sine_reg0   <= 36'sb110110101101011111110011101000100110;
        end
        3905: begin
            cosine_reg0 <= 36'sb11110101000101110010011010010000100;
            sine_reg0   <= 36'sb110110110000100000010000010111100010;
        end
        3906: begin
            cosine_reg0 <= 36'sb11110101001101000001110010011111001;
            sine_reg0   <= 36'sb110110110011100000110010110011010110;
        end
        3907: begin
            cosine_reg0 <= 36'sb11110101010100001110110011011101100;
            sine_reg0   <= 36'sb110110110110100001011010111010001010;
        end
        3908: begin
            cosine_reg0 <= 36'sb11110101011011011001011101000111001;
            sine_reg0   <= 36'sb110110111001100010001000101010001000;
        end
        3909: begin
            cosine_reg0 <= 36'sb11110101100010100001101111010111101;
            sine_reg0   <= 36'sb110110111100100010111100000001011001;
        end
        3910: begin
            cosine_reg0 <= 36'sb11110101101001100111101010001010110;
            sine_reg0   <= 36'sb110110111111100011110100111110000101;
        end
        3911: begin
            cosine_reg0 <= 36'sb11110101110000101011001101011011111;
            sine_reg0   <= 36'sb110111000010100100110011011110010111;
        end
        3912: begin
            cosine_reg0 <= 36'sb11110101110111101100011001000110111;
            sine_reg0   <= 36'sb110111000101100101110111100000010111;
        end
        3913: begin
            cosine_reg0 <= 36'sb11110101111110101011001101000111010;
            sine_reg0   <= 36'sb110111001000100111000001000010001101;
        end
        3914: begin
            cosine_reg0 <= 36'sb11110110000101100111101001011000110;
            sine_reg0   <= 36'sb110111001011101000010000000010000011;
        end
        3915: begin
            cosine_reg0 <= 36'sb11110110001100100001101101110111001;
            sine_reg0   <= 36'sb110111001110101001100100011110000010;
        end
        3916: begin
            cosine_reg0 <= 36'sb11110110010011011001011010011110000;
            sine_reg0   <= 36'sb110111010001101010111110010100010001;
        end
        3917: begin
            cosine_reg0 <= 36'sb11110110011010001110101111001001010;
            sine_reg0   <= 36'sb110111010100101100011101100010111011;
        end
        3918: begin
            cosine_reg0 <= 36'sb11110110100001000001101011110100101;
            sine_reg0   <= 36'sb110111010111101110000010001000000111;
        end
        3919: begin
            cosine_reg0 <= 36'sb11110110100111110010010000011100000;
            sine_reg0   <= 36'sb110111011010101111101100000001111111;
        end
        3920: begin
            cosine_reg0 <= 36'sb11110110101110100000011100111011001;
            sine_reg0   <= 36'sb110111011101110001011011001110101010;
        end
        3921: begin
            cosine_reg0 <= 36'sb11110110110101001100010001001101111;
            sine_reg0   <= 36'sb110111100000110011001111101100010001;
        end
        3922: begin
            cosine_reg0 <= 36'sb11110110111011110101101101010000001;
            sine_reg0   <= 36'sb110111100011110101001001011000111101;
        end
        3923: begin
            cosine_reg0 <= 36'sb11110111000010011100110000111101110;
            sine_reg0   <= 36'sb110111100110110111001000010010110110;
        end
        3924: begin
            cosine_reg0 <= 36'sb11110111001001000001011100010010110;
            sine_reg0   <= 36'sb110111101001111001001100011000000101;
        end
        3925: begin
            cosine_reg0 <= 36'sb11110111001111100011101111001010111;
            sine_reg0   <= 36'sb110111101100111011010101100110110001;
        end
        3926: begin
            cosine_reg0 <= 36'sb11110111010110000011101001100010011;
            sine_reg0   <= 36'sb110111101111111101100011111101000011;
        end
        3927: begin
            cosine_reg0 <= 36'sb11110111011100100001001011010101001;
            sine_reg0   <= 36'sb110111110010111111110111011001000011;
        end
        3928: begin
            cosine_reg0 <= 36'sb11110111100010111100010100011111000;
            sine_reg0   <= 36'sb110111110110000010001111111000111001;
        end
        3929: begin
            cosine_reg0 <= 36'sb11110111101001010101000100111100010;
            sine_reg0   <= 36'sb110111111001000100101101011010101110;
        end
        3930: begin
            cosine_reg0 <= 36'sb11110111101111101011011100101000110;
            sine_reg0   <= 36'sb110111111100000111001111111100101001;
        end
        3931: begin
            cosine_reg0 <= 36'sb11110111110101111111011011100000110;
            sine_reg0   <= 36'sb110111111111001001110111011100110010;
        end
        3932: begin
            cosine_reg0 <= 36'sb11110111111100010001000001100000010;
            sine_reg0   <= 36'sb111000000010001100100011111001010010;
        end
        3933: begin
            cosine_reg0 <= 36'sb11111000000010100000001110100011011;
            sine_reg0   <= 36'sb111000000101001111010101010000010000;
        end
        3934: begin
            cosine_reg0 <= 36'sb11111000001000101101000010100110011;
            sine_reg0   <= 36'sb111000001000010010001011011111110100;
        end
        3935: begin
            cosine_reg0 <= 36'sb11111000001110110111011101100101011;
            sine_reg0   <= 36'sb111000001011010101000110100110000110;
        end
        3936: begin
            cosine_reg0 <= 36'sb11111000010100111111011111011100100;
            sine_reg0   <= 36'sb111000001110011000000110100001001110;
        end
        3937: begin
            cosine_reg0 <= 36'sb11111000011011000101001000001000000;
            sine_reg0   <= 36'sb111000010001011011001011001111010011;
        end
        3938: begin
            cosine_reg0 <= 36'sb11111000100001001000010111100100001;
            sine_reg0   <= 36'sb111000010100011110010100101110011101;
        end
        3939: begin
            cosine_reg0 <= 36'sb11111000100111001001001101101101010;
            sine_reg0   <= 36'sb111000010111100001100010111100110100;
        end
        3940: begin
            cosine_reg0 <= 36'sb11111000101101000111101010011111101;
            sine_reg0   <= 36'sb111000011010100100110101111000011111;
        end
        3941: begin
            cosine_reg0 <= 36'sb11111000110011000011101101110111100;
            sine_reg0   <= 36'sb111000011101101000001101011111100110;
        end
        3942: begin
            cosine_reg0 <= 36'sb11111000111000111101010111110001001;
            sine_reg0   <= 36'sb111000100000101011101001110000010000;
        end
        3943: begin
            cosine_reg0 <= 36'sb11111000111110110100101000001001000;
            sine_reg0   <= 36'sb111000100011101111001010101000100101;
        end
        3944: begin
            cosine_reg0 <= 36'sb11111001000100101001011110111011101;
            sine_reg0   <= 36'sb111000100110110010110000000110101100;
        end
        3945: begin
            cosine_reg0 <= 36'sb11111001001010011011111100000101001;
            sine_reg0   <= 36'sb111000101001110110011010001000101100;
        end
        3946: begin
            cosine_reg0 <= 36'sb11111001010000001011111111100010001;
            sine_reg0   <= 36'sb111000101100111010001000101100101101;
        end
        3947: begin
            cosine_reg0 <= 36'sb11111001010101111001101001001110111;
            sine_reg0   <= 36'sb111000101111111101111011110000110111;
        end
        3948: begin
            cosine_reg0 <= 36'sb11111001011011100100111001001000001;
            sine_reg0   <= 36'sb111000110011000001110011010011001111;
        end
        3949: begin
            cosine_reg0 <= 36'sb11111001100001001101101111001010010;
            sine_reg0   <= 36'sb111000110110000101101111010001111110;
        end
        3950: begin
            cosine_reg0 <= 36'sb11111001100110110100001011010001110;
            sine_reg0   <= 36'sb111000111001001001101111101011001010;
        end
        3951: begin
            cosine_reg0 <= 36'sb11111001101100011000001101011011001;
            sine_reg0   <= 36'sb111000111100001101110100011100111011;
        end
        3952: begin
            cosine_reg0 <= 36'sb11111001110001111001110101100011000;
            sine_reg0   <= 36'sb111000111111010001111101100101011000;
        end
        3953: begin
            cosine_reg0 <= 36'sb11111001110111011001000011100110000;
            sine_reg0   <= 36'sb111001000010010110001011000010101000;
        end
        3954: begin
            cosine_reg0 <= 36'sb11111001111100110101110111100000110;
            sine_reg0   <= 36'sb111001000101011010011100110010110001;
        end
        3955: begin
            cosine_reg0 <= 36'sb11111010000010010000010001001111110;
            sine_reg0   <= 36'sb111001001000011110110010110011111011;
        end
        3956: begin
            cosine_reg0 <= 36'sb11111010000111101000010000101111111;
            sine_reg0   <= 36'sb111001001011100011001101000100001100;
        end
        3957: begin
            cosine_reg0 <= 36'sb11111010001100111101110101111101101;
            sine_reg0   <= 36'sb111001001110100111101011100001101100;
        end
        3958: begin
            cosine_reg0 <= 36'sb11111010010010010001000000110101110;
            sine_reg0   <= 36'sb111001010001101100001110001010100001;
        end
        3959: begin
            cosine_reg0 <= 36'sb11111010010111100001110001010101000;
            sine_reg0   <= 36'sb111001010100110000110100111100110010;
        end
        3960: begin
            cosine_reg0 <= 36'sb11111010011100110000000111011000010;
            sine_reg0   <= 36'sb111001010111110101011111110110100101;
        end
        3961: begin
            cosine_reg0 <= 36'sb11111010100001111100000010111100000;
            sine_reg0   <= 36'sb111001011010111010001110110110000010;
        end
        3962: begin
            cosine_reg0 <= 36'sb11111010100111000101100011111101011;
            sine_reg0   <= 36'sb111001011101111111000001111001001111;
        end
        3963: begin
            cosine_reg0 <= 36'sb11111010101100001100101010011000111;
            sine_reg0   <= 36'sb111001100001000011111000111110010010;
        end
        3964: begin
            cosine_reg0 <= 36'sb11111010110001010001010110001011101;
            sine_reg0   <= 36'sb111001100100001000110100000011010010;
        end
        3965: begin
            cosine_reg0 <= 36'sb11111010110110010011100111010010011;
            sine_reg0   <= 36'sb111001100111001101110011000110010111;
        end
        3966: begin
            cosine_reg0 <= 36'sb11111010111011010011011101101010000;
            sine_reg0   <= 36'sb111001101010010010110110000101100101;
        end
        3967: begin
            cosine_reg0 <= 36'sb11111011000000010000111001001111011;
            sine_reg0   <= 36'sb111001101101010111111100111111000100;
        end
        3968: begin
            cosine_reg0 <= 36'sb11111011000101001011111001111111101;
            sine_reg0   <= 36'sb111001110000011101000111110000111010;
        end
        3969: begin
            cosine_reg0 <= 36'sb11111011001010000100011111110111100;
            sine_reg0   <= 36'sb111001110011100010010110011001001101;
        end
        3970: begin
            cosine_reg0 <= 36'sb11111011001110111010101010110100001;
            sine_reg0   <= 36'sb111001110110100111101000110110000100;
        end
        3971: begin
            cosine_reg0 <= 36'sb11111011010011101110011010110010100;
            sine_reg0   <= 36'sb111001111001101100111111000101100101;
        end
        3972: begin
            cosine_reg0 <= 36'sb11111011011000011111101111101111100;
            sine_reg0   <= 36'sb111001111100110010011001000101110110;
        end
        3973: begin
            cosine_reg0 <= 36'sb11111011011101001110101001101000100;
            sine_reg0   <= 36'sb111001111111110111110110110100111110;
        end
        3974: begin
            cosine_reg0 <= 36'sb11111011100001111011001000011010010;
            sine_reg0   <= 36'sb111010000010111101011000010001000011;
        end
        3975: begin
            cosine_reg0 <= 36'sb11111011100110100101001100000010000;
            sine_reg0   <= 36'sb111010000110000010111101011000001011;
        end
        3976: begin
            cosine_reg0 <= 36'sb11111011101011001100110100011100111;
            sine_reg0   <= 36'sb111010001001001000100110001000011011;
        end
        3977: begin
            cosine_reg0 <= 36'sb11111011101111110010000001101000001;
            sine_reg0   <= 36'sb111010001100001110010010011111111011;
        end
        3978: begin
            cosine_reg0 <= 36'sb11111011110100010100110011100000110;
            sine_reg0   <= 36'sb111010001111010100000010011100110000;
        end
        3979: begin
            cosine_reg0 <= 36'sb11111011111000110101001010000100000;
            sine_reg0   <= 36'sb111010010010011001110101111101000000;
        end
        3980: begin
            cosine_reg0 <= 36'sb11111011111101010011000101001111001;
            sine_reg0   <= 36'sb111010010101011111101100111110110001;
        end
        3981: begin
            cosine_reg0 <= 36'sb11111100000001101110100100111111010;
            sine_reg0   <= 36'sb111010011000100101100111100000001001;
        end
        3982: begin
            cosine_reg0 <= 36'sb11111100000110000111101001010001111;
            sine_reg0   <= 36'sb111010011011101011100101011111001110;
        end
        3983: begin
            cosine_reg0 <= 36'sb11111100001010011110010010000100001;
            sine_reg0   <= 36'sb111010011110110001100110111010000111;
        end
        3984: begin
            cosine_reg0 <= 36'sb11111100001110110010011111010011011;
            sine_reg0   <= 36'sb111010100001110111101011101110110111;
        end
        3985: begin
            cosine_reg0 <= 36'sb11111100010011000100010000111101000;
            sine_reg0   <= 36'sb111010100100111101110011111011100111;
        end
        3986: begin
            cosine_reg0 <= 36'sb11111100010111010011100110111110010;
            sine_reg0   <= 36'sb111010101000000011111111011110011011;
        end
        3987: begin
            cosine_reg0 <= 36'sb11111100011011100000100001010100100;
            sine_reg0   <= 36'sb111010101011001010001110010101011001;
        end
        3988: begin
            cosine_reg0 <= 36'sb11111100011111101010111111111101011;
            sine_reg0   <= 36'sb111010101110010000100000011110100111;
        end
        3989: begin
            cosine_reg0 <= 36'sb11111100100011110011000010110110000;
            sine_reg0   <= 36'sb111010110001010110110101111000001010;
        end
        3990: begin
            cosine_reg0 <= 36'sb11111100100111111000101001111100000;
            sine_reg0   <= 36'sb111010110100011101001110100000001001;
        end
        3991: begin
            cosine_reg0 <= 36'sb11111100101011111011110101001100111;
            sine_reg0   <= 36'sb111010110111100011101010010100101000;
        end
        3992: begin
            cosine_reg0 <= 36'sb11111100101111111100100100100110001;
            sine_reg0   <= 36'sb111010111010101010001001010011101110;
        end
        3993: begin
            cosine_reg0 <= 36'sb11111100110011111010111000000101010;
            sine_reg0   <= 36'sb111010111101110000101011011011011111;
        end
        3994: begin
            cosine_reg0 <= 36'sb11111100110111110110101111100111110;
            sine_reg0   <= 36'sb111011000000110111010000101010000010;
        end
        3995: begin
            cosine_reg0 <= 36'sb11111100111011110000001011001011010;
            sine_reg0   <= 36'sb111011000011111101111000111101011101;
        end
        3996: begin
            cosine_reg0 <= 36'sb11111100111111100111001010101101010;
            sine_reg0   <= 36'sb111011000111000100100100010011110011;
        end
        3997: begin
            cosine_reg0 <= 36'sb11111101000011011011101110001011101;
            sine_reg0   <= 36'sb111011001010001011010010101011001100;
        end
        3998: begin
            cosine_reg0 <= 36'sb11111101000111001101110101100011110;
            sine_reg0   <= 36'sb111011001101010010000100000001101100;
        end
        3999: begin
            cosine_reg0 <= 36'sb11111101001010111101100000110011011;
            sine_reg0   <= 36'sb111011010000011000111000010101011000;
        end
        4000: begin
            cosine_reg0 <= 36'sb11111101001110101010101111111000001;
            sine_reg0   <= 36'sb111011010011011111101111100100010111;
        end
        4001: begin
            cosine_reg0 <= 36'sb11111101010010010101100010101111111;
            sine_reg0   <= 36'sb111011010110100110101001101100101101;
        end
        4002: begin
            cosine_reg0 <= 36'sb11111101010101111101111001011000010;
            sine_reg0   <= 36'sb111011011001101101100110101100100000;
        end
        4003: begin
            cosine_reg0 <= 36'sb11111101011001100011110011101111001;
            sine_reg0   <= 36'sb111011011100110100100110100001110101;
        end
        4004: begin
            cosine_reg0 <= 36'sb11111101011101000111010001110010001;
            sine_reg0   <= 36'sb111011011111111011101001001010110001;
        end
        4005: begin
            cosine_reg0 <= 36'sb11111101100000101000010011011111001;
            sine_reg0   <= 36'sb111011100011000010101110100101011010;
        end
        4006: begin
            cosine_reg0 <= 36'sb11111101100100000110111000110011111;
            sine_reg0   <= 36'sb111011100110001001110110101111110100;
        end
        4007: begin
            cosine_reg0 <= 36'sb11111101100111100011000001101110100;
            sine_reg0   <= 36'sb111011101001010001000001101000000101;
        end
        4008: begin
            cosine_reg0 <= 36'sb11111101101010111100101110001100100;
            sine_reg0   <= 36'sb111011101100011000001111001100010010;
        end
        4009: begin
            cosine_reg0 <= 36'sb11111101101110010011111110001100001;
            sine_reg0   <= 36'sb111011101111011111011111011010100001;
        end
        4010: begin
            cosine_reg0 <= 36'sb11111101110001101000110001101011001;
            sine_reg0   <= 36'sb111011110010100110110010010000110101;
        end
        4011: begin
            cosine_reg0 <= 36'sb11111101110100111011001000100111011;
            sine_reg0   <= 36'sb111011110101101110000111101101010101;
        end
        4012: begin
            cosine_reg0 <= 36'sb11111101111000001011000010111111000;
            sine_reg0   <= 36'sb111011111000110101011111101110000100;
        end
        4013: begin
            cosine_reg0 <= 36'sb11111101111011011000100000110000000;
            sine_reg0   <= 36'sb111011111011111100111010010001001010;
        end
        4014: begin
            cosine_reg0 <= 36'sb11111101111110100011100001111000010;
            sine_reg0   <= 36'sb111011111111000100010111010100101001;
        end
        4015: begin
            cosine_reg0 <= 36'sb11111110000001101100000110010101111;
            sine_reg0   <= 36'sb111100000010001011110110110110101000;
        end
        4016: begin
            cosine_reg0 <= 36'sb11111110000100110010001110000110111;
            sine_reg0   <= 36'sb111100000101010011011000110101001011;
        end
        4017: begin
            cosine_reg0 <= 36'sb11111110000111110101111001001001100;
            sine_reg0   <= 36'sb111100001000011010111101001110010111;
        end
        4018: begin
            cosine_reg0 <= 36'sb11111110001010110111000111011011110;
            sine_reg0   <= 36'sb111100001011100010100100000000010001;
        end
        4019: begin
            cosine_reg0 <= 36'sb11111110001101110101111000111011111;
            sine_reg0   <= 36'sb111100001110101010001101001000111110;
        end
        4020: begin
            cosine_reg0 <= 36'sb11111110010000110010001101100111111;
            sine_reg0   <= 36'sb111100010001110001111000100110100011;
        end
        4021: begin
            cosine_reg0 <= 36'sb11111110010011101100000101011110000;
            sine_reg0   <= 36'sb111100010100111001100110010111000100;
        end
        4022: begin
            cosine_reg0 <= 36'sb11111110010110100011100000011100011;
            sine_reg0   <= 36'sb111100011000000001010110011000100111;
        end
        4023: begin
            cosine_reg0 <= 36'sb11111110011001011000011110100001100;
            sine_reg0   <= 36'sb111100011011001001001000101001001111;
        end
        4024: begin
            cosine_reg0 <= 36'sb11111110011100001010111111101011010;
            sine_reg0   <= 36'sb111100011110010000111101000111000011;
        end
        4025: begin
            cosine_reg0 <= 36'sb11111110011110111011000011111000010;
            sine_reg0   <= 36'sb111100100001011000110011110000000111;
        end
        4026: begin
            cosine_reg0 <= 36'sb11111110100001101000101011000110101;
            sine_reg0   <= 36'sb111100100100100000101100100010011110;
        end
        4027: begin
            cosine_reg0 <= 36'sb11111110100100010011110101010100110;
            sine_reg0   <= 36'sb111100100111101000100111011100001111;
        end
        4028: begin
            cosine_reg0 <= 36'sb11111110100110111100100010100001000;
            sine_reg0   <= 36'sb111100101010110000100100011011011110;
        end
        4029: begin
            cosine_reg0 <= 36'sb11111110101001100010110010101001101;
            sine_reg0   <= 36'sb111100101101111000100011011110001111;
        end
        4030: begin
            cosine_reg0 <= 36'sb11111110101100000110100101101101001;
            sine_reg0   <= 36'sb111100110001000000100100100010100111;
        end
        4031: begin
            cosine_reg0 <= 36'sb11111110101110100111111011101001111;
            sine_reg0   <= 36'sb111100110100001000100111100110101011;
        end
        4032: begin
            cosine_reg0 <= 36'sb11111110110001000110110100011110011;
            sine_reg0   <= 36'sb111100110111010000101100101000011111;
        end
        4033: begin
            cosine_reg0 <= 36'sb11111110110011100011010000001001001;
            sine_reg0   <= 36'sb111100111010011000110011100110001000;
        end
        4034: begin
            cosine_reg0 <= 36'sb11111110110101111101001110101000100;
            sine_reg0   <= 36'sb111100111101100000111100011101101010;
        end
        4035: begin
            cosine_reg0 <= 36'sb11111110111000010100101111111011001;
            sine_reg0   <= 36'sb111101000000101001000111001101001010;
        end
        4036: begin
            cosine_reg0 <= 36'sb11111110111010101001110011111111011;
            sine_reg0   <= 36'sb111101000011110001010011110010101101;
        end
        4037: begin
            cosine_reg0 <= 36'sb11111110111100111100011010110100001;
            sine_reg0   <= 36'sb111101000110111001100010001100010111;
        end
        4038: begin
            cosine_reg0 <= 36'sb11111110111111001100100100010111101;
            sine_reg0   <= 36'sb111101001010000001110010011000001100;
        end
        4039: begin
            cosine_reg0 <= 36'sb11111111000001011010010000101000101;
            sine_reg0   <= 36'sb111101001101001010000100010100010010;
        end
        4040: begin
            cosine_reg0 <= 36'sb11111111000011100101011111100101110;
            sine_reg0   <= 36'sb111101010000010010010111111110101011;
        end
        4041: begin
            cosine_reg0 <= 36'sb11111111000101101110010001001101110;
            sine_reg0   <= 36'sb111101010011011010101101010101011110;
        end
        4042: begin
            cosine_reg0 <= 36'sb11111111000111110100100101011111001;
            sine_reg0   <= 36'sb111101010110100011000100010110101110;
        end
        4043: begin
            cosine_reg0 <= 36'sb11111111001001111000011100011000110;
            sine_reg0   <= 36'sb111101011001101011011101000000011111;
        end
        4044: begin
            cosine_reg0 <= 36'sb11111111001011111001110101111001011;
            sine_reg0   <= 36'sb111101011100110011110111010000110111;
        end
        4045: begin
            cosine_reg0 <= 36'sb11111111001101111000110001111111100;
            sine_reg0   <= 36'sb111101011111111100010011000101111001;
        end
        4046: begin
            cosine_reg0 <= 36'sb11111111001111110101010000101010001;
            sine_reg0   <= 36'sb111101100011000100110000011101101010;
        end
        4047: begin
            cosine_reg0 <= 36'sb11111111010001101111010001111000000;
            sine_reg0   <= 36'sb111101100110001101001111010110001110;
        end
        4048: begin
            cosine_reg0 <= 36'sb11111111010011100110110101100111111;
            sine_reg0   <= 36'sb111101101001010101101111101101101010;
        end
        4049: begin
            cosine_reg0 <= 36'sb11111111010101011011111011111000110;
            sine_reg0   <= 36'sb111101101100011110010001100010000001;
        end
        4050: begin
            cosine_reg0 <= 36'sb11111111010111001110100100101001011;
            sine_reg0   <= 36'sb111101101111100110110100110001011001;
        end
        4051: begin
            cosine_reg0 <= 36'sb11111111011000111110101111111000101;
            sine_reg0   <= 36'sb111101110010101111011001011001110101;
        end
        4052: begin
            cosine_reg0 <= 36'sb11111111011010101100011101100101101;
            sine_reg0   <= 36'sb111101110101110111111111011001011001;
        end
        4053: begin
            cosine_reg0 <= 36'sb11111111011100010111101101101111000;
            sine_reg0   <= 36'sb111101111001000000100110101110001011;
        end
        4054: begin
            cosine_reg0 <= 36'sb11111111011110000000100000010100000;
            sine_reg0   <= 36'sb111101111100001001001111010110001110;
        end
        4055: begin
            cosine_reg0 <= 36'sb11111111011111100110110101010011011;
            sine_reg0   <= 36'sb111101111111010001111001001111100110;
        end
        4056: begin
            cosine_reg0 <= 36'sb11111111100001001010101100101100011;
            sine_reg0   <= 36'sb111110000010011010100100011000011000;
        end
        4057: begin
            cosine_reg0 <= 36'sb11111111100010101100000110011101111;
            sine_reg0   <= 36'sb111110000101100011010000101110101000;
        end
        4058: begin
            cosine_reg0 <= 36'sb11111111100100001011000010100110111;
            sine_reg0   <= 36'sb111110001000101011111110010000011010;
        end
        4059: begin
            cosine_reg0 <= 36'sb11111111100101100111100001000110110;
            sine_reg0   <= 36'sb111110001011110100101100111011110010;
        end
        4060: begin
            cosine_reg0 <= 36'sb11111111100111000001100001111100010;
            sine_reg0   <= 36'sb111110001110111101011100101110110101;
        end
        4061: begin
            cosine_reg0 <= 36'sb11111111101000011001000101000110111;
            sine_reg0   <= 36'sb111110010010000110001101100111100110;
        end
        4062: begin
            cosine_reg0 <= 36'sb11111111101001101110001010100101011;
            sine_reg0   <= 36'sb111110010101001110111111100100001011;
        end
        4063: begin
            cosine_reg0 <= 36'sb11111111101011000000110010010111011;
            sine_reg0   <= 36'sb111110011000010111110010100010100110;
        end
        4064: begin
            cosine_reg0 <= 36'sb11111111101100010000111100011011101;
            sine_reg0   <= 36'sb111110011011100000100110100000111100;
        end
        4065: begin
            cosine_reg0 <= 36'sb11111111101101011110101000110001110;
            sine_reg0   <= 36'sb111110011110101001011011011101010001;
        end
        4066: begin
            cosine_reg0 <= 36'sb11111111101110101001110111011000110;
            sine_reg0   <= 36'sb111110100001110010010001010101101010;
        end
        4067: begin
            cosine_reg0 <= 36'sb11111111101111110010101000010000000;
            sine_reg0   <= 36'sb111110100100111011001000001000001010;
        end
        4068: begin
            cosine_reg0 <= 36'sb11111111110000111000111011010110110;
            sine_reg0   <= 36'sb111110101000000011111111110010110110;
        end
        4069: begin
            cosine_reg0 <= 36'sb11111111110001111100110000101100011;
            sine_reg0   <= 36'sb111110101011001100111000010011110001;
        end
        4070: begin
            cosine_reg0 <= 36'sb11111111110010111110001000010000001;
            sine_reg0   <= 36'sb111110101110010101110001101001000000;
        end
        4071: begin
            cosine_reg0 <= 36'sb11111111110011111101000010000001100;
            sine_reg0   <= 36'sb111110110001011110101011110000100111;
        end
        4072: begin
            cosine_reg0 <= 36'sb11111111110100111001011101111111111;
            sine_reg0   <= 36'sb111110110100100111100110101000101010;
        end
        4073: begin
            cosine_reg0 <= 36'sb11111111110101110011011100001010100;
            sine_reg0   <= 36'sb111110110111110000100010001111001100;
        end
        4074: begin
            cosine_reg0 <= 36'sb11111111110110101010111100100001000;
            sine_reg0   <= 36'sb111110111010111001011110100010010011;
        end
        4075: begin
            cosine_reg0 <= 36'sb11111111110111011111111111000010111;
            sine_reg0   <= 36'sb111110111110000010011011100000000010;
        end
        4076: begin
            cosine_reg0 <= 36'sb11111111111000010010100011101111011;
            sine_reg0   <= 36'sb111111000001001011011001000110011100;
        end
        4077: begin
            cosine_reg0 <= 36'sb11111111111001000010101010100110010;
            sine_reg0   <= 36'sb111111000100010100010111010011100111;
        end
        4078: begin
            cosine_reg0 <= 36'sb11111111111001110000010011100111000;
            sine_reg0   <= 36'sb111111000111011101010110000101100110;
        end
        4079: begin
            cosine_reg0 <= 36'sb11111111111010011011011110110001000;
            sine_reg0   <= 36'sb111111001010100110010101011010011101;
        end
        4080: begin
            cosine_reg0 <= 36'sb11111111111011000100001100000100000;
            sine_reg0   <= 36'sb111111001101101111010101010000010001;
        end
        4081: begin
            cosine_reg0 <= 36'sb11111111111011101010011011011111101;
            sine_reg0   <= 36'sb111111010000111000010101100101000100;
        end
        4082: begin
            cosine_reg0 <= 36'sb11111111111100001110001101000011011;
            sine_reg0   <= 36'sb111111010100000001010110010110111100;
        end
        4083: begin
            cosine_reg0 <= 36'sb11111111111100101111100000101111000;
            sine_reg0   <= 36'sb111111010111001010010111100011111100;
        end
        4084: begin
            cosine_reg0 <= 36'sb11111111111101001110010110100010010;
            sine_reg0   <= 36'sb111111011010010011011001001010001000;
        end
        4085: begin
            cosine_reg0 <= 36'sb11111111111101101010101110011100101;
            sine_reg0   <= 36'sb111111011101011100011011000111100101;
        end
        4086: begin
            cosine_reg0 <= 36'sb11111111111110000100101000011110000;
            sine_reg0   <= 36'sb111111100000100101011101011010010101;
        end
        4087: begin
            cosine_reg0 <= 36'sb11111111111110011100000100100110001;
            sine_reg0   <= 36'sb111111100011101110100000000000011110;
        end
        4088: begin
            cosine_reg0 <= 36'sb11111111111110110001000010110100110;
            sine_reg0   <= 36'sb111111100110110111100010111000000011;
        end
        4089: begin
            cosine_reg0 <= 36'sb11111111111111000011100011001001101;
            sine_reg0   <= 36'sb111111101010000000100101111111001000;
        end
        4090: begin
            cosine_reg0 <= 36'sb11111111111111010011100101100100101;
            sine_reg0   <= 36'sb111111101101001001101001010011110010;
        end
        4091: begin
            cosine_reg0 <= 36'sb11111111111111100001001010000101100;
            sine_reg0   <= 36'sb111111110000010010101100110100000011;
        end
        4092: begin
            cosine_reg0 <= 36'sb11111111111111101100010000101100011;
            sine_reg0   <= 36'sb111111110011011011110000011110000001;
        end
        4093: begin
            cosine_reg0 <= 36'sb11111111111111110100111001011000111;
            sine_reg0   <= 36'sb111111110110100100110100001111101111;
        end
        4094: begin
            cosine_reg0 <= 36'sb11111111111111111011000100001011000;
            sine_reg0   <= 36'sb111111111001101101111000000111010000;
        end
        default: begin
            cosine_reg0 <= 36'sb11111111111111111110110001000010101;
            sine_reg0   <= 36'sb111111111100110110111100000010101010;
        end
        endcase
        // Compute residual (value not obtained from table * 2*pi) // unsigned mult okay
        // residual_reg0 <= phase_accum[32-12-1:0] * 16'b110010010000111111;
    end
end

// Perform Correction
logic signed [WIDTH-1:0]                cosine_reg1;
logic signed [WIDTH-1:0]                sine_reg1;
// logic signed [RESIDUAL_WIDTH-1:0]       residual_reg1;

logic signed [WIDTH-1:0]                cosine_reg2;
logic signed [WIDTH-1:0]                sine_reg2;

always_ff @ (posedge i_clock) begin
    if (i_ready == 1'b1) begin
        // Pipeline Stage 1
        cosine_reg1 <= cosine_reg0;
        sine_reg1 <= sine_reg0;
        // residual_reg1 <= (residual_reg0[12+RESIDUAL_WIDTH-1:11] + 1'b1) >> 1;
        // Pipeline Stage 2
        cosine_reg2 <= cosine_reg1;
        sine_reg2 <= sine_reg1;

        // Pipeline Stage 3
        o_cosine_data <= cosine_reg2;
        o_sine_data <= sine_reg2;
    end
end

endmodule: chmod_dds

`default_nettype wire
