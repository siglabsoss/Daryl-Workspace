// Generated from template at 01/31/2017
`timescale 10ps / 10ps

`default_nettype none

module ldpc_column_to_row_rom #(
	parameter integer INPUT_LENGTH = 1152,
    parameter integer EXPANSION_FACTOR = 96
) (
    input  wire logic                                   i_valid,
    output      logic [$clog2(12*EXPANSION_FACTOR)-1:0] o_index_for_a0,
    output      logic [$clog2(12*EXPANSION_FACTOR)-1:0] o_index_for_a1,
    output      logic [$clog2(12*EXPANSION_FACTOR)-1:0] o_index_for_a2,
    output      logic [$clog2(12*EXPANSION_FACTOR)-1:0] o_index_for_a3,
    output      logic [$clog2(12*EXPANSION_FACTOR)-1:0] o_index_for_a4,
    output      logic [$clog2(12*EXPANSION_FACTOR)-1:0] o_index_for_a5, 
    output      logic [$clog2(8)-1:0]                   o_branch_for_a0,
    output      logic [$clog2(8)-1:0]                   o_branch_for_a1,
    output      logic [$clog2(8)-1:0]                   o_branch_for_a2,
    output      logic [$clog2(8)-1:0]                   o_branch_for_a3,
    output      logic [$clog2(8)-1:0]                   o_branch_for_a4,
    output      logic [$clog2(8)-1:0]                   o_branch_for_a5,
    input  wire logic                                   i_clock,
	input  wire logic                                   i_reset
);

logic [$clog2(INPUT_LENGTH)-1:0] count;

always_ff @(posedge i_clock) begin
    if (i_reset == 1'b1) begin
        count <= 0;
    end else if (i_valid) begin
        if (count == INPUT_LENGTH-1) begin
            count <= 0;
        end else begin
            count <= count + 1;
        end
    end

    case (count)
    0: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 349;
        o_index_for_a1 <= 780;
        o_index_for_a2 <= 1099;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 350;
        o_index_for_a1 <= 781;
        o_index_for_a2 <= 1100;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 351;
        o_index_for_a1 <= 782;
        o_index_for_a2 <= 1101;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    3: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 352;
        o_index_for_a1 <= 783;
        o_index_for_a2 <= 1102;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    4: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 353;
        o_index_for_a1 <= 784;
        o_index_for_a2 <= 1103;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    5: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 354;
        o_index_for_a1 <= 785;
        o_index_for_a2 <= 1104;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    6: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 355;
        o_index_for_a1 <= 786;
        o_index_for_a2 <= 1105;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    7: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 356;
        o_index_for_a1 <= 787;
        o_index_for_a2 <= 1106;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    8: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 357;
        o_index_for_a1 <= 788;
        o_index_for_a2 <= 1107;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    9: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 358;
        o_index_for_a1 <= 789;
        o_index_for_a2 <= 1108;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    10: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 359;
        o_index_for_a1 <= 790;
        o_index_for_a2 <= 1109;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    11: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 360;
        o_index_for_a1 <= 791;
        o_index_for_a2 <= 1110;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    12: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 361;
        o_index_for_a1 <= 792;
        o_index_for_a2 <= 1111;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    13: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 362;
        o_index_for_a1 <= 793;
        o_index_for_a2 <= 1112;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    14: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 363;
        o_index_for_a1 <= 794;
        o_index_for_a2 <= 1113;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    15: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 364;
        o_index_for_a1 <= 795;
        o_index_for_a2 <= 1114;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    16: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 365;
        o_index_for_a1 <= 796;
        o_index_for_a2 <= 1115;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    17: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 366;
        o_index_for_a1 <= 797;
        o_index_for_a2 <= 1116;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    18: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 367;
        o_index_for_a1 <= 798;
        o_index_for_a2 <= 1117;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    19: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 368;
        o_index_for_a1 <= 799;
        o_index_for_a2 <= 1118;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    20: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 369;
        o_index_for_a1 <= 800;
        o_index_for_a2 <= 1119;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    21: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 370;
        o_index_for_a1 <= 801;
        o_index_for_a2 <= 1120;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    22: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 371;
        o_index_for_a1 <= 802;
        o_index_for_a2 <= 1121;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    23: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 372;
        o_index_for_a1 <= 803;
        o_index_for_a2 <= 1122;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    24: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 373;
        o_index_for_a1 <= 804;
        o_index_for_a2 <= 1123;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    25: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 374;
        o_index_for_a1 <= 805;
        o_index_for_a2 <= 1124;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    26: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 375;
        o_index_for_a1 <= 806;
        o_index_for_a2 <= 1125;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    27: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 376;
        o_index_for_a1 <= 807;
        o_index_for_a2 <= 1126;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    28: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 377;
        o_index_for_a1 <= 808;
        o_index_for_a2 <= 1127;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    29: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 378;
        o_index_for_a1 <= 809;
        o_index_for_a2 <= 1128;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    30: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 379;
        o_index_for_a1 <= 810;
        o_index_for_a2 <= 1129;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    31: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 380;
        o_index_for_a1 <= 811;
        o_index_for_a2 <= 1130;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    32: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 381;
        o_index_for_a1 <= 812;
        o_index_for_a2 <= 1131;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    33: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 382;
        o_index_for_a1 <= 813;
        o_index_for_a2 <= 1132;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    34: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 383;
        o_index_for_a1 <= 814;
        o_index_for_a2 <= 1133;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    35: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 288;
        o_index_for_a1 <= 815;
        o_index_for_a2 <= 1134;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    36: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 289;
        o_index_for_a1 <= 816;
        o_index_for_a2 <= 1135;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    37: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 290;
        o_index_for_a1 <= 817;
        o_index_for_a2 <= 1136;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    38: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 291;
        o_index_for_a1 <= 818;
        o_index_for_a2 <= 1137;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    39: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 292;
        o_index_for_a1 <= 819;
        o_index_for_a2 <= 1138;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    40: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 293;
        o_index_for_a1 <= 820;
        o_index_for_a2 <= 1139;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    41: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 294;
        o_index_for_a1 <= 821;
        o_index_for_a2 <= 1140;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    42: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 295;
        o_index_for_a1 <= 822;
        o_index_for_a2 <= 1141;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    43: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 296;
        o_index_for_a1 <= 823;
        o_index_for_a2 <= 1142;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    44: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 297;
        o_index_for_a1 <= 824;
        o_index_for_a2 <= 1143;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    45: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 298;
        o_index_for_a1 <= 825;
        o_index_for_a2 <= 1144;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    46: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 299;
        o_index_for_a1 <= 826;
        o_index_for_a2 <= 1145;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    47: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 300;
        o_index_for_a1 <= 827;
        o_index_for_a2 <= 1146;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    48: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 301;
        o_index_for_a1 <= 828;
        o_index_for_a2 <= 1147;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    49: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 302;
        o_index_for_a1 <= 829;
        o_index_for_a2 <= 1148;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    50: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 303;
        o_index_for_a1 <= 830;
        o_index_for_a2 <= 1149;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    51: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 304;
        o_index_for_a1 <= 831;
        o_index_for_a2 <= 1150;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    52: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 305;
        o_index_for_a1 <= 832;
        o_index_for_a2 <= 1151;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    53: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 306;
        o_index_for_a1 <= 833;
        o_index_for_a2 <= 1056;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    54: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 307;
        o_index_for_a1 <= 834;
        o_index_for_a2 <= 1057;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    55: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 308;
        o_index_for_a1 <= 835;
        o_index_for_a2 <= 1058;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    56: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 309;
        o_index_for_a1 <= 836;
        o_index_for_a2 <= 1059;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    57: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 310;
        o_index_for_a1 <= 837;
        o_index_for_a2 <= 1060;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    58: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 311;
        o_index_for_a1 <= 838;
        o_index_for_a2 <= 1061;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    59: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 312;
        o_index_for_a1 <= 839;
        o_index_for_a2 <= 1062;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    60: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 313;
        o_index_for_a1 <= 840;
        o_index_for_a2 <= 1063;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    61: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 314;
        o_index_for_a1 <= 841;
        o_index_for_a2 <= 1064;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    62: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 315;
        o_index_for_a1 <= 842;
        o_index_for_a2 <= 1065;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    63: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 316;
        o_index_for_a1 <= 843;
        o_index_for_a2 <= 1066;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    64: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 317;
        o_index_for_a1 <= 844;
        o_index_for_a2 <= 1067;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    65: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 318;
        o_index_for_a1 <= 845;
        o_index_for_a2 <= 1068;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    66: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 319;
        o_index_for_a1 <= 846;
        o_index_for_a2 <= 1069;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    67: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 320;
        o_index_for_a1 <= 847;
        o_index_for_a2 <= 1070;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    68: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 321;
        o_index_for_a1 <= 848;
        o_index_for_a2 <= 1071;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    69: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 322;
        o_index_for_a1 <= 849;
        o_index_for_a2 <= 1072;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    70: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 323;
        o_index_for_a1 <= 850;
        o_index_for_a2 <= 1073;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    71: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 324;
        o_index_for_a1 <= 851;
        o_index_for_a2 <= 1074;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    72: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 325;
        o_index_for_a1 <= 852;
        o_index_for_a2 <= 1075;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    73: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 326;
        o_index_for_a1 <= 853;
        o_index_for_a2 <= 1076;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    74: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 327;
        o_index_for_a1 <= 854;
        o_index_for_a2 <= 1077;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    75: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 328;
        o_index_for_a1 <= 855;
        o_index_for_a2 <= 1078;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    76: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 329;
        o_index_for_a1 <= 856;
        o_index_for_a2 <= 1079;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    77: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 330;
        o_index_for_a1 <= 857;
        o_index_for_a2 <= 1080;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    78: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 331;
        o_index_for_a1 <= 858;
        o_index_for_a2 <= 1081;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    79: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 332;
        o_index_for_a1 <= 859;
        o_index_for_a2 <= 1082;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    80: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 333;
        o_index_for_a1 <= 860;
        o_index_for_a2 <= 1083;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    81: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 334;
        o_index_for_a1 <= 861;
        o_index_for_a2 <= 1084;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    82: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 335;
        o_index_for_a1 <= 862;
        o_index_for_a2 <= 1085;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    83: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 336;
        o_index_for_a1 <= 863;
        o_index_for_a2 <= 1086;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    84: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 337;
        o_index_for_a1 <= 768;
        o_index_for_a2 <= 1087;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    85: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 338;
        o_index_for_a1 <= 769;
        o_index_for_a2 <= 1088;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    86: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 339;
        o_index_for_a1 <= 770;
        o_index_for_a2 <= 1089;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    87: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 340;
        o_index_for_a1 <= 771;
        o_index_for_a2 <= 1090;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    88: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 341;
        o_index_for_a1 <= 772;
        o_index_for_a2 <= 1091;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    89: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 342;
        o_index_for_a1 <= 773;
        o_index_for_a2 <= 1092;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    90: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 343;
        o_index_for_a1 <= 774;
        o_index_for_a2 <= 1093;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    91: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 344;
        o_index_for_a1 <= 775;
        o_index_for_a2 <= 1094;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    92: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 345;
        o_index_for_a1 <= 776;
        o_index_for_a2 <= 1095;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    93: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 346;
        o_index_for_a1 <= 777;
        o_index_for_a2 <= 1096;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    94: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 347;
        o_index_for_a1 <= 778;
        o_index_for_a2 <= 1097;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    95: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 348;
        o_index_for_a1 <= 779;
        o_index_for_a2 <= 1098;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    96: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 94;
        o_index_for_a1 <= 123;
        o_index_for_a2 <= 683;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    97: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 95;
        o_index_for_a1 <= 124;
        o_index_for_a2 <= 684;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    98: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 0;
        o_index_for_a1 <= 125;
        o_index_for_a2 <= 685;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    99: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1;
        o_index_for_a1 <= 126;
        o_index_for_a2 <= 686;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    100: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 2;
        o_index_for_a1 <= 127;
        o_index_for_a2 <= 687;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    101: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 3;
        o_index_for_a1 <= 128;
        o_index_for_a2 <= 688;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    102: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 4;
        o_index_for_a1 <= 129;
        o_index_for_a2 <= 689;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    103: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 5;
        o_index_for_a1 <= 130;
        o_index_for_a2 <= 690;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    104: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 6;
        o_index_for_a1 <= 131;
        o_index_for_a2 <= 691;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    105: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 7;
        o_index_for_a1 <= 132;
        o_index_for_a2 <= 692;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    106: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 8;
        o_index_for_a1 <= 133;
        o_index_for_a2 <= 693;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    107: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 9;
        o_index_for_a1 <= 134;
        o_index_for_a2 <= 694;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    108: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 10;
        o_index_for_a1 <= 135;
        o_index_for_a2 <= 695;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    109: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 11;
        o_index_for_a1 <= 136;
        o_index_for_a2 <= 696;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    110: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 12;
        o_index_for_a1 <= 137;
        o_index_for_a2 <= 697;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    111: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 13;
        o_index_for_a1 <= 138;
        o_index_for_a2 <= 698;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    112: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 14;
        o_index_for_a1 <= 139;
        o_index_for_a2 <= 699;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    113: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 15;
        o_index_for_a1 <= 140;
        o_index_for_a2 <= 700;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    114: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 16;
        o_index_for_a1 <= 141;
        o_index_for_a2 <= 701;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    115: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 17;
        o_index_for_a1 <= 142;
        o_index_for_a2 <= 702;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    116: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 18;
        o_index_for_a1 <= 143;
        o_index_for_a2 <= 703;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    117: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 19;
        o_index_for_a1 <= 144;
        o_index_for_a2 <= 704;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    118: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 20;
        o_index_for_a1 <= 145;
        o_index_for_a2 <= 705;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    119: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 21;
        o_index_for_a1 <= 146;
        o_index_for_a2 <= 706;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    120: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 22;
        o_index_for_a1 <= 147;
        o_index_for_a2 <= 707;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    121: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 23;
        o_index_for_a1 <= 148;
        o_index_for_a2 <= 708;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    122: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 24;
        o_index_for_a1 <= 149;
        o_index_for_a2 <= 709;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    123: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 25;
        o_index_for_a1 <= 150;
        o_index_for_a2 <= 710;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    124: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 26;
        o_index_for_a1 <= 151;
        o_index_for_a2 <= 711;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    125: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 27;
        o_index_for_a1 <= 152;
        o_index_for_a2 <= 712;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    126: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 28;
        o_index_for_a1 <= 153;
        o_index_for_a2 <= 713;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    127: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 29;
        o_index_for_a1 <= 154;
        o_index_for_a2 <= 714;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    128: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 30;
        o_index_for_a1 <= 155;
        o_index_for_a2 <= 715;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    129: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 31;
        o_index_for_a1 <= 156;
        o_index_for_a2 <= 716;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    130: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 32;
        o_index_for_a1 <= 157;
        o_index_for_a2 <= 717;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    131: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 33;
        o_index_for_a1 <= 158;
        o_index_for_a2 <= 718;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    132: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 34;
        o_index_for_a1 <= 159;
        o_index_for_a2 <= 719;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    133: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 35;
        o_index_for_a1 <= 160;
        o_index_for_a2 <= 720;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    134: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 36;
        o_index_for_a1 <= 161;
        o_index_for_a2 <= 721;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    135: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 37;
        o_index_for_a1 <= 162;
        o_index_for_a2 <= 722;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    136: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 38;
        o_index_for_a1 <= 163;
        o_index_for_a2 <= 723;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    137: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 39;
        o_index_for_a1 <= 164;
        o_index_for_a2 <= 724;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    138: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 40;
        o_index_for_a1 <= 165;
        o_index_for_a2 <= 725;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    139: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 41;
        o_index_for_a1 <= 166;
        o_index_for_a2 <= 726;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    140: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 42;
        o_index_for_a1 <= 167;
        o_index_for_a2 <= 727;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    141: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 43;
        o_index_for_a1 <= 168;
        o_index_for_a2 <= 728;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    142: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 44;
        o_index_for_a1 <= 169;
        o_index_for_a2 <= 729;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    143: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 45;
        o_index_for_a1 <= 170;
        o_index_for_a2 <= 730;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    144: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 46;
        o_index_for_a1 <= 171;
        o_index_for_a2 <= 731;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    145: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 47;
        o_index_for_a1 <= 172;
        o_index_for_a2 <= 732;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    146: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 48;
        o_index_for_a1 <= 173;
        o_index_for_a2 <= 733;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    147: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 49;
        o_index_for_a1 <= 174;
        o_index_for_a2 <= 734;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    148: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 50;
        o_index_for_a1 <= 175;
        o_index_for_a2 <= 735;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    149: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 51;
        o_index_for_a1 <= 176;
        o_index_for_a2 <= 736;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    150: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 52;
        o_index_for_a1 <= 177;
        o_index_for_a2 <= 737;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    151: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 53;
        o_index_for_a1 <= 178;
        o_index_for_a2 <= 738;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    152: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 54;
        o_index_for_a1 <= 179;
        o_index_for_a2 <= 739;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    153: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 55;
        o_index_for_a1 <= 180;
        o_index_for_a2 <= 740;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    154: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 56;
        o_index_for_a1 <= 181;
        o_index_for_a2 <= 741;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    155: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 57;
        o_index_for_a1 <= 182;
        o_index_for_a2 <= 742;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    156: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 58;
        o_index_for_a1 <= 183;
        o_index_for_a2 <= 743;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    157: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 59;
        o_index_for_a1 <= 184;
        o_index_for_a2 <= 744;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    158: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 60;
        o_index_for_a1 <= 185;
        o_index_for_a2 <= 745;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    159: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 61;
        o_index_for_a1 <= 186;
        o_index_for_a2 <= 746;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    160: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 62;
        o_index_for_a1 <= 187;
        o_index_for_a2 <= 747;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    161: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 63;
        o_index_for_a1 <= 188;
        o_index_for_a2 <= 748;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    162: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 64;
        o_index_for_a1 <= 189;
        o_index_for_a2 <= 749;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    163: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 65;
        o_index_for_a1 <= 190;
        o_index_for_a2 <= 750;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    164: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 66;
        o_index_for_a1 <= 191;
        o_index_for_a2 <= 751;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    165: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 67;
        o_index_for_a1 <= 96;
        o_index_for_a2 <= 752;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    166: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 68;
        o_index_for_a1 <= 97;
        o_index_for_a2 <= 753;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    167: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 69;
        o_index_for_a1 <= 98;
        o_index_for_a2 <= 754;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    168: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 70;
        o_index_for_a1 <= 99;
        o_index_for_a2 <= 755;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    169: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 71;
        o_index_for_a1 <= 100;
        o_index_for_a2 <= 756;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    170: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 72;
        o_index_for_a1 <= 101;
        o_index_for_a2 <= 757;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    171: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 73;
        o_index_for_a1 <= 102;
        o_index_for_a2 <= 758;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    172: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 74;
        o_index_for_a1 <= 103;
        o_index_for_a2 <= 759;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    173: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 75;
        o_index_for_a1 <= 104;
        o_index_for_a2 <= 760;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    174: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 76;
        o_index_for_a1 <= 105;
        o_index_for_a2 <= 761;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    175: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 77;
        o_index_for_a1 <= 106;
        o_index_for_a2 <= 762;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    176: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 78;
        o_index_for_a1 <= 107;
        o_index_for_a2 <= 763;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    177: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 79;
        o_index_for_a1 <= 108;
        o_index_for_a2 <= 764;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    178: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 80;
        o_index_for_a1 <= 109;
        o_index_for_a2 <= 765;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    179: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 81;
        o_index_for_a1 <= 110;
        o_index_for_a2 <= 766;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    180: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 82;
        o_index_for_a1 <= 111;
        o_index_for_a2 <= 767;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    181: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 83;
        o_index_for_a1 <= 112;
        o_index_for_a2 <= 672;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    182: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 84;
        o_index_for_a1 <= 113;
        o_index_for_a2 <= 673;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    183: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 85;
        o_index_for_a1 <= 114;
        o_index_for_a2 <= 674;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    184: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 86;
        o_index_for_a1 <= 115;
        o_index_for_a2 <= 675;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    185: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 87;
        o_index_for_a1 <= 116;
        o_index_for_a2 <= 676;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    186: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 88;
        o_index_for_a1 <= 117;
        o_index_for_a2 <= 677;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    187: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 89;
        o_index_for_a1 <= 118;
        o_index_for_a2 <= 678;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    188: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 90;
        o_index_for_a1 <= 119;
        o_index_for_a2 <= 679;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    189: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 91;
        o_index_for_a1 <= 120;
        o_index_for_a2 <= 680;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    190: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 92;
        o_index_for_a1 <= 121;
        o_index_for_a2 <= 681;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    191: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 93;
        o_index_for_a1 <= 122;
        o_index_for_a2 <= 682;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    192: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 73;
        o_index_for_a1 <= 335;
        o_index_for_a2 <= 423;
        o_index_for_a3 <= 671;
        o_index_for_a4 <= 745;
        o_index_for_a5 <= 967; 
    end
    193: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 74;
        o_index_for_a1 <= 336;
        o_index_for_a2 <= 424;
        o_index_for_a3 <= 576;
        o_index_for_a4 <= 746;
        o_index_for_a5 <= 968; 
    end
    194: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 75;
        o_index_for_a1 <= 337;
        o_index_for_a2 <= 425;
        o_index_for_a3 <= 577;
        o_index_for_a4 <= 747;
        o_index_for_a5 <= 969; 
    end
    195: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 76;
        o_index_for_a1 <= 338;
        o_index_for_a2 <= 426;
        o_index_for_a3 <= 578;
        o_index_for_a4 <= 748;
        o_index_for_a5 <= 970; 
    end
    196: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 77;
        o_index_for_a1 <= 339;
        o_index_for_a2 <= 427;
        o_index_for_a3 <= 579;
        o_index_for_a4 <= 749;
        o_index_for_a5 <= 971; 
    end
    197: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 78;
        o_index_for_a1 <= 340;
        o_index_for_a2 <= 428;
        o_index_for_a3 <= 580;
        o_index_for_a4 <= 750;
        o_index_for_a5 <= 972; 
    end
    198: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 79;
        o_index_for_a1 <= 341;
        o_index_for_a2 <= 429;
        o_index_for_a3 <= 581;
        o_index_for_a4 <= 751;
        o_index_for_a5 <= 973; 
    end
    199: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 80;
        o_index_for_a1 <= 342;
        o_index_for_a2 <= 430;
        o_index_for_a3 <= 582;
        o_index_for_a4 <= 752;
        o_index_for_a5 <= 974; 
    end
    200: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 81;
        o_index_for_a1 <= 343;
        o_index_for_a2 <= 431;
        o_index_for_a3 <= 583;
        o_index_for_a4 <= 753;
        o_index_for_a5 <= 975; 
    end
    201: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 82;
        o_index_for_a1 <= 344;
        o_index_for_a2 <= 432;
        o_index_for_a3 <= 584;
        o_index_for_a4 <= 754;
        o_index_for_a5 <= 976; 
    end
    202: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 83;
        o_index_for_a1 <= 345;
        o_index_for_a2 <= 433;
        o_index_for_a3 <= 585;
        o_index_for_a4 <= 755;
        o_index_for_a5 <= 977; 
    end
    203: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 84;
        o_index_for_a1 <= 346;
        o_index_for_a2 <= 434;
        o_index_for_a3 <= 586;
        o_index_for_a4 <= 756;
        o_index_for_a5 <= 978; 
    end
    204: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 85;
        o_index_for_a1 <= 347;
        o_index_for_a2 <= 435;
        o_index_for_a3 <= 587;
        o_index_for_a4 <= 757;
        o_index_for_a5 <= 979; 
    end
    205: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 86;
        o_index_for_a1 <= 348;
        o_index_for_a2 <= 436;
        o_index_for_a3 <= 588;
        o_index_for_a4 <= 758;
        o_index_for_a5 <= 980; 
    end
    206: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 87;
        o_index_for_a1 <= 349;
        o_index_for_a2 <= 437;
        o_index_for_a3 <= 589;
        o_index_for_a4 <= 759;
        o_index_for_a5 <= 981; 
    end
    207: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 88;
        o_index_for_a1 <= 350;
        o_index_for_a2 <= 438;
        o_index_for_a3 <= 590;
        o_index_for_a4 <= 760;
        o_index_for_a5 <= 982; 
    end
    208: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 89;
        o_index_for_a1 <= 351;
        o_index_for_a2 <= 439;
        o_index_for_a3 <= 591;
        o_index_for_a4 <= 761;
        o_index_for_a5 <= 983; 
    end
    209: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 90;
        o_index_for_a1 <= 352;
        o_index_for_a2 <= 440;
        o_index_for_a3 <= 592;
        o_index_for_a4 <= 762;
        o_index_for_a5 <= 984; 
    end
    210: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 91;
        o_index_for_a1 <= 353;
        o_index_for_a2 <= 441;
        o_index_for_a3 <= 593;
        o_index_for_a4 <= 763;
        o_index_for_a5 <= 985; 
    end
    211: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 92;
        o_index_for_a1 <= 354;
        o_index_for_a2 <= 442;
        o_index_for_a3 <= 594;
        o_index_for_a4 <= 764;
        o_index_for_a5 <= 986; 
    end
    212: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 93;
        o_index_for_a1 <= 355;
        o_index_for_a2 <= 443;
        o_index_for_a3 <= 595;
        o_index_for_a4 <= 765;
        o_index_for_a5 <= 987; 
    end
    213: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 94;
        o_index_for_a1 <= 356;
        o_index_for_a2 <= 444;
        o_index_for_a3 <= 596;
        o_index_for_a4 <= 766;
        o_index_for_a5 <= 988; 
    end
    214: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 95;
        o_index_for_a1 <= 357;
        o_index_for_a2 <= 445;
        o_index_for_a3 <= 597;
        o_index_for_a4 <= 767;
        o_index_for_a5 <= 989; 
    end
    215: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 0;
        o_index_for_a1 <= 358;
        o_index_for_a2 <= 446;
        o_index_for_a3 <= 598;
        o_index_for_a4 <= 672;
        o_index_for_a5 <= 990; 
    end
    216: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 1;
        o_index_for_a1 <= 359;
        o_index_for_a2 <= 447;
        o_index_for_a3 <= 599;
        o_index_for_a4 <= 673;
        o_index_for_a5 <= 991; 
    end
    217: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 2;
        o_index_for_a1 <= 360;
        o_index_for_a2 <= 448;
        o_index_for_a3 <= 600;
        o_index_for_a4 <= 674;
        o_index_for_a5 <= 992; 
    end
    218: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 3;
        o_index_for_a1 <= 361;
        o_index_for_a2 <= 449;
        o_index_for_a3 <= 601;
        o_index_for_a4 <= 675;
        o_index_for_a5 <= 993; 
    end
    219: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 4;
        o_index_for_a1 <= 362;
        o_index_for_a2 <= 450;
        o_index_for_a3 <= 602;
        o_index_for_a4 <= 676;
        o_index_for_a5 <= 994; 
    end
    220: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 5;
        o_index_for_a1 <= 363;
        o_index_for_a2 <= 451;
        o_index_for_a3 <= 603;
        o_index_for_a4 <= 677;
        o_index_for_a5 <= 995; 
    end
    221: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 6;
        o_index_for_a1 <= 364;
        o_index_for_a2 <= 452;
        o_index_for_a3 <= 604;
        o_index_for_a4 <= 678;
        o_index_for_a5 <= 996; 
    end
    222: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 7;
        o_index_for_a1 <= 365;
        o_index_for_a2 <= 453;
        o_index_for_a3 <= 605;
        o_index_for_a4 <= 679;
        o_index_for_a5 <= 997; 
    end
    223: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 8;
        o_index_for_a1 <= 366;
        o_index_for_a2 <= 454;
        o_index_for_a3 <= 606;
        o_index_for_a4 <= 680;
        o_index_for_a5 <= 998; 
    end
    224: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 9;
        o_index_for_a1 <= 367;
        o_index_for_a2 <= 455;
        o_index_for_a3 <= 607;
        o_index_for_a4 <= 681;
        o_index_for_a5 <= 999; 
    end
    225: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 10;
        o_index_for_a1 <= 368;
        o_index_for_a2 <= 456;
        o_index_for_a3 <= 608;
        o_index_for_a4 <= 682;
        o_index_for_a5 <= 1000; 
    end
    226: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 11;
        o_index_for_a1 <= 369;
        o_index_for_a2 <= 457;
        o_index_for_a3 <= 609;
        o_index_for_a4 <= 683;
        o_index_for_a5 <= 1001; 
    end
    227: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 12;
        o_index_for_a1 <= 370;
        o_index_for_a2 <= 458;
        o_index_for_a3 <= 610;
        o_index_for_a4 <= 684;
        o_index_for_a5 <= 1002; 
    end
    228: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 13;
        o_index_for_a1 <= 371;
        o_index_for_a2 <= 459;
        o_index_for_a3 <= 611;
        o_index_for_a4 <= 685;
        o_index_for_a5 <= 1003; 
    end
    229: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 14;
        o_index_for_a1 <= 372;
        o_index_for_a2 <= 460;
        o_index_for_a3 <= 612;
        o_index_for_a4 <= 686;
        o_index_for_a5 <= 1004; 
    end
    230: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 15;
        o_index_for_a1 <= 373;
        o_index_for_a2 <= 461;
        o_index_for_a3 <= 613;
        o_index_for_a4 <= 687;
        o_index_for_a5 <= 1005; 
    end
    231: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 16;
        o_index_for_a1 <= 374;
        o_index_for_a2 <= 462;
        o_index_for_a3 <= 614;
        o_index_for_a4 <= 688;
        o_index_for_a5 <= 1006; 
    end
    232: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 17;
        o_index_for_a1 <= 375;
        o_index_for_a2 <= 463;
        o_index_for_a3 <= 615;
        o_index_for_a4 <= 689;
        o_index_for_a5 <= 1007; 
    end
    233: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 18;
        o_index_for_a1 <= 376;
        o_index_for_a2 <= 464;
        o_index_for_a3 <= 616;
        o_index_for_a4 <= 690;
        o_index_for_a5 <= 1008; 
    end
    234: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 19;
        o_index_for_a1 <= 377;
        o_index_for_a2 <= 465;
        o_index_for_a3 <= 617;
        o_index_for_a4 <= 691;
        o_index_for_a5 <= 1009; 
    end
    235: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 20;
        o_index_for_a1 <= 378;
        o_index_for_a2 <= 466;
        o_index_for_a3 <= 618;
        o_index_for_a4 <= 692;
        o_index_for_a5 <= 1010; 
    end
    236: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 21;
        o_index_for_a1 <= 379;
        o_index_for_a2 <= 467;
        o_index_for_a3 <= 619;
        o_index_for_a4 <= 693;
        o_index_for_a5 <= 1011; 
    end
    237: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 22;
        o_index_for_a1 <= 380;
        o_index_for_a2 <= 468;
        o_index_for_a3 <= 620;
        o_index_for_a4 <= 694;
        o_index_for_a5 <= 1012; 
    end
    238: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 23;
        o_index_for_a1 <= 381;
        o_index_for_a2 <= 469;
        o_index_for_a3 <= 621;
        o_index_for_a4 <= 695;
        o_index_for_a5 <= 1013; 
    end
    239: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 24;
        o_index_for_a1 <= 382;
        o_index_for_a2 <= 470;
        o_index_for_a3 <= 622;
        o_index_for_a4 <= 696;
        o_index_for_a5 <= 1014; 
    end
    240: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 25;
        o_index_for_a1 <= 383;
        o_index_for_a2 <= 471;
        o_index_for_a3 <= 623;
        o_index_for_a4 <= 697;
        o_index_for_a5 <= 1015; 
    end
    241: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 26;
        o_index_for_a1 <= 288;
        o_index_for_a2 <= 472;
        o_index_for_a3 <= 624;
        o_index_for_a4 <= 698;
        o_index_for_a5 <= 1016; 
    end
    242: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 27;
        o_index_for_a1 <= 289;
        o_index_for_a2 <= 473;
        o_index_for_a3 <= 625;
        o_index_for_a4 <= 699;
        o_index_for_a5 <= 1017; 
    end
    243: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 28;
        o_index_for_a1 <= 290;
        o_index_for_a2 <= 474;
        o_index_for_a3 <= 626;
        o_index_for_a4 <= 700;
        o_index_for_a5 <= 1018; 
    end
    244: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 29;
        o_index_for_a1 <= 291;
        o_index_for_a2 <= 475;
        o_index_for_a3 <= 627;
        o_index_for_a4 <= 701;
        o_index_for_a5 <= 1019; 
    end
    245: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 30;
        o_index_for_a1 <= 292;
        o_index_for_a2 <= 476;
        o_index_for_a3 <= 628;
        o_index_for_a4 <= 702;
        o_index_for_a5 <= 1020; 
    end
    246: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 31;
        o_index_for_a1 <= 293;
        o_index_for_a2 <= 477;
        o_index_for_a3 <= 629;
        o_index_for_a4 <= 703;
        o_index_for_a5 <= 1021; 
    end
    247: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 32;
        o_index_for_a1 <= 294;
        o_index_for_a2 <= 478;
        o_index_for_a3 <= 630;
        o_index_for_a4 <= 704;
        o_index_for_a5 <= 1022; 
    end
    248: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 33;
        o_index_for_a1 <= 295;
        o_index_for_a2 <= 479;
        o_index_for_a3 <= 631;
        o_index_for_a4 <= 705;
        o_index_for_a5 <= 1023; 
    end
    249: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 34;
        o_index_for_a1 <= 296;
        o_index_for_a2 <= 384;
        o_index_for_a3 <= 632;
        o_index_for_a4 <= 706;
        o_index_for_a5 <= 1024; 
    end
    250: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 35;
        o_index_for_a1 <= 297;
        o_index_for_a2 <= 385;
        o_index_for_a3 <= 633;
        o_index_for_a4 <= 707;
        o_index_for_a5 <= 1025; 
    end
    251: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 36;
        o_index_for_a1 <= 298;
        o_index_for_a2 <= 386;
        o_index_for_a3 <= 634;
        o_index_for_a4 <= 708;
        o_index_for_a5 <= 1026; 
    end
    252: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 37;
        o_index_for_a1 <= 299;
        o_index_for_a2 <= 387;
        o_index_for_a3 <= 635;
        o_index_for_a4 <= 709;
        o_index_for_a5 <= 1027; 
    end
    253: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 38;
        o_index_for_a1 <= 300;
        o_index_for_a2 <= 388;
        o_index_for_a3 <= 636;
        o_index_for_a4 <= 710;
        o_index_for_a5 <= 1028; 
    end
    254: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 39;
        o_index_for_a1 <= 301;
        o_index_for_a2 <= 389;
        o_index_for_a3 <= 637;
        o_index_for_a4 <= 711;
        o_index_for_a5 <= 1029; 
    end
    255: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 40;
        o_index_for_a1 <= 302;
        o_index_for_a2 <= 390;
        o_index_for_a3 <= 638;
        o_index_for_a4 <= 712;
        o_index_for_a5 <= 1030; 
    end
    256: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 41;
        o_index_for_a1 <= 303;
        o_index_for_a2 <= 391;
        o_index_for_a3 <= 639;
        o_index_for_a4 <= 713;
        o_index_for_a5 <= 1031; 
    end
    257: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 42;
        o_index_for_a1 <= 304;
        o_index_for_a2 <= 392;
        o_index_for_a3 <= 640;
        o_index_for_a4 <= 714;
        o_index_for_a5 <= 1032; 
    end
    258: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 43;
        o_index_for_a1 <= 305;
        o_index_for_a2 <= 393;
        o_index_for_a3 <= 641;
        o_index_for_a4 <= 715;
        o_index_for_a5 <= 1033; 
    end
    259: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 44;
        o_index_for_a1 <= 306;
        o_index_for_a2 <= 394;
        o_index_for_a3 <= 642;
        o_index_for_a4 <= 716;
        o_index_for_a5 <= 1034; 
    end
    260: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 45;
        o_index_for_a1 <= 307;
        o_index_for_a2 <= 395;
        o_index_for_a3 <= 643;
        o_index_for_a4 <= 717;
        o_index_for_a5 <= 1035; 
    end
    261: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 46;
        o_index_for_a1 <= 308;
        o_index_for_a2 <= 396;
        o_index_for_a3 <= 644;
        o_index_for_a4 <= 718;
        o_index_for_a5 <= 1036; 
    end
    262: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 47;
        o_index_for_a1 <= 309;
        o_index_for_a2 <= 397;
        o_index_for_a3 <= 645;
        o_index_for_a4 <= 719;
        o_index_for_a5 <= 1037; 
    end
    263: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 48;
        o_index_for_a1 <= 310;
        o_index_for_a2 <= 398;
        o_index_for_a3 <= 646;
        o_index_for_a4 <= 720;
        o_index_for_a5 <= 1038; 
    end
    264: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 49;
        o_index_for_a1 <= 311;
        o_index_for_a2 <= 399;
        o_index_for_a3 <= 647;
        o_index_for_a4 <= 721;
        o_index_for_a5 <= 1039; 
    end
    265: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 50;
        o_index_for_a1 <= 312;
        o_index_for_a2 <= 400;
        o_index_for_a3 <= 648;
        o_index_for_a4 <= 722;
        o_index_for_a5 <= 1040; 
    end
    266: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 51;
        o_index_for_a1 <= 313;
        o_index_for_a2 <= 401;
        o_index_for_a3 <= 649;
        o_index_for_a4 <= 723;
        o_index_for_a5 <= 1041; 
    end
    267: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 52;
        o_index_for_a1 <= 314;
        o_index_for_a2 <= 402;
        o_index_for_a3 <= 650;
        o_index_for_a4 <= 724;
        o_index_for_a5 <= 1042; 
    end
    268: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 53;
        o_index_for_a1 <= 315;
        o_index_for_a2 <= 403;
        o_index_for_a3 <= 651;
        o_index_for_a4 <= 725;
        o_index_for_a5 <= 1043; 
    end
    269: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 54;
        o_index_for_a1 <= 316;
        o_index_for_a2 <= 404;
        o_index_for_a3 <= 652;
        o_index_for_a4 <= 726;
        o_index_for_a5 <= 1044; 
    end
    270: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 55;
        o_index_for_a1 <= 317;
        o_index_for_a2 <= 405;
        o_index_for_a3 <= 653;
        o_index_for_a4 <= 727;
        o_index_for_a5 <= 1045; 
    end
    271: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 56;
        o_index_for_a1 <= 318;
        o_index_for_a2 <= 406;
        o_index_for_a3 <= 654;
        o_index_for_a4 <= 728;
        o_index_for_a5 <= 1046; 
    end
    272: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 57;
        o_index_for_a1 <= 319;
        o_index_for_a2 <= 407;
        o_index_for_a3 <= 655;
        o_index_for_a4 <= 729;
        o_index_for_a5 <= 1047; 
    end
    273: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 58;
        o_index_for_a1 <= 320;
        o_index_for_a2 <= 408;
        o_index_for_a3 <= 656;
        o_index_for_a4 <= 730;
        o_index_for_a5 <= 1048; 
    end
    274: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 59;
        o_index_for_a1 <= 321;
        o_index_for_a2 <= 409;
        o_index_for_a3 <= 657;
        o_index_for_a4 <= 731;
        o_index_for_a5 <= 1049; 
    end
    275: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 60;
        o_index_for_a1 <= 322;
        o_index_for_a2 <= 410;
        o_index_for_a3 <= 658;
        o_index_for_a4 <= 732;
        o_index_for_a5 <= 1050; 
    end
    276: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 61;
        o_index_for_a1 <= 323;
        o_index_for_a2 <= 411;
        o_index_for_a3 <= 659;
        o_index_for_a4 <= 733;
        o_index_for_a5 <= 1051; 
    end
    277: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 62;
        o_index_for_a1 <= 324;
        o_index_for_a2 <= 412;
        o_index_for_a3 <= 660;
        o_index_for_a4 <= 734;
        o_index_for_a5 <= 1052; 
    end
    278: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 63;
        o_index_for_a1 <= 325;
        o_index_for_a2 <= 413;
        o_index_for_a3 <= 661;
        o_index_for_a4 <= 735;
        o_index_for_a5 <= 1053; 
    end
    279: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 64;
        o_index_for_a1 <= 326;
        o_index_for_a2 <= 414;
        o_index_for_a3 <= 662;
        o_index_for_a4 <= 736;
        o_index_for_a5 <= 1054; 
    end
    280: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 65;
        o_index_for_a1 <= 327;
        o_index_for_a2 <= 415;
        o_index_for_a3 <= 663;
        o_index_for_a4 <= 737;
        o_index_for_a5 <= 1055; 
    end
    281: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 66;
        o_index_for_a1 <= 328;
        o_index_for_a2 <= 416;
        o_index_for_a3 <= 664;
        o_index_for_a4 <= 738;
        o_index_for_a5 <= 960; 
    end
    282: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 67;
        o_index_for_a1 <= 329;
        o_index_for_a2 <= 417;
        o_index_for_a3 <= 665;
        o_index_for_a4 <= 739;
        o_index_for_a5 <= 961; 
    end
    283: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 68;
        o_index_for_a1 <= 330;
        o_index_for_a2 <= 418;
        o_index_for_a3 <= 666;
        o_index_for_a4 <= 740;
        o_index_for_a5 <= 962; 
    end
    284: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 69;
        o_index_for_a1 <= 331;
        o_index_for_a2 <= 419;
        o_index_for_a3 <= 667;
        o_index_for_a4 <= 741;
        o_index_for_a5 <= 963; 
    end
    285: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 70;
        o_index_for_a1 <= 332;
        o_index_for_a2 <= 420;
        o_index_for_a3 <= 668;
        o_index_for_a4 <= 742;
        o_index_for_a5 <= 964; 
    end
    286: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 71;
        o_index_for_a1 <= 333;
        o_index_for_a2 <= 421;
        o_index_for_a3 <= 669;
        o_index_for_a4 <= 743;
        o_index_for_a5 <= 965; 
    end
    287: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_index_for_a0 <= 72;
        o_index_for_a1 <= 334;
        o_index_for_a2 <= 422;
        o_index_for_a3 <= 670;
        o_index_for_a4 <= 744;
        o_index_for_a5 <= 966; 
    end
    288: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 216;
        o_index_for_a1 <= 629;
        o_index_for_a2 <= 1025;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    289: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 217;
        o_index_for_a1 <= 630;
        o_index_for_a2 <= 1026;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    290: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 218;
        o_index_for_a1 <= 631;
        o_index_for_a2 <= 1027;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    291: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 219;
        o_index_for_a1 <= 632;
        o_index_for_a2 <= 1028;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    292: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 220;
        o_index_for_a1 <= 633;
        o_index_for_a2 <= 1029;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    293: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 221;
        o_index_for_a1 <= 634;
        o_index_for_a2 <= 1030;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    294: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 222;
        o_index_for_a1 <= 635;
        o_index_for_a2 <= 1031;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    295: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 223;
        o_index_for_a1 <= 636;
        o_index_for_a2 <= 1032;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    296: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 224;
        o_index_for_a1 <= 637;
        o_index_for_a2 <= 1033;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    297: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 225;
        o_index_for_a1 <= 638;
        o_index_for_a2 <= 1034;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    298: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 226;
        o_index_for_a1 <= 639;
        o_index_for_a2 <= 1035;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    299: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 227;
        o_index_for_a1 <= 640;
        o_index_for_a2 <= 1036;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    300: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 228;
        o_index_for_a1 <= 641;
        o_index_for_a2 <= 1037;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    301: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 229;
        o_index_for_a1 <= 642;
        o_index_for_a2 <= 1038;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    302: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 230;
        o_index_for_a1 <= 643;
        o_index_for_a2 <= 1039;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    303: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 231;
        o_index_for_a1 <= 644;
        o_index_for_a2 <= 1040;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    304: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 232;
        o_index_for_a1 <= 645;
        o_index_for_a2 <= 1041;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    305: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 233;
        o_index_for_a1 <= 646;
        o_index_for_a2 <= 1042;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    306: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 234;
        o_index_for_a1 <= 647;
        o_index_for_a2 <= 1043;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    307: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 235;
        o_index_for_a1 <= 648;
        o_index_for_a2 <= 1044;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    308: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 236;
        o_index_for_a1 <= 649;
        o_index_for_a2 <= 1045;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    309: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 237;
        o_index_for_a1 <= 650;
        o_index_for_a2 <= 1046;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    310: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 238;
        o_index_for_a1 <= 651;
        o_index_for_a2 <= 1047;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    311: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 239;
        o_index_for_a1 <= 652;
        o_index_for_a2 <= 1048;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    312: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 240;
        o_index_for_a1 <= 653;
        o_index_for_a2 <= 1049;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    313: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 241;
        o_index_for_a1 <= 654;
        o_index_for_a2 <= 1050;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    314: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 242;
        o_index_for_a1 <= 655;
        o_index_for_a2 <= 1051;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    315: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 243;
        o_index_for_a1 <= 656;
        o_index_for_a2 <= 1052;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    316: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 244;
        o_index_for_a1 <= 657;
        o_index_for_a2 <= 1053;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    317: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 245;
        o_index_for_a1 <= 658;
        o_index_for_a2 <= 1054;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    318: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 246;
        o_index_for_a1 <= 659;
        o_index_for_a2 <= 1055;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    319: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 247;
        o_index_for_a1 <= 660;
        o_index_for_a2 <= 960;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    320: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 248;
        o_index_for_a1 <= 661;
        o_index_for_a2 <= 961;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    321: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 249;
        o_index_for_a1 <= 662;
        o_index_for_a2 <= 962;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    322: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 250;
        o_index_for_a1 <= 663;
        o_index_for_a2 <= 963;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    323: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 251;
        o_index_for_a1 <= 664;
        o_index_for_a2 <= 964;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    324: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 252;
        o_index_for_a1 <= 665;
        o_index_for_a2 <= 965;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    325: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 253;
        o_index_for_a1 <= 666;
        o_index_for_a2 <= 966;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    326: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 254;
        o_index_for_a1 <= 667;
        o_index_for_a2 <= 967;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    327: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 255;
        o_index_for_a1 <= 668;
        o_index_for_a2 <= 968;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    328: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 256;
        o_index_for_a1 <= 669;
        o_index_for_a2 <= 969;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    329: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 257;
        o_index_for_a1 <= 670;
        o_index_for_a2 <= 970;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    330: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 258;
        o_index_for_a1 <= 671;
        o_index_for_a2 <= 971;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    331: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 259;
        o_index_for_a1 <= 576;
        o_index_for_a2 <= 972;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    332: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 260;
        o_index_for_a1 <= 577;
        o_index_for_a2 <= 973;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    333: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 261;
        o_index_for_a1 <= 578;
        o_index_for_a2 <= 974;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    334: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 262;
        o_index_for_a1 <= 579;
        o_index_for_a2 <= 975;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    335: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 263;
        o_index_for_a1 <= 580;
        o_index_for_a2 <= 976;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    336: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 264;
        o_index_for_a1 <= 581;
        o_index_for_a2 <= 977;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    337: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 265;
        o_index_for_a1 <= 582;
        o_index_for_a2 <= 978;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    338: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 266;
        o_index_for_a1 <= 583;
        o_index_for_a2 <= 979;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    339: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 267;
        o_index_for_a1 <= 584;
        o_index_for_a2 <= 980;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    340: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 268;
        o_index_for_a1 <= 585;
        o_index_for_a2 <= 981;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    341: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 269;
        o_index_for_a1 <= 586;
        o_index_for_a2 <= 982;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    342: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 270;
        o_index_for_a1 <= 587;
        o_index_for_a2 <= 983;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    343: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 271;
        o_index_for_a1 <= 588;
        o_index_for_a2 <= 984;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    344: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 272;
        o_index_for_a1 <= 589;
        o_index_for_a2 <= 985;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    345: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 273;
        o_index_for_a1 <= 590;
        o_index_for_a2 <= 986;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    346: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 274;
        o_index_for_a1 <= 591;
        o_index_for_a2 <= 987;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    347: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 275;
        o_index_for_a1 <= 592;
        o_index_for_a2 <= 988;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    348: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 276;
        o_index_for_a1 <= 593;
        o_index_for_a2 <= 989;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    349: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 277;
        o_index_for_a1 <= 594;
        o_index_for_a2 <= 990;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    350: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 278;
        o_index_for_a1 <= 595;
        o_index_for_a2 <= 991;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    351: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 279;
        o_index_for_a1 <= 596;
        o_index_for_a2 <= 992;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    352: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 280;
        o_index_for_a1 <= 597;
        o_index_for_a2 <= 993;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    353: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 281;
        o_index_for_a1 <= 598;
        o_index_for_a2 <= 994;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    354: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 282;
        o_index_for_a1 <= 599;
        o_index_for_a2 <= 995;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    355: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 283;
        o_index_for_a1 <= 600;
        o_index_for_a2 <= 996;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    356: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 284;
        o_index_for_a1 <= 601;
        o_index_for_a2 <= 997;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    357: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 285;
        o_index_for_a1 <= 602;
        o_index_for_a2 <= 998;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    358: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 286;
        o_index_for_a1 <= 603;
        o_index_for_a2 <= 999;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    359: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 287;
        o_index_for_a1 <= 604;
        o_index_for_a2 <= 1000;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    360: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 192;
        o_index_for_a1 <= 605;
        o_index_for_a2 <= 1001;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    361: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 193;
        o_index_for_a1 <= 606;
        o_index_for_a2 <= 1002;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    362: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 194;
        o_index_for_a1 <= 607;
        o_index_for_a2 <= 1003;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    363: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 195;
        o_index_for_a1 <= 608;
        o_index_for_a2 <= 1004;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    364: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 196;
        o_index_for_a1 <= 609;
        o_index_for_a2 <= 1005;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    365: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 197;
        o_index_for_a1 <= 610;
        o_index_for_a2 <= 1006;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    366: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 198;
        o_index_for_a1 <= 611;
        o_index_for_a2 <= 1007;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    367: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 199;
        o_index_for_a1 <= 612;
        o_index_for_a2 <= 1008;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    368: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 200;
        o_index_for_a1 <= 613;
        o_index_for_a2 <= 1009;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    369: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 201;
        o_index_for_a1 <= 614;
        o_index_for_a2 <= 1010;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    370: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 202;
        o_index_for_a1 <= 615;
        o_index_for_a2 <= 1011;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    371: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 203;
        o_index_for_a1 <= 616;
        o_index_for_a2 <= 1012;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    372: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 204;
        o_index_for_a1 <= 617;
        o_index_for_a2 <= 1013;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    373: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 205;
        o_index_for_a1 <= 618;
        o_index_for_a2 <= 1014;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    374: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 206;
        o_index_for_a1 <= 619;
        o_index_for_a2 <= 1015;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    375: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 207;
        o_index_for_a1 <= 620;
        o_index_for_a2 <= 1016;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    376: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 208;
        o_index_for_a1 <= 621;
        o_index_for_a2 <= 1017;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    377: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 209;
        o_index_for_a1 <= 622;
        o_index_for_a2 <= 1018;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    378: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 210;
        o_index_for_a1 <= 623;
        o_index_for_a2 <= 1019;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    379: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 211;
        o_index_for_a1 <= 624;
        o_index_for_a2 <= 1020;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    380: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 212;
        o_index_for_a1 <= 625;
        o_index_for_a2 <= 1021;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    381: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 213;
        o_index_for_a1 <= 626;
        o_index_for_a2 <= 1022;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    382: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 214;
        o_index_for_a1 <= 627;
        o_index_for_a2 <= 1023;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    383: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 215;
        o_index_for_a1 <= 628;
        o_index_for_a2 <= 1024;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    384: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 214;
        o_index_for_a1 <= 526;
        o_index_for_a2 <= 851;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    385: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 215;
        o_index_for_a1 <= 527;
        o_index_for_a2 <= 852;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    386: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 216;
        o_index_for_a1 <= 528;
        o_index_for_a2 <= 853;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    387: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 217;
        o_index_for_a1 <= 529;
        o_index_for_a2 <= 854;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    388: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 218;
        o_index_for_a1 <= 530;
        o_index_for_a2 <= 855;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    389: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 219;
        o_index_for_a1 <= 531;
        o_index_for_a2 <= 856;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    390: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 220;
        o_index_for_a1 <= 532;
        o_index_for_a2 <= 857;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    391: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 221;
        o_index_for_a1 <= 533;
        o_index_for_a2 <= 858;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    392: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 222;
        o_index_for_a1 <= 534;
        o_index_for_a2 <= 859;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    393: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 223;
        o_index_for_a1 <= 535;
        o_index_for_a2 <= 860;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    394: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 224;
        o_index_for_a1 <= 536;
        o_index_for_a2 <= 861;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    395: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 225;
        o_index_for_a1 <= 537;
        o_index_for_a2 <= 862;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    396: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 226;
        o_index_for_a1 <= 538;
        o_index_for_a2 <= 863;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    397: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 227;
        o_index_for_a1 <= 539;
        o_index_for_a2 <= 768;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    398: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 228;
        o_index_for_a1 <= 540;
        o_index_for_a2 <= 769;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    399: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 229;
        o_index_for_a1 <= 541;
        o_index_for_a2 <= 770;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    400: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 230;
        o_index_for_a1 <= 542;
        o_index_for_a2 <= 771;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    401: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 231;
        o_index_for_a1 <= 543;
        o_index_for_a2 <= 772;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    402: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 232;
        o_index_for_a1 <= 544;
        o_index_for_a2 <= 773;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    403: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 233;
        o_index_for_a1 <= 545;
        o_index_for_a2 <= 774;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    404: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 234;
        o_index_for_a1 <= 546;
        o_index_for_a2 <= 775;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    405: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 235;
        o_index_for_a1 <= 547;
        o_index_for_a2 <= 776;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    406: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 236;
        o_index_for_a1 <= 548;
        o_index_for_a2 <= 777;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    407: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 237;
        o_index_for_a1 <= 549;
        o_index_for_a2 <= 778;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    408: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 238;
        o_index_for_a1 <= 550;
        o_index_for_a2 <= 779;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    409: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 239;
        o_index_for_a1 <= 551;
        o_index_for_a2 <= 780;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    410: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 240;
        o_index_for_a1 <= 552;
        o_index_for_a2 <= 781;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    411: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 241;
        o_index_for_a1 <= 553;
        o_index_for_a2 <= 782;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    412: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 242;
        o_index_for_a1 <= 554;
        o_index_for_a2 <= 783;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    413: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 243;
        o_index_for_a1 <= 555;
        o_index_for_a2 <= 784;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    414: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 244;
        o_index_for_a1 <= 556;
        o_index_for_a2 <= 785;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    415: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 245;
        o_index_for_a1 <= 557;
        o_index_for_a2 <= 786;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    416: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 246;
        o_index_for_a1 <= 558;
        o_index_for_a2 <= 787;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    417: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 247;
        o_index_for_a1 <= 559;
        o_index_for_a2 <= 788;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    418: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 248;
        o_index_for_a1 <= 560;
        o_index_for_a2 <= 789;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    419: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 249;
        o_index_for_a1 <= 561;
        o_index_for_a2 <= 790;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    420: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 250;
        o_index_for_a1 <= 562;
        o_index_for_a2 <= 791;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    421: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 251;
        o_index_for_a1 <= 563;
        o_index_for_a2 <= 792;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    422: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 252;
        o_index_for_a1 <= 564;
        o_index_for_a2 <= 793;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    423: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 253;
        o_index_for_a1 <= 565;
        o_index_for_a2 <= 794;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    424: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 254;
        o_index_for_a1 <= 566;
        o_index_for_a2 <= 795;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    425: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 255;
        o_index_for_a1 <= 567;
        o_index_for_a2 <= 796;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    426: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 256;
        o_index_for_a1 <= 568;
        o_index_for_a2 <= 797;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    427: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 257;
        o_index_for_a1 <= 569;
        o_index_for_a2 <= 798;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    428: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 258;
        o_index_for_a1 <= 570;
        o_index_for_a2 <= 799;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    429: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 259;
        o_index_for_a1 <= 571;
        o_index_for_a2 <= 800;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    430: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 260;
        o_index_for_a1 <= 572;
        o_index_for_a2 <= 801;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    431: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 261;
        o_index_for_a1 <= 573;
        o_index_for_a2 <= 802;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    432: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 262;
        o_index_for_a1 <= 574;
        o_index_for_a2 <= 803;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    433: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 263;
        o_index_for_a1 <= 575;
        o_index_for_a2 <= 804;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    434: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 264;
        o_index_for_a1 <= 480;
        o_index_for_a2 <= 805;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    435: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 265;
        o_index_for_a1 <= 481;
        o_index_for_a2 <= 806;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    436: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 266;
        o_index_for_a1 <= 482;
        o_index_for_a2 <= 807;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    437: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 267;
        o_index_for_a1 <= 483;
        o_index_for_a2 <= 808;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    438: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 268;
        o_index_for_a1 <= 484;
        o_index_for_a2 <= 809;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    439: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 269;
        o_index_for_a1 <= 485;
        o_index_for_a2 <= 810;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    440: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 270;
        o_index_for_a1 <= 486;
        o_index_for_a2 <= 811;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    441: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 271;
        o_index_for_a1 <= 487;
        o_index_for_a2 <= 812;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    442: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 272;
        o_index_for_a1 <= 488;
        o_index_for_a2 <= 813;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    443: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 273;
        o_index_for_a1 <= 489;
        o_index_for_a2 <= 814;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    444: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 274;
        o_index_for_a1 <= 490;
        o_index_for_a2 <= 815;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    445: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 275;
        o_index_for_a1 <= 491;
        o_index_for_a2 <= 816;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    446: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 276;
        o_index_for_a1 <= 492;
        o_index_for_a2 <= 817;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    447: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 277;
        o_index_for_a1 <= 493;
        o_index_for_a2 <= 818;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    448: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 278;
        o_index_for_a1 <= 494;
        o_index_for_a2 <= 819;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    449: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 279;
        o_index_for_a1 <= 495;
        o_index_for_a2 <= 820;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    450: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 280;
        o_index_for_a1 <= 496;
        o_index_for_a2 <= 821;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    451: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 281;
        o_index_for_a1 <= 497;
        o_index_for_a2 <= 822;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    452: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 282;
        o_index_for_a1 <= 498;
        o_index_for_a2 <= 823;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    453: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 283;
        o_index_for_a1 <= 499;
        o_index_for_a2 <= 824;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    454: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 284;
        o_index_for_a1 <= 500;
        o_index_for_a2 <= 825;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    455: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 285;
        o_index_for_a1 <= 501;
        o_index_for_a2 <= 826;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    456: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 286;
        o_index_for_a1 <= 502;
        o_index_for_a2 <= 827;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    457: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 287;
        o_index_for_a1 <= 503;
        o_index_for_a2 <= 828;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    458: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 192;
        o_index_for_a1 <= 504;
        o_index_for_a2 <= 829;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    459: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 193;
        o_index_for_a1 <= 505;
        o_index_for_a2 <= 830;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    460: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 194;
        o_index_for_a1 <= 506;
        o_index_for_a2 <= 831;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    461: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 195;
        o_index_for_a1 <= 507;
        o_index_for_a2 <= 832;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    462: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 196;
        o_index_for_a1 <= 508;
        o_index_for_a2 <= 833;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    463: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 197;
        o_index_for_a1 <= 509;
        o_index_for_a2 <= 834;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    464: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 198;
        o_index_for_a1 <= 510;
        o_index_for_a2 <= 835;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    465: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 199;
        o_index_for_a1 <= 511;
        o_index_for_a2 <= 836;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    466: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 200;
        o_index_for_a1 <= 512;
        o_index_for_a2 <= 837;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    467: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 201;
        o_index_for_a1 <= 513;
        o_index_for_a2 <= 838;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    468: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 202;
        o_index_for_a1 <= 514;
        o_index_for_a2 <= 839;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    469: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 203;
        o_index_for_a1 <= 515;
        o_index_for_a2 <= 840;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    470: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 204;
        o_index_for_a1 <= 516;
        o_index_for_a2 <= 841;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    471: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 205;
        o_index_for_a1 <= 517;
        o_index_for_a2 <= 842;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    472: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 206;
        o_index_for_a1 <= 518;
        o_index_for_a2 <= 843;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    473: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 207;
        o_index_for_a1 <= 519;
        o_index_for_a2 <= 844;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    474: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 208;
        o_index_for_a1 <= 520;
        o_index_for_a2 <= 845;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    475: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 209;
        o_index_for_a1 <= 521;
        o_index_for_a2 <= 846;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    476: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 210;
        o_index_for_a1 <= 522;
        o_index_for_a2 <= 847;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    477: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 211;
        o_index_for_a1 <= 523;
        o_index_for_a2 <= 848;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    478: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 212;
        o_index_for_a1 <= 524;
        o_index_for_a2 <= 849;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    479: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 213;
        o_index_for_a1 <= 525;
        o_index_for_a2 <= 850;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    480: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 118;
        o_index_for_a1 <= 273;
        o_index_for_a2 <= 520;
        o_index_for_a3 <= 792;
        o_index_for_a4 <= 958;
        o_index_for_a5 <= 1122; 
    end
    481: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 119;
        o_index_for_a1 <= 274;
        o_index_for_a2 <= 521;
        o_index_for_a3 <= 793;
        o_index_for_a4 <= 959;
        o_index_for_a5 <= 1123; 
    end
    482: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 120;
        o_index_for_a1 <= 275;
        o_index_for_a2 <= 522;
        o_index_for_a3 <= 794;
        o_index_for_a4 <= 864;
        o_index_for_a5 <= 1124; 
    end
    483: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 121;
        o_index_for_a1 <= 276;
        o_index_for_a2 <= 523;
        o_index_for_a3 <= 795;
        o_index_for_a4 <= 865;
        o_index_for_a5 <= 1125; 
    end
    484: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 122;
        o_index_for_a1 <= 277;
        o_index_for_a2 <= 524;
        o_index_for_a3 <= 796;
        o_index_for_a4 <= 866;
        o_index_for_a5 <= 1126; 
    end
    485: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 123;
        o_index_for_a1 <= 278;
        o_index_for_a2 <= 525;
        o_index_for_a3 <= 797;
        o_index_for_a4 <= 867;
        o_index_for_a5 <= 1127; 
    end
    486: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 124;
        o_index_for_a1 <= 279;
        o_index_for_a2 <= 526;
        o_index_for_a3 <= 798;
        o_index_for_a4 <= 868;
        o_index_for_a5 <= 1128; 
    end
    487: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 125;
        o_index_for_a1 <= 280;
        o_index_for_a2 <= 527;
        o_index_for_a3 <= 799;
        o_index_for_a4 <= 869;
        o_index_for_a5 <= 1129; 
    end
    488: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 126;
        o_index_for_a1 <= 281;
        o_index_for_a2 <= 528;
        o_index_for_a3 <= 800;
        o_index_for_a4 <= 870;
        o_index_for_a5 <= 1130; 
    end
    489: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 127;
        o_index_for_a1 <= 282;
        o_index_for_a2 <= 529;
        o_index_for_a3 <= 801;
        o_index_for_a4 <= 871;
        o_index_for_a5 <= 1131; 
    end
    490: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 128;
        o_index_for_a1 <= 283;
        o_index_for_a2 <= 530;
        o_index_for_a3 <= 802;
        o_index_for_a4 <= 872;
        o_index_for_a5 <= 1132; 
    end
    491: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 129;
        o_index_for_a1 <= 284;
        o_index_for_a2 <= 531;
        o_index_for_a3 <= 803;
        o_index_for_a4 <= 873;
        o_index_for_a5 <= 1133; 
    end
    492: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 130;
        o_index_for_a1 <= 285;
        o_index_for_a2 <= 532;
        o_index_for_a3 <= 804;
        o_index_for_a4 <= 874;
        o_index_for_a5 <= 1134; 
    end
    493: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 131;
        o_index_for_a1 <= 286;
        o_index_for_a2 <= 533;
        o_index_for_a3 <= 805;
        o_index_for_a4 <= 875;
        o_index_for_a5 <= 1135; 
    end
    494: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 132;
        o_index_for_a1 <= 287;
        o_index_for_a2 <= 534;
        o_index_for_a3 <= 806;
        o_index_for_a4 <= 876;
        o_index_for_a5 <= 1136; 
    end
    495: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 133;
        o_index_for_a1 <= 192;
        o_index_for_a2 <= 535;
        o_index_for_a3 <= 807;
        o_index_for_a4 <= 877;
        o_index_for_a5 <= 1137; 
    end
    496: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 134;
        o_index_for_a1 <= 193;
        o_index_for_a2 <= 536;
        o_index_for_a3 <= 808;
        o_index_for_a4 <= 878;
        o_index_for_a5 <= 1138; 
    end
    497: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 135;
        o_index_for_a1 <= 194;
        o_index_for_a2 <= 537;
        o_index_for_a3 <= 809;
        o_index_for_a4 <= 879;
        o_index_for_a5 <= 1139; 
    end
    498: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 136;
        o_index_for_a1 <= 195;
        o_index_for_a2 <= 538;
        o_index_for_a3 <= 810;
        o_index_for_a4 <= 880;
        o_index_for_a5 <= 1140; 
    end
    499: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 137;
        o_index_for_a1 <= 196;
        o_index_for_a2 <= 539;
        o_index_for_a3 <= 811;
        o_index_for_a4 <= 881;
        o_index_for_a5 <= 1141; 
    end
    500: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 138;
        o_index_for_a1 <= 197;
        o_index_for_a2 <= 540;
        o_index_for_a3 <= 812;
        o_index_for_a4 <= 882;
        o_index_for_a5 <= 1142; 
    end
    501: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 139;
        o_index_for_a1 <= 198;
        o_index_for_a2 <= 541;
        o_index_for_a3 <= 813;
        o_index_for_a4 <= 883;
        o_index_for_a5 <= 1143; 
    end
    502: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 140;
        o_index_for_a1 <= 199;
        o_index_for_a2 <= 542;
        o_index_for_a3 <= 814;
        o_index_for_a4 <= 884;
        o_index_for_a5 <= 1144; 
    end
    503: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 141;
        o_index_for_a1 <= 200;
        o_index_for_a2 <= 543;
        o_index_for_a3 <= 815;
        o_index_for_a4 <= 885;
        o_index_for_a5 <= 1145; 
    end
    504: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 142;
        o_index_for_a1 <= 201;
        o_index_for_a2 <= 544;
        o_index_for_a3 <= 816;
        o_index_for_a4 <= 886;
        o_index_for_a5 <= 1146; 
    end
    505: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 143;
        o_index_for_a1 <= 202;
        o_index_for_a2 <= 545;
        o_index_for_a3 <= 817;
        o_index_for_a4 <= 887;
        o_index_for_a5 <= 1147; 
    end
    506: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 144;
        o_index_for_a1 <= 203;
        o_index_for_a2 <= 546;
        o_index_for_a3 <= 818;
        o_index_for_a4 <= 888;
        o_index_for_a5 <= 1148; 
    end
    507: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 145;
        o_index_for_a1 <= 204;
        o_index_for_a2 <= 547;
        o_index_for_a3 <= 819;
        o_index_for_a4 <= 889;
        o_index_for_a5 <= 1149; 
    end
    508: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 146;
        o_index_for_a1 <= 205;
        o_index_for_a2 <= 548;
        o_index_for_a3 <= 820;
        o_index_for_a4 <= 890;
        o_index_for_a5 <= 1150; 
    end
    509: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 147;
        o_index_for_a1 <= 206;
        o_index_for_a2 <= 549;
        o_index_for_a3 <= 821;
        o_index_for_a4 <= 891;
        o_index_for_a5 <= 1151; 
    end
    510: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 148;
        o_index_for_a1 <= 207;
        o_index_for_a2 <= 550;
        o_index_for_a3 <= 822;
        o_index_for_a4 <= 892;
        o_index_for_a5 <= 1056; 
    end
    511: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 149;
        o_index_for_a1 <= 208;
        o_index_for_a2 <= 551;
        o_index_for_a3 <= 823;
        o_index_for_a4 <= 893;
        o_index_for_a5 <= 1057; 
    end
    512: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 150;
        o_index_for_a1 <= 209;
        o_index_for_a2 <= 552;
        o_index_for_a3 <= 824;
        o_index_for_a4 <= 894;
        o_index_for_a5 <= 1058; 
    end
    513: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 151;
        o_index_for_a1 <= 210;
        o_index_for_a2 <= 553;
        o_index_for_a3 <= 825;
        o_index_for_a4 <= 895;
        o_index_for_a5 <= 1059; 
    end
    514: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 152;
        o_index_for_a1 <= 211;
        o_index_for_a2 <= 554;
        o_index_for_a3 <= 826;
        o_index_for_a4 <= 896;
        o_index_for_a5 <= 1060; 
    end
    515: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 153;
        o_index_for_a1 <= 212;
        o_index_for_a2 <= 555;
        o_index_for_a3 <= 827;
        o_index_for_a4 <= 897;
        o_index_for_a5 <= 1061; 
    end
    516: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 154;
        o_index_for_a1 <= 213;
        o_index_for_a2 <= 556;
        o_index_for_a3 <= 828;
        o_index_for_a4 <= 898;
        o_index_for_a5 <= 1062; 
    end
    517: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 155;
        o_index_for_a1 <= 214;
        o_index_for_a2 <= 557;
        o_index_for_a3 <= 829;
        o_index_for_a4 <= 899;
        o_index_for_a5 <= 1063; 
    end
    518: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 156;
        o_index_for_a1 <= 215;
        o_index_for_a2 <= 558;
        o_index_for_a3 <= 830;
        o_index_for_a4 <= 900;
        o_index_for_a5 <= 1064; 
    end
    519: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 157;
        o_index_for_a1 <= 216;
        o_index_for_a2 <= 559;
        o_index_for_a3 <= 831;
        o_index_for_a4 <= 901;
        o_index_for_a5 <= 1065; 
    end
    520: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 158;
        o_index_for_a1 <= 217;
        o_index_for_a2 <= 560;
        o_index_for_a3 <= 832;
        o_index_for_a4 <= 902;
        o_index_for_a5 <= 1066; 
    end
    521: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 159;
        o_index_for_a1 <= 218;
        o_index_for_a2 <= 561;
        o_index_for_a3 <= 833;
        o_index_for_a4 <= 903;
        o_index_for_a5 <= 1067; 
    end
    522: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 160;
        o_index_for_a1 <= 219;
        o_index_for_a2 <= 562;
        o_index_for_a3 <= 834;
        o_index_for_a4 <= 904;
        o_index_for_a5 <= 1068; 
    end
    523: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 161;
        o_index_for_a1 <= 220;
        o_index_for_a2 <= 563;
        o_index_for_a3 <= 835;
        o_index_for_a4 <= 905;
        o_index_for_a5 <= 1069; 
    end
    524: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 162;
        o_index_for_a1 <= 221;
        o_index_for_a2 <= 564;
        o_index_for_a3 <= 836;
        o_index_for_a4 <= 906;
        o_index_for_a5 <= 1070; 
    end
    525: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 163;
        o_index_for_a1 <= 222;
        o_index_for_a2 <= 565;
        o_index_for_a3 <= 837;
        o_index_for_a4 <= 907;
        o_index_for_a5 <= 1071; 
    end
    526: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 164;
        o_index_for_a1 <= 223;
        o_index_for_a2 <= 566;
        o_index_for_a3 <= 838;
        o_index_for_a4 <= 908;
        o_index_for_a5 <= 1072; 
    end
    527: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 165;
        o_index_for_a1 <= 224;
        o_index_for_a2 <= 567;
        o_index_for_a3 <= 839;
        o_index_for_a4 <= 909;
        o_index_for_a5 <= 1073; 
    end
    528: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 166;
        o_index_for_a1 <= 225;
        o_index_for_a2 <= 568;
        o_index_for_a3 <= 840;
        o_index_for_a4 <= 910;
        o_index_for_a5 <= 1074; 
    end
    529: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 167;
        o_index_for_a1 <= 226;
        o_index_for_a2 <= 569;
        o_index_for_a3 <= 841;
        o_index_for_a4 <= 911;
        o_index_for_a5 <= 1075; 
    end
    530: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 168;
        o_index_for_a1 <= 227;
        o_index_for_a2 <= 570;
        o_index_for_a3 <= 842;
        o_index_for_a4 <= 912;
        o_index_for_a5 <= 1076; 
    end
    531: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 169;
        o_index_for_a1 <= 228;
        o_index_for_a2 <= 571;
        o_index_for_a3 <= 843;
        o_index_for_a4 <= 913;
        o_index_for_a5 <= 1077; 
    end
    532: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 170;
        o_index_for_a1 <= 229;
        o_index_for_a2 <= 572;
        o_index_for_a3 <= 844;
        o_index_for_a4 <= 914;
        o_index_for_a5 <= 1078; 
    end
    533: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 171;
        o_index_for_a1 <= 230;
        o_index_for_a2 <= 573;
        o_index_for_a3 <= 845;
        o_index_for_a4 <= 915;
        o_index_for_a5 <= 1079; 
    end
    534: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 172;
        o_index_for_a1 <= 231;
        o_index_for_a2 <= 574;
        o_index_for_a3 <= 846;
        o_index_for_a4 <= 916;
        o_index_for_a5 <= 1080; 
    end
    535: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 173;
        o_index_for_a1 <= 232;
        o_index_for_a2 <= 575;
        o_index_for_a3 <= 847;
        o_index_for_a4 <= 917;
        o_index_for_a5 <= 1081; 
    end
    536: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 174;
        o_index_for_a1 <= 233;
        o_index_for_a2 <= 480;
        o_index_for_a3 <= 848;
        o_index_for_a4 <= 918;
        o_index_for_a5 <= 1082; 
    end
    537: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 175;
        o_index_for_a1 <= 234;
        o_index_for_a2 <= 481;
        o_index_for_a3 <= 849;
        o_index_for_a4 <= 919;
        o_index_for_a5 <= 1083; 
    end
    538: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 176;
        o_index_for_a1 <= 235;
        o_index_for_a2 <= 482;
        o_index_for_a3 <= 850;
        o_index_for_a4 <= 920;
        o_index_for_a5 <= 1084; 
    end
    539: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 177;
        o_index_for_a1 <= 236;
        o_index_for_a2 <= 483;
        o_index_for_a3 <= 851;
        o_index_for_a4 <= 921;
        o_index_for_a5 <= 1085; 
    end
    540: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 178;
        o_index_for_a1 <= 237;
        o_index_for_a2 <= 484;
        o_index_for_a3 <= 852;
        o_index_for_a4 <= 922;
        o_index_for_a5 <= 1086; 
    end
    541: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 179;
        o_index_for_a1 <= 238;
        o_index_for_a2 <= 485;
        o_index_for_a3 <= 853;
        o_index_for_a4 <= 923;
        o_index_for_a5 <= 1087; 
    end
    542: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 180;
        o_index_for_a1 <= 239;
        o_index_for_a2 <= 486;
        o_index_for_a3 <= 854;
        o_index_for_a4 <= 924;
        o_index_for_a5 <= 1088; 
    end
    543: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 181;
        o_index_for_a1 <= 240;
        o_index_for_a2 <= 487;
        o_index_for_a3 <= 855;
        o_index_for_a4 <= 925;
        o_index_for_a5 <= 1089; 
    end
    544: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 182;
        o_index_for_a1 <= 241;
        o_index_for_a2 <= 488;
        o_index_for_a3 <= 856;
        o_index_for_a4 <= 926;
        o_index_for_a5 <= 1090; 
    end
    545: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 183;
        o_index_for_a1 <= 242;
        o_index_for_a2 <= 489;
        o_index_for_a3 <= 857;
        o_index_for_a4 <= 927;
        o_index_for_a5 <= 1091; 
    end
    546: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 184;
        o_index_for_a1 <= 243;
        o_index_for_a2 <= 490;
        o_index_for_a3 <= 858;
        o_index_for_a4 <= 928;
        o_index_for_a5 <= 1092; 
    end
    547: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 185;
        o_index_for_a1 <= 244;
        o_index_for_a2 <= 491;
        o_index_for_a3 <= 859;
        o_index_for_a4 <= 929;
        o_index_for_a5 <= 1093; 
    end
    548: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 186;
        o_index_for_a1 <= 245;
        o_index_for_a2 <= 492;
        o_index_for_a3 <= 860;
        o_index_for_a4 <= 930;
        o_index_for_a5 <= 1094; 
    end
    549: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 187;
        o_index_for_a1 <= 246;
        o_index_for_a2 <= 493;
        o_index_for_a3 <= 861;
        o_index_for_a4 <= 931;
        o_index_for_a5 <= 1095; 
    end
    550: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 188;
        o_index_for_a1 <= 247;
        o_index_for_a2 <= 494;
        o_index_for_a3 <= 862;
        o_index_for_a4 <= 932;
        o_index_for_a5 <= 1096; 
    end
    551: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 189;
        o_index_for_a1 <= 248;
        o_index_for_a2 <= 495;
        o_index_for_a3 <= 863;
        o_index_for_a4 <= 933;
        o_index_for_a5 <= 1097; 
    end
    552: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 190;
        o_index_for_a1 <= 249;
        o_index_for_a2 <= 496;
        o_index_for_a3 <= 768;
        o_index_for_a4 <= 934;
        o_index_for_a5 <= 1098; 
    end
    553: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 191;
        o_index_for_a1 <= 250;
        o_index_for_a2 <= 497;
        o_index_for_a3 <= 769;
        o_index_for_a4 <= 935;
        o_index_for_a5 <= 1099; 
    end
    554: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 96;
        o_index_for_a1 <= 251;
        o_index_for_a2 <= 498;
        o_index_for_a3 <= 770;
        o_index_for_a4 <= 936;
        o_index_for_a5 <= 1100; 
    end
    555: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 97;
        o_index_for_a1 <= 252;
        o_index_for_a2 <= 499;
        o_index_for_a3 <= 771;
        o_index_for_a4 <= 937;
        o_index_for_a5 <= 1101; 
    end
    556: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 98;
        o_index_for_a1 <= 253;
        o_index_for_a2 <= 500;
        o_index_for_a3 <= 772;
        o_index_for_a4 <= 938;
        o_index_for_a5 <= 1102; 
    end
    557: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 99;
        o_index_for_a1 <= 254;
        o_index_for_a2 <= 501;
        o_index_for_a3 <= 773;
        o_index_for_a4 <= 939;
        o_index_for_a5 <= 1103; 
    end
    558: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 100;
        o_index_for_a1 <= 255;
        o_index_for_a2 <= 502;
        o_index_for_a3 <= 774;
        o_index_for_a4 <= 940;
        o_index_for_a5 <= 1104; 
    end
    559: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 101;
        o_index_for_a1 <= 256;
        o_index_for_a2 <= 503;
        o_index_for_a3 <= 775;
        o_index_for_a4 <= 941;
        o_index_for_a5 <= 1105; 
    end
    560: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 102;
        o_index_for_a1 <= 257;
        o_index_for_a2 <= 504;
        o_index_for_a3 <= 776;
        o_index_for_a4 <= 942;
        o_index_for_a5 <= 1106; 
    end
    561: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 103;
        o_index_for_a1 <= 258;
        o_index_for_a2 <= 505;
        o_index_for_a3 <= 777;
        o_index_for_a4 <= 943;
        o_index_for_a5 <= 1107; 
    end
    562: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 104;
        o_index_for_a1 <= 259;
        o_index_for_a2 <= 506;
        o_index_for_a3 <= 778;
        o_index_for_a4 <= 944;
        o_index_for_a5 <= 1108; 
    end
    563: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 105;
        o_index_for_a1 <= 260;
        o_index_for_a2 <= 507;
        o_index_for_a3 <= 779;
        o_index_for_a4 <= 945;
        o_index_for_a5 <= 1109; 
    end
    564: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 106;
        o_index_for_a1 <= 261;
        o_index_for_a2 <= 508;
        o_index_for_a3 <= 780;
        o_index_for_a4 <= 946;
        o_index_for_a5 <= 1110; 
    end
    565: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 107;
        o_index_for_a1 <= 262;
        o_index_for_a2 <= 509;
        o_index_for_a3 <= 781;
        o_index_for_a4 <= 947;
        o_index_for_a5 <= 1111; 
    end
    566: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 108;
        o_index_for_a1 <= 263;
        o_index_for_a2 <= 510;
        o_index_for_a3 <= 782;
        o_index_for_a4 <= 948;
        o_index_for_a5 <= 1112; 
    end
    567: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 109;
        o_index_for_a1 <= 264;
        o_index_for_a2 <= 511;
        o_index_for_a3 <= 783;
        o_index_for_a4 <= 949;
        o_index_for_a5 <= 1113; 
    end
    568: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 110;
        o_index_for_a1 <= 265;
        o_index_for_a2 <= 512;
        o_index_for_a3 <= 784;
        o_index_for_a4 <= 950;
        o_index_for_a5 <= 1114; 
    end
    569: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 111;
        o_index_for_a1 <= 266;
        o_index_for_a2 <= 513;
        o_index_for_a3 <= 785;
        o_index_for_a4 <= 951;
        o_index_for_a5 <= 1115; 
    end
    570: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 112;
        o_index_for_a1 <= 267;
        o_index_for_a2 <= 514;
        o_index_for_a3 <= 786;
        o_index_for_a4 <= 952;
        o_index_for_a5 <= 1116; 
    end
    571: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 113;
        o_index_for_a1 <= 268;
        o_index_for_a2 <= 515;
        o_index_for_a3 <= 787;
        o_index_for_a4 <= 953;
        o_index_for_a5 <= 1117; 
    end
    572: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 114;
        o_index_for_a1 <= 269;
        o_index_for_a2 <= 516;
        o_index_for_a3 <= 788;
        o_index_for_a4 <= 954;
        o_index_for_a5 <= 1118; 
    end
    573: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 115;
        o_index_for_a1 <= 270;
        o_index_for_a2 <= 517;
        o_index_for_a3 <= 789;
        o_index_for_a4 <= 955;
        o_index_for_a5 <= 1119; 
    end
    574: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 116;
        o_index_for_a1 <= 271;
        o_index_for_a2 <= 518;
        o_index_for_a3 <= 790;
        o_index_for_a4 <= 956;
        o_index_for_a5 <= 1120; 
    end
    575: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_index_for_a0 <= 117;
        o_index_for_a1 <= 272;
        o_index_for_a2 <= 519;
        o_index_for_a3 <= 791;
        o_index_for_a4 <= 957;
        o_index_for_a5 <= 1121; 
    end
    576: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 175;
        o_index_for_a1 <= 468;
        o_index_for_a2 <= 674;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    577: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 176;
        o_index_for_a1 <= 469;
        o_index_for_a2 <= 675;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    578: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 177;
        o_index_for_a1 <= 470;
        o_index_for_a2 <= 676;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    579: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 178;
        o_index_for_a1 <= 471;
        o_index_for_a2 <= 677;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    580: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 179;
        o_index_for_a1 <= 472;
        o_index_for_a2 <= 678;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    581: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 180;
        o_index_for_a1 <= 473;
        o_index_for_a2 <= 679;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    582: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 181;
        o_index_for_a1 <= 474;
        o_index_for_a2 <= 680;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    583: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 182;
        o_index_for_a1 <= 475;
        o_index_for_a2 <= 681;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    584: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 183;
        o_index_for_a1 <= 476;
        o_index_for_a2 <= 682;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    585: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 184;
        o_index_for_a1 <= 477;
        o_index_for_a2 <= 683;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    586: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 185;
        o_index_for_a1 <= 478;
        o_index_for_a2 <= 684;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    587: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 186;
        o_index_for_a1 <= 479;
        o_index_for_a2 <= 685;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    588: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 187;
        o_index_for_a1 <= 384;
        o_index_for_a2 <= 686;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    589: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 188;
        o_index_for_a1 <= 385;
        o_index_for_a2 <= 687;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    590: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 189;
        o_index_for_a1 <= 386;
        o_index_for_a2 <= 688;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    591: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 190;
        o_index_for_a1 <= 387;
        o_index_for_a2 <= 689;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    592: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 191;
        o_index_for_a1 <= 388;
        o_index_for_a2 <= 690;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    593: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 96;
        o_index_for_a1 <= 389;
        o_index_for_a2 <= 691;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    594: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 97;
        o_index_for_a1 <= 390;
        o_index_for_a2 <= 692;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    595: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 98;
        o_index_for_a1 <= 391;
        o_index_for_a2 <= 693;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    596: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 99;
        o_index_for_a1 <= 392;
        o_index_for_a2 <= 694;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    597: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 100;
        o_index_for_a1 <= 393;
        o_index_for_a2 <= 695;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    598: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 101;
        o_index_for_a1 <= 394;
        o_index_for_a2 <= 696;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    599: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 102;
        o_index_for_a1 <= 395;
        o_index_for_a2 <= 697;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    600: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 103;
        o_index_for_a1 <= 396;
        o_index_for_a2 <= 698;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    601: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 104;
        o_index_for_a1 <= 397;
        o_index_for_a2 <= 699;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    602: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 105;
        o_index_for_a1 <= 398;
        o_index_for_a2 <= 700;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    603: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 106;
        o_index_for_a1 <= 399;
        o_index_for_a2 <= 701;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    604: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 107;
        o_index_for_a1 <= 400;
        o_index_for_a2 <= 702;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    605: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 108;
        o_index_for_a1 <= 401;
        o_index_for_a2 <= 703;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    606: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 109;
        o_index_for_a1 <= 402;
        o_index_for_a2 <= 704;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    607: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 110;
        o_index_for_a1 <= 403;
        o_index_for_a2 <= 705;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    608: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 111;
        o_index_for_a1 <= 404;
        o_index_for_a2 <= 706;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    609: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 112;
        o_index_for_a1 <= 405;
        o_index_for_a2 <= 707;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    610: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 113;
        o_index_for_a1 <= 406;
        o_index_for_a2 <= 708;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    611: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 114;
        o_index_for_a1 <= 407;
        o_index_for_a2 <= 709;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    612: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 115;
        o_index_for_a1 <= 408;
        o_index_for_a2 <= 710;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    613: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 116;
        o_index_for_a1 <= 409;
        o_index_for_a2 <= 711;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    614: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 117;
        o_index_for_a1 <= 410;
        o_index_for_a2 <= 712;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    615: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 118;
        o_index_for_a1 <= 411;
        o_index_for_a2 <= 713;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    616: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 119;
        o_index_for_a1 <= 412;
        o_index_for_a2 <= 714;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    617: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 120;
        o_index_for_a1 <= 413;
        o_index_for_a2 <= 715;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    618: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 121;
        o_index_for_a1 <= 414;
        o_index_for_a2 <= 716;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    619: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 122;
        o_index_for_a1 <= 415;
        o_index_for_a2 <= 717;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    620: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 123;
        o_index_for_a1 <= 416;
        o_index_for_a2 <= 718;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    621: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 124;
        o_index_for_a1 <= 417;
        o_index_for_a2 <= 719;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    622: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 125;
        o_index_for_a1 <= 418;
        o_index_for_a2 <= 720;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    623: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 126;
        o_index_for_a1 <= 419;
        o_index_for_a2 <= 721;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    624: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 127;
        o_index_for_a1 <= 420;
        o_index_for_a2 <= 722;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    625: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 128;
        o_index_for_a1 <= 421;
        o_index_for_a2 <= 723;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    626: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 129;
        o_index_for_a1 <= 422;
        o_index_for_a2 <= 724;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    627: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 130;
        o_index_for_a1 <= 423;
        o_index_for_a2 <= 725;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    628: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 131;
        o_index_for_a1 <= 424;
        o_index_for_a2 <= 726;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    629: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 132;
        o_index_for_a1 <= 425;
        o_index_for_a2 <= 727;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    630: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 133;
        o_index_for_a1 <= 426;
        o_index_for_a2 <= 728;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    631: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 134;
        o_index_for_a1 <= 427;
        o_index_for_a2 <= 729;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    632: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 135;
        o_index_for_a1 <= 428;
        o_index_for_a2 <= 730;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    633: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 136;
        o_index_for_a1 <= 429;
        o_index_for_a2 <= 731;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    634: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 137;
        o_index_for_a1 <= 430;
        o_index_for_a2 <= 732;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    635: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 138;
        o_index_for_a1 <= 431;
        o_index_for_a2 <= 733;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    636: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 139;
        o_index_for_a1 <= 432;
        o_index_for_a2 <= 734;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    637: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 140;
        o_index_for_a1 <= 433;
        o_index_for_a2 <= 735;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    638: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 141;
        o_index_for_a1 <= 434;
        o_index_for_a2 <= 736;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    639: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 142;
        o_index_for_a1 <= 435;
        o_index_for_a2 <= 737;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    640: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 143;
        o_index_for_a1 <= 436;
        o_index_for_a2 <= 738;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    641: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 144;
        o_index_for_a1 <= 437;
        o_index_for_a2 <= 739;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    642: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 145;
        o_index_for_a1 <= 438;
        o_index_for_a2 <= 740;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    643: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 146;
        o_index_for_a1 <= 439;
        o_index_for_a2 <= 741;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    644: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 147;
        o_index_for_a1 <= 440;
        o_index_for_a2 <= 742;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    645: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 148;
        o_index_for_a1 <= 441;
        o_index_for_a2 <= 743;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    646: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 149;
        o_index_for_a1 <= 442;
        o_index_for_a2 <= 744;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    647: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 150;
        o_index_for_a1 <= 443;
        o_index_for_a2 <= 745;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    648: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 151;
        o_index_for_a1 <= 444;
        o_index_for_a2 <= 746;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    649: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 152;
        o_index_for_a1 <= 445;
        o_index_for_a2 <= 747;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    650: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 153;
        o_index_for_a1 <= 446;
        o_index_for_a2 <= 748;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    651: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 154;
        o_index_for_a1 <= 447;
        o_index_for_a2 <= 749;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    652: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 155;
        o_index_for_a1 <= 448;
        o_index_for_a2 <= 750;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    653: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 156;
        o_index_for_a1 <= 449;
        o_index_for_a2 <= 751;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    654: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 157;
        o_index_for_a1 <= 450;
        o_index_for_a2 <= 752;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    655: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 158;
        o_index_for_a1 <= 451;
        o_index_for_a2 <= 753;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    656: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 159;
        o_index_for_a1 <= 452;
        o_index_for_a2 <= 754;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    657: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 160;
        o_index_for_a1 <= 453;
        o_index_for_a2 <= 755;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    658: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 161;
        o_index_for_a1 <= 454;
        o_index_for_a2 <= 756;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    659: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 162;
        o_index_for_a1 <= 455;
        o_index_for_a2 <= 757;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    660: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 163;
        o_index_for_a1 <= 456;
        o_index_for_a2 <= 758;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    661: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 164;
        o_index_for_a1 <= 457;
        o_index_for_a2 <= 759;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    662: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 165;
        o_index_for_a1 <= 458;
        o_index_for_a2 <= 760;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    663: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 166;
        o_index_for_a1 <= 459;
        o_index_for_a2 <= 761;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    664: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 167;
        o_index_for_a1 <= 460;
        o_index_for_a2 <= 762;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    665: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 168;
        o_index_for_a1 <= 461;
        o_index_for_a2 <= 763;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    666: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 169;
        o_index_for_a1 <= 462;
        o_index_for_a2 <= 764;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    667: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 170;
        o_index_for_a1 <= 463;
        o_index_for_a2 <= 765;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    668: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 171;
        o_index_for_a1 <= 464;
        o_index_for_a2 <= 766;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    669: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 172;
        o_index_for_a1 <= 465;
        o_index_for_a2 <= 767;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    670: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 173;
        o_index_for_a1 <= 466;
        o_index_for_a2 <= 672;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    671: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 174;
        o_index_for_a1 <= 467;
        o_index_for_a2 <= 673;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    672: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 105;
        o_index_for_a1 <= 225;
        o_index_for_a2 <= 562;
        o_index_for_a3 <= 811;
        o_index_for_a4 <= 923;
        o_index_for_a5 <= 1097; 
    end
    673: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 106;
        o_index_for_a1 <= 226;
        o_index_for_a2 <= 563;
        o_index_for_a3 <= 812;
        o_index_for_a4 <= 924;
        o_index_for_a5 <= 1098; 
    end
    674: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 107;
        o_index_for_a1 <= 227;
        o_index_for_a2 <= 564;
        o_index_for_a3 <= 813;
        o_index_for_a4 <= 925;
        o_index_for_a5 <= 1099; 
    end
    675: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 108;
        o_index_for_a1 <= 228;
        o_index_for_a2 <= 565;
        o_index_for_a3 <= 814;
        o_index_for_a4 <= 926;
        o_index_for_a5 <= 1100; 
    end
    676: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 109;
        o_index_for_a1 <= 229;
        o_index_for_a2 <= 566;
        o_index_for_a3 <= 815;
        o_index_for_a4 <= 927;
        o_index_for_a5 <= 1101; 
    end
    677: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 110;
        o_index_for_a1 <= 230;
        o_index_for_a2 <= 567;
        o_index_for_a3 <= 816;
        o_index_for_a4 <= 928;
        o_index_for_a5 <= 1102; 
    end
    678: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 111;
        o_index_for_a1 <= 231;
        o_index_for_a2 <= 568;
        o_index_for_a3 <= 817;
        o_index_for_a4 <= 929;
        o_index_for_a5 <= 1103; 
    end
    679: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 112;
        o_index_for_a1 <= 232;
        o_index_for_a2 <= 569;
        o_index_for_a3 <= 818;
        o_index_for_a4 <= 930;
        o_index_for_a5 <= 1104; 
    end
    680: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 113;
        o_index_for_a1 <= 233;
        o_index_for_a2 <= 570;
        o_index_for_a3 <= 819;
        o_index_for_a4 <= 931;
        o_index_for_a5 <= 1105; 
    end
    681: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 114;
        o_index_for_a1 <= 234;
        o_index_for_a2 <= 571;
        o_index_for_a3 <= 820;
        o_index_for_a4 <= 932;
        o_index_for_a5 <= 1106; 
    end
    682: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 115;
        o_index_for_a1 <= 235;
        o_index_for_a2 <= 572;
        o_index_for_a3 <= 821;
        o_index_for_a4 <= 933;
        o_index_for_a5 <= 1107; 
    end
    683: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 116;
        o_index_for_a1 <= 236;
        o_index_for_a2 <= 573;
        o_index_for_a3 <= 822;
        o_index_for_a4 <= 934;
        o_index_for_a5 <= 1108; 
    end
    684: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 117;
        o_index_for_a1 <= 237;
        o_index_for_a2 <= 574;
        o_index_for_a3 <= 823;
        o_index_for_a4 <= 935;
        o_index_for_a5 <= 1109; 
    end
    685: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 118;
        o_index_for_a1 <= 238;
        o_index_for_a2 <= 575;
        o_index_for_a3 <= 824;
        o_index_for_a4 <= 936;
        o_index_for_a5 <= 1110; 
    end
    686: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 119;
        o_index_for_a1 <= 239;
        o_index_for_a2 <= 480;
        o_index_for_a3 <= 825;
        o_index_for_a4 <= 937;
        o_index_for_a5 <= 1111; 
    end
    687: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 120;
        o_index_for_a1 <= 240;
        o_index_for_a2 <= 481;
        o_index_for_a3 <= 826;
        o_index_for_a4 <= 938;
        o_index_for_a5 <= 1112; 
    end
    688: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 121;
        o_index_for_a1 <= 241;
        o_index_for_a2 <= 482;
        o_index_for_a3 <= 827;
        o_index_for_a4 <= 939;
        o_index_for_a5 <= 1113; 
    end
    689: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 122;
        o_index_for_a1 <= 242;
        o_index_for_a2 <= 483;
        o_index_for_a3 <= 828;
        o_index_for_a4 <= 940;
        o_index_for_a5 <= 1114; 
    end
    690: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 123;
        o_index_for_a1 <= 243;
        o_index_for_a2 <= 484;
        o_index_for_a3 <= 829;
        o_index_for_a4 <= 941;
        o_index_for_a5 <= 1115; 
    end
    691: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 124;
        o_index_for_a1 <= 244;
        o_index_for_a2 <= 485;
        o_index_for_a3 <= 830;
        o_index_for_a4 <= 942;
        o_index_for_a5 <= 1116; 
    end
    692: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 125;
        o_index_for_a1 <= 245;
        o_index_for_a2 <= 486;
        o_index_for_a3 <= 831;
        o_index_for_a4 <= 943;
        o_index_for_a5 <= 1117; 
    end
    693: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 126;
        o_index_for_a1 <= 246;
        o_index_for_a2 <= 487;
        o_index_for_a3 <= 832;
        o_index_for_a4 <= 944;
        o_index_for_a5 <= 1118; 
    end
    694: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 127;
        o_index_for_a1 <= 247;
        o_index_for_a2 <= 488;
        o_index_for_a3 <= 833;
        o_index_for_a4 <= 945;
        o_index_for_a5 <= 1119; 
    end
    695: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 128;
        o_index_for_a1 <= 248;
        o_index_for_a2 <= 489;
        o_index_for_a3 <= 834;
        o_index_for_a4 <= 946;
        o_index_for_a5 <= 1120; 
    end
    696: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 129;
        o_index_for_a1 <= 249;
        o_index_for_a2 <= 490;
        o_index_for_a3 <= 835;
        o_index_for_a4 <= 947;
        o_index_for_a5 <= 1121; 
    end
    697: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 130;
        o_index_for_a1 <= 250;
        o_index_for_a2 <= 491;
        o_index_for_a3 <= 836;
        o_index_for_a4 <= 948;
        o_index_for_a5 <= 1122; 
    end
    698: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 131;
        o_index_for_a1 <= 251;
        o_index_for_a2 <= 492;
        o_index_for_a3 <= 837;
        o_index_for_a4 <= 949;
        o_index_for_a5 <= 1123; 
    end
    699: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 132;
        o_index_for_a1 <= 252;
        o_index_for_a2 <= 493;
        o_index_for_a3 <= 838;
        o_index_for_a4 <= 950;
        o_index_for_a5 <= 1124; 
    end
    700: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 133;
        o_index_for_a1 <= 253;
        o_index_for_a2 <= 494;
        o_index_for_a3 <= 839;
        o_index_for_a4 <= 951;
        o_index_for_a5 <= 1125; 
    end
    701: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 134;
        o_index_for_a1 <= 254;
        o_index_for_a2 <= 495;
        o_index_for_a3 <= 840;
        o_index_for_a4 <= 952;
        o_index_for_a5 <= 1126; 
    end
    702: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 135;
        o_index_for_a1 <= 255;
        o_index_for_a2 <= 496;
        o_index_for_a3 <= 841;
        o_index_for_a4 <= 953;
        o_index_for_a5 <= 1127; 
    end
    703: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 136;
        o_index_for_a1 <= 256;
        o_index_for_a2 <= 497;
        o_index_for_a3 <= 842;
        o_index_for_a4 <= 954;
        o_index_for_a5 <= 1128; 
    end
    704: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 137;
        o_index_for_a1 <= 257;
        o_index_for_a2 <= 498;
        o_index_for_a3 <= 843;
        o_index_for_a4 <= 955;
        o_index_for_a5 <= 1129; 
    end
    705: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 138;
        o_index_for_a1 <= 258;
        o_index_for_a2 <= 499;
        o_index_for_a3 <= 844;
        o_index_for_a4 <= 956;
        o_index_for_a5 <= 1130; 
    end
    706: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 139;
        o_index_for_a1 <= 259;
        o_index_for_a2 <= 500;
        o_index_for_a3 <= 845;
        o_index_for_a4 <= 957;
        o_index_for_a5 <= 1131; 
    end
    707: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 140;
        o_index_for_a1 <= 260;
        o_index_for_a2 <= 501;
        o_index_for_a3 <= 846;
        o_index_for_a4 <= 958;
        o_index_for_a5 <= 1132; 
    end
    708: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 141;
        o_index_for_a1 <= 261;
        o_index_for_a2 <= 502;
        o_index_for_a3 <= 847;
        o_index_for_a4 <= 959;
        o_index_for_a5 <= 1133; 
    end
    709: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 142;
        o_index_for_a1 <= 262;
        o_index_for_a2 <= 503;
        o_index_for_a3 <= 848;
        o_index_for_a4 <= 864;
        o_index_for_a5 <= 1134; 
    end
    710: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 143;
        o_index_for_a1 <= 263;
        o_index_for_a2 <= 504;
        o_index_for_a3 <= 849;
        o_index_for_a4 <= 865;
        o_index_for_a5 <= 1135; 
    end
    711: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 144;
        o_index_for_a1 <= 264;
        o_index_for_a2 <= 505;
        o_index_for_a3 <= 850;
        o_index_for_a4 <= 866;
        o_index_for_a5 <= 1136; 
    end
    712: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 145;
        o_index_for_a1 <= 265;
        o_index_for_a2 <= 506;
        o_index_for_a3 <= 851;
        o_index_for_a4 <= 867;
        o_index_for_a5 <= 1137; 
    end
    713: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 146;
        o_index_for_a1 <= 266;
        o_index_for_a2 <= 507;
        o_index_for_a3 <= 852;
        o_index_for_a4 <= 868;
        o_index_for_a5 <= 1138; 
    end
    714: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 147;
        o_index_for_a1 <= 267;
        o_index_for_a2 <= 508;
        o_index_for_a3 <= 853;
        o_index_for_a4 <= 869;
        o_index_for_a5 <= 1139; 
    end
    715: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 148;
        o_index_for_a1 <= 268;
        o_index_for_a2 <= 509;
        o_index_for_a3 <= 854;
        o_index_for_a4 <= 870;
        o_index_for_a5 <= 1140; 
    end
    716: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 149;
        o_index_for_a1 <= 269;
        o_index_for_a2 <= 510;
        o_index_for_a3 <= 855;
        o_index_for_a4 <= 871;
        o_index_for_a5 <= 1141; 
    end
    717: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 150;
        o_index_for_a1 <= 270;
        o_index_for_a2 <= 511;
        o_index_for_a3 <= 856;
        o_index_for_a4 <= 872;
        o_index_for_a5 <= 1142; 
    end
    718: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 151;
        o_index_for_a1 <= 271;
        o_index_for_a2 <= 512;
        o_index_for_a3 <= 857;
        o_index_for_a4 <= 873;
        o_index_for_a5 <= 1143; 
    end
    719: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 152;
        o_index_for_a1 <= 272;
        o_index_for_a2 <= 513;
        o_index_for_a3 <= 858;
        o_index_for_a4 <= 874;
        o_index_for_a5 <= 1144; 
    end
    720: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 153;
        o_index_for_a1 <= 273;
        o_index_for_a2 <= 514;
        o_index_for_a3 <= 859;
        o_index_for_a4 <= 875;
        o_index_for_a5 <= 1145; 
    end
    721: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 154;
        o_index_for_a1 <= 274;
        o_index_for_a2 <= 515;
        o_index_for_a3 <= 860;
        o_index_for_a4 <= 876;
        o_index_for_a5 <= 1146; 
    end
    722: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 155;
        o_index_for_a1 <= 275;
        o_index_for_a2 <= 516;
        o_index_for_a3 <= 861;
        o_index_for_a4 <= 877;
        o_index_for_a5 <= 1147; 
    end
    723: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 156;
        o_index_for_a1 <= 276;
        o_index_for_a2 <= 517;
        o_index_for_a3 <= 862;
        o_index_for_a4 <= 878;
        o_index_for_a5 <= 1148; 
    end
    724: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 157;
        o_index_for_a1 <= 277;
        o_index_for_a2 <= 518;
        o_index_for_a3 <= 863;
        o_index_for_a4 <= 879;
        o_index_for_a5 <= 1149; 
    end
    725: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 158;
        o_index_for_a1 <= 278;
        o_index_for_a2 <= 519;
        o_index_for_a3 <= 768;
        o_index_for_a4 <= 880;
        o_index_for_a5 <= 1150; 
    end
    726: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 159;
        o_index_for_a1 <= 279;
        o_index_for_a2 <= 520;
        o_index_for_a3 <= 769;
        o_index_for_a4 <= 881;
        o_index_for_a5 <= 1151; 
    end
    727: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 160;
        o_index_for_a1 <= 280;
        o_index_for_a2 <= 521;
        o_index_for_a3 <= 770;
        o_index_for_a4 <= 882;
        o_index_for_a5 <= 1056; 
    end
    728: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 161;
        o_index_for_a1 <= 281;
        o_index_for_a2 <= 522;
        o_index_for_a3 <= 771;
        o_index_for_a4 <= 883;
        o_index_for_a5 <= 1057; 
    end
    729: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 162;
        o_index_for_a1 <= 282;
        o_index_for_a2 <= 523;
        o_index_for_a3 <= 772;
        o_index_for_a4 <= 884;
        o_index_for_a5 <= 1058; 
    end
    730: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 163;
        o_index_for_a1 <= 283;
        o_index_for_a2 <= 524;
        o_index_for_a3 <= 773;
        o_index_for_a4 <= 885;
        o_index_for_a5 <= 1059; 
    end
    731: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 164;
        o_index_for_a1 <= 284;
        o_index_for_a2 <= 525;
        o_index_for_a3 <= 774;
        o_index_for_a4 <= 886;
        o_index_for_a5 <= 1060; 
    end
    732: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 165;
        o_index_for_a1 <= 285;
        o_index_for_a2 <= 526;
        o_index_for_a3 <= 775;
        o_index_for_a4 <= 887;
        o_index_for_a5 <= 1061; 
    end
    733: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 166;
        o_index_for_a1 <= 286;
        o_index_for_a2 <= 527;
        o_index_for_a3 <= 776;
        o_index_for_a4 <= 888;
        o_index_for_a5 <= 1062; 
    end
    734: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 167;
        o_index_for_a1 <= 287;
        o_index_for_a2 <= 528;
        o_index_for_a3 <= 777;
        o_index_for_a4 <= 889;
        o_index_for_a5 <= 1063; 
    end
    735: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 168;
        o_index_for_a1 <= 192;
        o_index_for_a2 <= 529;
        o_index_for_a3 <= 778;
        o_index_for_a4 <= 890;
        o_index_for_a5 <= 1064; 
    end
    736: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 169;
        o_index_for_a1 <= 193;
        o_index_for_a2 <= 530;
        o_index_for_a3 <= 779;
        o_index_for_a4 <= 891;
        o_index_for_a5 <= 1065; 
    end
    737: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 170;
        o_index_for_a1 <= 194;
        o_index_for_a2 <= 531;
        o_index_for_a3 <= 780;
        o_index_for_a4 <= 892;
        o_index_for_a5 <= 1066; 
    end
    738: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 171;
        o_index_for_a1 <= 195;
        o_index_for_a2 <= 532;
        o_index_for_a3 <= 781;
        o_index_for_a4 <= 893;
        o_index_for_a5 <= 1067; 
    end
    739: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 172;
        o_index_for_a1 <= 196;
        o_index_for_a2 <= 533;
        o_index_for_a3 <= 782;
        o_index_for_a4 <= 894;
        o_index_for_a5 <= 1068; 
    end
    740: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 173;
        o_index_for_a1 <= 197;
        o_index_for_a2 <= 534;
        o_index_for_a3 <= 783;
        o_index_for_a4 <= 895;
        o_index_for_a5 <= 1069; 
    end
    741: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 174;
        o_index_for_a1 <= 198;
        o_index_for_a2 <= 535;
        o_index_for_a3 <= 784;
        o_index_for_a4 <= 896;
        o_index_for_a5 <= 1070; 
    end
    742: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 175;
        o_index_for_a1 <= 199;
        o_index_for_a2 <= 536;
        o_index_for_a3 <= 785;
        o_index_for_a4 <= 897;
        o_index_for_a5 <= 1071; 
    end
    743: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 176;
        o_index_for_a1 <= 200;
        o_index_for_a2 <= 537;
        o_index_for_a3 <= 786;
        o_index_for_a4 <= 898;
        o_index_for_a5 <= 1072; 
    end
    744: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 177;
        o_index_for_a1 <= 201;
        o_index_for_a2 <= 538;
        o_index_for_a3 <= 787;
        o_index_for_a4 <= 899;
        o_index_for_a5 <= 1073; 
    end
    745: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 178;
        o_index_for_a1 <= 202;
        o_index_for_a2 <= 539;
        o_index_for_a3 <= 788;
        o_index_for_a4 <= 900;
        o_index_for_a5 <= 1074; 
    end
    746: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 179;
        o_index_for_a1 <= 203;
        o_index_for_a2 <= 540;
        o_index_for_a3 <= 789;
        o_index_for_a4 <= 901;
        o_index_for_a5 <= 1075; 
    end
    747: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 180;
        o_index_for_a1 <= 204;
        o_index_for_a2 <= 541;
        o_index_for_a3 <= 790;
        o_index_for_a4 <= 902;
        o_index_for_a5 <= 1076; 
    end
    748: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 181;
        o_index_for_a1 <= 205;
        o_index_for_a2 <= 542;
        o_index_for_a3 <= 791;
        o_index_for_a4 <= 903;
        o_index_for_a5 <= 1077; 
    end
    749: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 182;
        o_index_for_a1 <= 206;
        o_index_for_a2 <= 543;
        o_index_for_a3 <= 792;
        o_index_for_a4 <= 904;
        o_index_for_a5 <= 1078; 
    end
    750: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 183;
        o_index_for_a1 <= 207;
        o_index_for_a2 <= 544;
        o_index_for_a3 <= 793;
        o_index_for_a4 <= 905;
        o_index_for_a5 <= 1079; 
    end
    751: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 184;
        o_index_for_a1 <= 208;
        o_index_for_a2 <= 545;
        o_index_for_a3 <= 794;
        o_index_for_a4 <= 906;
        o_index_for_a5 <= 1080; 
    end
    752: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 185;
        o_index_for_a1 <= 209;
        o_index_for_a2 <= 546;
        o_index_for_a3 <= 795;
        o_index_for_a4 <= 907;
        o_index_for_a5 <= 1081; 
    end
    753: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 186;
        o_index_for_a1 <= 210;
        o_index_for_a2 <= 547;
        o_index_for_a3 <= 796;
        o_index_for_a4 <= 908;
        o_index_for_a5 <= 1082; 
    end
    754: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 187;
        o_index_for_a1 <= 211;
        o_index_for_a2 <= 548;
        o_index_for_a3 <= 797;
        o_index_for_a4 <= 909;
        o_index_for_a5 <= 1083; 
    end
    755: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 188;
        o_index_for_a1 <= 212;
        o_index_for_a2 <= 549;
        o_index_for_a3 <= 798;
        o_index_for_a4 <= 910;
        o_index_for_a5 <= 1084; 
    end
    756: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 189;
        o_index_for_a1 <= 213;
        o_index_for_a2 <= 550;
        o_index_for_a3 <= 799;
        o_index_for_a4 <= 911;
        o_index_for_a5 <= 1085; 
    end
    757: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 190;
        o_index_for_a1 <= 214;
        o_index_for_a2 <= 551;
        o_index_for_a3 <= 800;
        o_index_for_a4 <= 912;
        o_index_for_a5 <= 1086; 
    end
    758: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 191;
        o_index_for_a1 <= 215;
        o_index_for_a2 <= 552;
        o_index_for_a3 <= 801;
        o_index_for_a4 <= 913;
        o_index_for_a5 <= 1087; 
    end
    759: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 96;
        o_index_for_a1 <= 216;
        o_index_for_a2 <= 553;
        o_index_for_a3 <= 802;
        o_index_for_a4 <= 914;
        o_index_for_a5 <= 1088; 
    end
    760: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 97;
        o_index_for_a1 <= 217;
        o_index_for_a2 <= 554;
        o_index_for_a3 <= 803;
        o_index_for_a4 <= 915;
        o_index_for_a5 <= 1089; 
    end
    761: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 98;
        o_index_for_a1 <= 218;
        o_index_for_a2 <= 555;
        o_index_for_a3 <= 804;
        o_index_for_a4 <= 916;
        o_index_for_a5 <= 1090; 
    end
    762: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 99;
        o_index_for_a1 <= 219;
        o_index_for_a2 <= 556;
        o_index_for_a3 <= 805;
        o_index_for_a4 <= 917;
        o_index_for_a5 <= 1091; 
    end
    763: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 100;
        o_index_for_a1 <= 220;
        o_index_for_a2 <= 557;
        o_index_for_a3 <= 806;
        o_index_for_a4 <= 918;
        o_index_for_a5 <= 1092; 
    end
    764: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 101;
        o_index_for_a1 <= 221;
        o_index_for_a2 <= 558;
        o_index_for_a3 <= 807;
        o_index_for_a4 <= 919;
        o_index_for_a5 <= 1093; 
    end
    765: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 102;
        o_index_for_a1 <= 222;
        o_index_for_a2 <= 559;
        o_index_for_a3 <= 808;
        o_index_for_a4 <= 920;
        o_index_for_a5 <= 1094; 
    end
    766: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 103;
        o_index_for_a1 <= 223;
        o_index_for_a2 <= 560;
        o_index_for_a3 <= 809;
        o_index_for_a4 <= 921;
        o_index_for_a5 <= 1095; 
    end
    767: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 2; 
        o_index_for_a0 <= 104;
        o_index_for_a1 <= 224;
        o_index_for_a2 <= 561;
        o_index_for_a3 <= 810;
        o_index_for_a4 <= 922;
        o_index_for_a5 <= 1096; 
    end
    768: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 55;
        o_index_for_a1 <= 353;
        o_index_for_a2 <= 999;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    769: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 56;
        o_index_for_a1 <= 354;
        o_index_for_a2 <= 1000;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    770: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 57;
        o_index_for_a1 <= 355;
        o_index_for_a2 <= 1001;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    771: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 58;
        o_index_for_a1 <= 356;
        o_index_for_a2 <= 1002;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    772: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 59;
        o_index_for_a1 <= 357;
        o_index_for_a2 <= 1003;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    773: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 60;
        o_index_for_a1 <= 358;
        o_index_for_a2 <= 1004;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    774: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 61;
        o_index_for_a1 <= 359;
        o_index_for_a2 <= 1005;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    775: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 62;
        o_index_for_a1 <= 360;
        o_index_for_a2 <= 1006;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    776: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 63;
        o_index_for_a1 <= 361;
        o_index_for_a2 <= 1007;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    777: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 64;
        o_index_for_a1 <= 362;
        o_index_for_a2 <= 1008;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    778: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 65;
        o_index_for_a1 <= 363;
        o_index_for_a2 <= 1009;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    779: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 66;
        o_index_for_a1 <= 364;
        o_index_for_a2 <= 1010;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    780: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 67;
        o_index_for_a1 <= 365;
        o_index_for_a2 <= 1011;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    781: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 68;
        o_index_for_a1 <= 366;
        o_index_for_a2 <= 1012;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    782: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 69;
        o_index_for_a1 <= 367;
        o_index_for_a2 <= 1013;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    783: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 70;
        o_index_for_a1 <= 368;
        o_index_for_a2 <= 1014;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    784: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 71;
        o_index_for_a1 <= 369;
        o_index_for_a2 <= 1015;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    785: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 72;
        o_index_for_a1 <= 370;
        o_index_for_a2 <= 1016;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    786: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 73;
        o_index_for_a1 <= 371;
        o_index_for_a2 <= 1017;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    787: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 74;
        o_index_for_a1 <= 372;
        o_index_for_a2 <= 1018;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    788: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 75;
        o_index_for_a1 <= 373;
        o_index_for_a2 <= 1019;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    789: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 76;
        o_index_for_a1 <= 374;
        o_index_for_a2 <= 1020;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    790: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 77;
        o_index_for_a1 <= 375;
        o_index_for_a2 <= 1021;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    791: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 78;
        o_index_for_a1 <= 376;
        o_index_for_a2 <= 1022;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    792: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 79;
        o_index_for_a1 <= 377;
        o_index_for_a2 <= 1023;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    793: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 80;
        o_index_for_a1 <= 378;
        o_index_for_a2 <= 1024;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    794: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 81;
        o_index_for_a1 <= 379;
        o_index_for_a2 <= 1025;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    795: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 82;
        o_index_for_a1 <= 380;
        o_index_for_a2 <= 1026;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    796: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 83;
        o_index_for_a1 <= 381;
        o_index_for_a2 <= 1027;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    797: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 84;
        o_index_for_a1 <= 382;
        o_index_for_a2 <= 1028;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    798: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 85;
        o_index_for_a1 <= 383;
        o_index_for_a2 <= 1029;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    799: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 86;
        o_index_for_a1 <= 288;
        o_index_for_a2 <= 1030;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    800: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 87;
        o_index_for_a1 <= 289;
        o_index_for_a2 <= 1031;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    801: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 88;
        o_index_for_a1 <= 290;
        o_index_for_a2 <= 1032;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    802: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 89;
        o_index_for_a1 <= 291;
        o_index_for_a2 <= 1033;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    803: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 90;
        o_index_for_a1 <= 292;
        o_index_for_a2 <= 1034;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    804: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 91;
        o_index_for_a1 <= 293;
        o_index_for_a2 <= 1035;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    805: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 92;
        o_index_for_a1 <= 294;
        o_index_for_a2 <= 1036;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    806: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 93;
        o_index_for_a1 <= 295;
        o_index_for_a2 <= 1037;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    807: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 94;
        o_index_for_a1 <= 296;
        o_index_for_a2 <= 1038;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    808: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 95;
        o_index_for_a1 <= 297;
        o_index_for_a2 <= 1039;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    809: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 0;
        o_index_for_a1 <= 298;
        o_index_for_a2 <= 1040;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    810: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1;
        o_index_for_a1 <= 299;
        o_index_for_a2 <= 1041;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    811: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 2;
        o_index_for_a1 <= 300;
        o_index_for_a2 <= 1042;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    812: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 3;
        o_index_for_a1 <= 301;
        o_index_for_a2 <= 1043;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    813: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 4;
        o_index_for_a1 <= 302;
        o_index_for_a2 <= 1044;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    814: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 5;
        o_index_for_a1 <= 303;
        o_index_for_a2 <= 1045;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    815: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 6;
        o_index_for_a1 <= 304;
        o_index_for_a2 <= 1046;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    816: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 7;
        o_index_for_a1 <= 305;
        o_index_for_a2 <= 1047;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    817: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 8;
        o_index_for_a1 <= 306;
        o_index_for_a2 <= 1048;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    818: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 9;
        o_index_for_a1 <= 307;
        o_index_for_a2 <= 1049;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    819: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 10;
        o_index_for_a1 <= 308;
        o_index_for_a2 <= 1050;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    820: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 11;
        o_index_for_a1 <= 309;
        o_index_for_a2 <= 1051;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    821: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 12;
        o_index_for_a1 <= 310;
        o_index_for_a2 <= 1052;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    822: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 13;
        o_index_for_a1 <= 311;
        o_index_for_a2 <= 1053;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    823: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 14;
        o_index_for_a1 <= 312;
        o_index_for_a2 <= 1054;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    824: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 15;
        o_index_for_a1 <= 313;
        o_index_for_a2 <= 1055;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    825: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 16;
        o_index_for_a1 <= 314;
        o_index_for_a2 <= 960;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    826: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 17;
        o_index_for_a1 <= 315;
        o_index_for_a2 <= 961;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    827: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 18;
        o_index_for_a1 <= 316;
        o_index_for_a2 <= 962;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    828: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 19;
        o_index_for_a1 <= 317;
        o_index_for_a2 <= 963;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    829: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 20;
        o_index_for_a1 <= 318;
        o_index_for_a2 <= 964;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    830: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 21;
        o_index_for_a1 <= 319;
        o_index_for_a2 <= 965;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    831: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 22;
        o_index_for_a1 <= 320;
        o_index_for_a2 <= 966;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    832: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 23;
        o_index_for_a1 <= 321;
        o_index_for_a2 <= 967;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    833: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 24;
        o_index_for_a1 <= 322;
        o_index_for_a2 <= 968;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    834: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 25;
        o_index_for_a1 <= 323;
        o_index_for_a2 <= 969;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    835: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 26;
        o_index_for_a1 <= 324;
        o_index_for_a2 <= 970;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    836: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 27;
        o_index_for_a1 <= 325;
        o_index_for_a2 <= 971;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    837: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 28;
        o_index_for_a1 <= 326;
        o_index_for_a2 <= 972;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    838: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 29;
        o_index_for_a1 <= 327;
        o_index_for_a2 <= 973;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    839: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 30;
        o_index_for_a1 <= 328;
        o_index_for_a2 <= 974;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    840: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 31;
        o_index_for_a1 <= 329;
        o_index_for_a2 <= 975;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    841: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 32;
        o_index_for_a1 <= 330;
        o_index_for_a2 <= 976;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    842: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 33;
        o_index_for_a1 <= 331;
        o_index_for_a2 <= 977;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    843: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 34;
        o_index_for_a1 <= 332;
        o_index_for_a2 <= 978;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    844: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 35;
        o_index_for_a1 <= 333;
        o_index_for_a2 <= 979;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    845: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 36;
        o_index_for_a1 <= 334;
        o_index_for_a2 <= 980;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    846: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 37;
        o_index_for_a1 <= 335;
        o_index_for_a2 <= 981;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    847: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 38;
        o_index_for_a1 <= 336;
        o_index_for_a2 <= 982;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    848: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 39;
        o_index_for_a1 <= 337;
        o_index_for_a2 <= 983;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    849: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 40;
        o_index_for_a1 <= 338;
        o_index_for_a2 <= 984;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    850: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 41;
        o_index_for_a1 <= 339;
        o_index_for_a2 <= 985;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    851: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 42;
        o_index_for_a1 <= 340;
        o_index_for_a2 <= 986;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    852: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 43;
        o_index_for_a1 <= 341;
        o_index_for_a2 <= 987;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    853: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 44;
        o_index_for_a1 <= 342;
        o_index_for_a2 <= 988;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    854: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 45;
        o_index_for_a1 <= 343;
        o_index_for_a2 <= 989;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    855: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 46;
        o_index_for_a1 <= 344;
        o_index_for_a2 <= 990;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    856: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 47;
        o_index_for_a1 <= 345;
        o_index_for_a2 <= 991;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    857: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 48;
        o_index_for_a1 <= 346;
        o_index_for_a2 <= 992;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    858: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 49;
        o_index_for_a1 <= 347;
        o_index_for_a2 <= 993;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    859: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 50;
        o_index_for_a1 <= 348;
        o_index_for_a2 <= 994;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    860: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 51;
        o_index_for_a1 <= 349;
        o_index_for_a2 <= 995;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    861: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 52;
        o_index_for_a1 <= 350;
        o_index_for_a2 <= 996;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    862: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 53;
        o_index_for_a1 <= 351;
        o_index_for_a2 <= 997;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    863: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 54;
        o_index_for_a1 <= 352;
        o_index_for_a2 <= 998;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    864: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 83;
        o_index_for_a1 <= 313;
        o_index_for_a2 <= 425;
        o_index_for_a3 <= 590;
        o_index_for_a4 <= 719;
        o_index_for_a5 <= 1009; 
    end
    865: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 84;
        o_index_for_a1 <= 314;
        o_index_for_a2 <= 426;
        o_index_for_a3 <= 591;
        o_index_for_a4 <= 720;
        o_index_for_a5 <= 1010; 
    end
    866: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 85;
        o_index_for_a1 <= 315;
        o_index_for_a2 <= 427;
        o_index_for_a3 <= 592;
        o_index_for_a4 <= 721;
        o_index_for_a5 <= 1011; 
    end
    867: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 86;
        o_index_for_a1 <= 316;
        o_index_for_a2 <= 428;
        o_index_for_a3 <= 593;
        o_index_for_a4 <= 722;
        o_index_for_a5 <= 1012; 
    end
    868: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 87;
        o_index_for_a1 <= 317;
        o_index_for_a2 <= 429;
        o_index_for_a3 <= 594;
        o_index_for_a4 <= 723;
        o_index_for_a5 <= 1013; 
    end
    869: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 88;
        o_index_for_a1 <= 318;
        o_index_for_a2 <= 430;
        o_index_for_a3 <= 595;
        o_index_for_a4 <= 724;
        o_index_for_a5 <= 1014; 
    end
    870: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 89;
        o_index_for_a1 <= 319;
        o_index_for_a2 <= 431;
        o_index_for_a3 <= 596;
        o_index_for_a4 <= 725;
        o_index_for_a5 <= 1015; 
    end
    871: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 90;
        o_index_for_a1 <= 320;
        o_index_for_a2 <= 432;
        o_index_for_a3 <= 597;
        o_index_for_a4 <= 726;
        o_index_for_a5 <= 1016; 
    end
    872: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 91;
        o_index_for_a1 <= 321;
        o_index_for_a2 <= 433;
        o_index_for_a3 <= 598;
        o_index_for_a4 <= 727;
        o_index_for_a5 <= 1017; 
    end
    873: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 92;
        o_index_for_a1 <= 322;
        o_index_for_a2 <= 434;
        o_index_for_a3 <= 599;
        o_index_for_a4 <= 728;
        o_index_for_a5 <= 1018; 
    end
    874: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 93;
        o_index_for_a1 <= 323;
        o_index_for_a2 <= 435;
        o_index_for_a3 <= 600;
        o_index_for_a4 <= 729;
        o_index_for_a5 <= 1019; 
    end
    875: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 94;
        o_index_for_a1 <= 324;
        o_index_for_a2 <= 436;
        o_index_for_a3 <= 601;
        o_index_for_a4 <= 730;
        o_index_for_a5 <= 1020; 
    end
    876: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 95;
        o_index_for_a1 <= 325;
        o_index_for_a2 <= 437;
        o_index_for_a3 <= 602;
        o_index_for_a4 <= 731;
        o_index_for_a5 <= 1021; 
    end
    877: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 0;
        o_index_for_a1 <= 326;
        o_index_for_a2 <= 438;
        o_index_for_a3 <= 603;
        o_index_for_a4 <= 732;
        o_index_for_a5 <= 1022; 
    end
    878: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 1;
        o_index_for_a1 <= 327;
        o_index_for_a2 <= 439;
        o_index_for_a3 <= 604;
        o_index_for_a4 <= 733;
        o_index_for_a5 <= 1023; 
    end
    879: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 2;
        o_index_for_a1 <= 328;
        o_index_for_a2 <= 440;
        o_index_for_a3 <= 605;
        o_index_for_a4 <= 734;
        o_index_for_a5 <= 1024; 
    end
    880: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 3;
        o_index_for_a1 <= 329;
        o_index_for_a2 <= 441;
        o_index_for_a3 <= 606;
        o_index_for_a4 <= 735;
        o_index_for_a5 <= 1025; 
    end
    881: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 4;
        o_index_for_a1 <= 330;
        o_index_for_a2 <= 442;
        o_index_for_a3 <= 607;
        o_index_for_a4 <= 736;
        o_index_for_a5 <= 1026; 
    end
    882: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 5;
        o_index_for_a1 <= 331;
        o_index_for_a2 <= 443;
        o_index_for_a3 <= 608;
        o_index_for_a4 <= 737;
        o_index_for_a5 <= 1027; 
    end
    883: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 6;
        o_index_for_a1 <= 332;
        o_index_for_a2 <= 444;
        o_index_for_a3 <= 609;
        o_index_for_a4 <= 738;
        o_index_for_a5 <= 1028; 
    end
    884: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 7;
        o_index_for_a1 <= 333;
        o_index_for_a2 <= 445;
        o_index_for_a3 <= 610;
        o_index_for_a4 <= 739;
        o_index_for_a5 <= 1029; 
    end
    885: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 8;
        o_index_for_a1 <= 334;
        o_index_for_a2 <= 446;
        o_index_for_a3 <= 611;
        o_index_for_a4 <= 740;
        o_index_for_a5 <= 1030; 
    end
    886: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 9;
        o_index_for_a1 <= 335;
        o_index_for_a2 <= 447;
        o_index_for_a3 <= 612;
        o_index_for_a4 <= 741;
        o_index_for_a5 <= 1031; 
    end
    887: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 10;
        o_index_for_a1 <= 336;
        o_index_for_a2 <= 448;
        o_index_for_a3 <= 613;
        o_index_for_a4 <= 742;
        o_index_for_a5 <= 1032; 
    end
    888: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 11;
        o_index_for_a1 <= 337;
        o_index_for_a2 <= 449;
        o_index_for_a3 <= 614;
        o_index_for_a4 <= 743;
        o_index_for_a5 <= 1033; 
    end
    889: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 12;
        o_index_for_a1 <= 338;
        o_index_for_a2 <= 450;
        o_index_for_a3 <= 615;
        o_index_for_a4 <= 744;
        o_index_for_a5 <= 1034; 
    end
    890: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 13;
        o_index_for_a1 <= 339;
        o_index_for_a2 <= 451;
        o_index_for_a3 <= 616;
        o_index_for_a4 <= 745;
        o_index_for_a5 <= 1035; 
    end
    891: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 14;
        o_index_for_a1 <= 340;
        o_index_for_a2 <= 452;
        o_index_for_a3 <= 617;
        o_index_for_a4 <= 746;
        o_index_for_a5 <= 1036; 
    end
    892: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 15;
        o_index_for_a1 <= 341;
        o_index_for_a2 <= 453;
        o_index_for_a3 <= 618;
        o_index_for_a4 <= 747;
        o_index_for_a5 <= 1037; 
    end
    893: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 16;
        o_index_for_a1 <= 342;
        o_index_for_a2 <= 454;
        o_index_for_a3 <= 619;
        o_index_for_a4 <= 748;
        o_index_for_a5 <= 1038; 
    end
    894: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 17;
        o_index_for_a1 <= 343;
        o_index_for_a2 <= 455;
        o_index_for_a3 <= 620;
        o_index_for_a4 <= 749;
        o_index_for_a5 <= 1039; 
    end
    895: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 18;
        o_index_for_a1 <= 344;
        o_index_for_a2 <= 456;
        o_index_for_a3 <= 621;
        o_index_for_a4 <= 750;
        o_index_for_a5 <= 1040; 
    end
    896: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 19;
        o_index_for_a1 <= 345;
        o_index_for_a2 <= 457;
        o_index_for_a3 <= 622;
        o_index_for_a4 <= 751;
        o_index_for_a5 <= 1041; 
    end
    897: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 20;
        o_index_for_a1 <= 346;
        o_index_for_a2 <= 458;
        o_index_for_a3 <= 623;
        o_index_for_a4 <= 752;
        o_index_for_a5 <= 1042; 
    end
    898: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 21;
        o_index_for_a1 <= 347;
        o_index_for_a2 <= 459;
        o_index_for_a3 <= 624;
        o_index_for_a4 <= 753;
        o_index_for_a5 <= 1043; 
    end
    899: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 22;
        o_index_for_a1 <= 348;
        o_index_for_a2 <= 460;
        o_index_for_a3 <= 625;
        o_index_for_a4 <= 754;
        o_index_for_a5 <= 1044; 
    end
    900: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 23;
        o_index_for_a1 <= 349;
        o_index_for_a2 <= 461;
        o_index_for_a3 <= 626;
        o_index_for_a4 <= 755;
        o_index_for_a5 <= 1045; 
    end
    901: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 24;
        o_index_for_a1 <= 350;
        o_index_for_a2 <= 462;
        o_index_for_a3 <= 627;
        o_index_for_a4 <= 756;
        o_index_for_a5 <= 1046; 
    end
    902: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 25;
        o_index_for_a1 <= 351;
        o_index_for_a2 <= 463;
        o_index_for_a3 <= 628;
        o_index_for_a4 <= 757;
        o_index_for_a5 <= 1047; 
    end
    903: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 26;
        o_index_for_a1 <= 352;
        o_index_for_a2 <= 464;
        o_index_for_a3 <= 629;
        o_index_for_a4 <= 758;
        o_index_for_a5 <= 1048; 
    end
    904: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 27;
        o_index_for_a1 <= 353;
        o_index_for_a2 <= 465;
        o_index_for_a3 <= 630;
        o_index_for_a4 <= 759;
        o_index_for_a5 <= 1049; 
    end
    905: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 28;
        o_index_for_a1 <= 354;
        o_index_for_a2 <= 466;
        o_index_for_a3 <= 631;
        o_index_for_a4 <= 760;
        o_index_for_a5 <= 1050; 
    end
    906: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 29;
        o_index_for_a1 <= 355;
        o_index_for_a2 <= 467;
        o_index_for_a3 <= 632;
        o_index_for_a4 <= 761;
        o_index_for_a5 <= 1051; 
    end
    907: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 30;
        o_index_for_a1 <= 356;
        o_index_for_a2 <= 468;
        o_index_for_a3 <= 633;
        o_index_for_a4 <= 762;
        o_index_for_a5 <= 1052; 
    end
    908: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 31;
        o_index_for_a1 <= 357;
        o_index_for_a2 <= 469;
        o_index_for_a3 <= 634;
        o_index_for_a4 <= 763;
        o_index_for_a5 <= 1053; 
    end
    909: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 32;
        o_index_for_a1 <= 358;
        o_index_for_a2 <= 470;
        o_index_for_a3 <= 635;
        o_index_for_a4 <= 764;
        o_index_for_a5 <= 1054; 
    end
    910: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 33;
        o_index_for_a1 <= 359;
        o_index_for_a2 <= 471;
        o_index_for_a3 <= 636;
        o_index_for_a4 <= 765;
        o_index_for_a5 <= 1055; 
    end
    911: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 34;
        o_index_for_a1 <= 360;
        o_index_for_a2 <= 472;
        o_index_for_a3 <= 637;
        o_index_for_a4 <= 766;
        o_index_for_a5 <= 960; 
    end
    912: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 35;
        o_index_for_a1 <= 361;
        o_index_for_a2 <= 473;
        o_index_for_a3 <= 638;
        o_index_for_a4 <= 767;
        o_index_for_a5 <= 961; 
    end
    913: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 36;
        o_index_for_a1 <= 362;
        o_index_for_a2 <= 474;
        o_index_for_a3 <= 639;
        o_index_for_a4 <= 672;
        o_index_for_a5 <= 962; 
    end
    914: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 37;
        o_index_for_a1 <= 363;
        o_index_for_a2 <= 475;
        o_index_for_a3 <= 640;
        o_index_for_a4 <= 673;
        o_index_for_a5 <= 963; 
    end
    915: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 38;
        o_index_for_a1 <= 364;
        o_index_for_a2 <= 476;
        o_index_for_a3 <= 641;
        o_index_for_a4 <= 674;
        o_index_for_a5 <= 964; 
    end
    916: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 39;
        o_index_for_a1 <= 365;
        o_index_for_a2 <= 477;
        o_index_for_a3 <= 642;
        o_index_for_a4 <= 675;
        o_index_for_a5 <= 965; 
    end
    917: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 40;
        o_index_for_a1 <= 366;
        o_index_for_a2 <= 478;
        o_index_for_a3 <= 643;
        o_index_for_a4 <= 676;
        o_index_for_a5 <= 966; 
    end
    918: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 41;
        o_index_for_a1 <= 367;
        o_index_for_a2 <= 479;
        o_index_for_a3 <= 644;
        o_index_for_a4 <= 677;
        o_index_for_a5 <= 967; 
    end
    919: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 42;
        o_index_for_a1 <= 368;
        o_index_for_a2 <= 384;
        o_index_for_a3 <= 645;
        o_index_for_a4 <= 678;
        o_index_for_a5 <= 968; 
    end
    920: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 43;
        o_index_for_a1 <= 369;
        o_index_for_a2 <= 385;
        o_index_for_a3 <= 646;
        o_index_for_a4 <= 679;
        o_index_for_a5 <= 969; 
    end
    921: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 44;
        o_index_for_a1 <= 370;
        o_index_for_a2 <= 386;
        o_index_for_a3 <= 647;
        o_index_for_a4 <= 680;
        o_index_for_a5 <= 970; 
    end
    922: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 45;
        o_index_for_a1 <= 371;
        o_index_for_a2 <= 387;
        o_index_for_a3 <= 648;
        o_index_for_a4 <= 681;
        o_index_for_a5 <= 971; 
    end
    923: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 46;
        o_index_for_a1 <= 372;
        o_index_for_a2 <= 388;
        o_index_for_a3 <= 649;
        o_index_for_a4 <= 682;
        o_index_for_a5 <= 972; 
    end
    924: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 47;
        o_index_for_a1 <= 373;
        o_index_for_a2 <= 389;
        o_index_for_a3 <= 650;
        o_index_for_a4 <= 683;
        o_index_for_a5 <= 973; 
    end
    925: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 48;
        o_index_for_a1 <= 374;
        o_index_for_a2 <= 390;
        o_index_for_a3 <= 651;
        o_index_for_a4 <= 684;
        o_index_for_a5 <= 974; 
    end
    926: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 49;
        o_index_for_a1 <= 375;
        o_index_for_a2 <= 391;
        o_index_for_a3 <= 652;
        o_index_for_a4 <= 685;
        o_index_for_a5 <= 975; 
    end
    927: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 50;
        o_index_for_a1 <= 376;
        o_index_for_a2 <= 392;
        o_index_for_a3 <= 653;
        o_index_for_a4 <= 686;
        o_index_for_a5 <= 976; 
    end
    928: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 51;
        o_index_for_a1 <= 377;
        o_index_for_a2 <= 393;
        o_index_for_a3 <= 654;
        o_index_for_a4 <= 687;
        o_index_for_a5 <= 977; 
    end
    929: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 52;
        o_index_for_a1 <= 378;
        o_index_for_a2 <= 394;
        o_index_for_a3 <= 655;
        o_index_for_a4 <= 688;
        o_index_for_a5 <= 978; 
    end
    930: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 53;
        o_index_for_a1 <= 379;
        o_index_for_a2 <= 395;
        o_index_for_a3 <= 656;
        o_index_for_a4 <= 689;
        o_index_for_a5 <= 979; 
    end
    931: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 54;
        o_index_for_a1 <= 380;
        o_index_for_a2 <= 396;
        o_index_for_a3 <= 657;
        o_index_for_a4 <= 690;
        o_index_for_a5 <= 980; 
    end
    932: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 55;
        o_index_for_a1 <= 381;
        o_index_for_a2 <= 397;
        o_index_for_a3 <= 658;
        o_index_for_a4 <= 691;
        o_index_for_a5 <= 981; 
    end
    933: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 56;
        o_index_for_a1 <= 382;
        o_index_for_a2 <= 398;
        o_index_for_a3 <= 659;
        o_index_for_a4 <= 692;
        o_index_for_a5 <= 982; 
    end
    934: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 57;
        o_index_for_a1 <= 383;
        o_index_for_a2 <= 399;
        o_index_for_a3 <= 660;
        o_index_for_a4 <= 693;
        o_index_for_a5 <= 983; 
    end
    935: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 58;
        o_index_for_a1 <= 288;
        o_index_for_a2 <= 400;
        o_index_for_a3 <= 661;
        o_index_for_a4 <= 694;
        o_index_for_a5 <= 984; 
    end
    936: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 59;
        o_index_for_a1 <= 289;
        o_index_for_a2 <= 401;
        o_index_for_a3 <= 662;
        o_index_for_a4 <= 695;
        o_index_for_a5 <= 985; 
    end
    937: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 60;
        o_index_for_a1 <= 290;
        o_index_for_a2 <= 402;
        o_index_for_a3 <= 663;
        o_index_for_a4 <= 696;
        o_index_for_a5 <= 986; 
    end
    938: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 61;
        o_index_for_a1 <= 291;
        o_index_for_a2 <= 403;
        o_index_for_a3 <= 664;
        o_index_for_a4 <= 697;
        o_index_for_a5 <= 987; 
    end
    939: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 62;
        o_index_for_a1 <= 292;
        o_index_for_a2 <= 404;
        o_index_for_a3 <= 665;
        o_index_for_a4 <= 698;
        o_index_for_a5 <= 988; 
    end
    940: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 63;
        o_index_for_a1 <= 293;
        o_index_for_a2 <= 405;
        o_index_for_a3 <= 666;
        o_index_for_a4 <= 699;
        o_index_for_a5 <= 989; 
    end
    941: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 64;
        o_index_for_a1 <= 294;
        o_index_for_a2 <= 406;
        o_index_for_a3 <= 667;
        o_index_for_a4 <= 700;
        o_index_for_a5 <= 990; 
    end
    942: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 65;
        o_index_for_a1 <= 295;
        o_index_for_a2 <= 407;
        o_index_for_a3 <= 668;
        o_index_for_a4 <= 701;
        o_index_for_a5 <= 991; 
    end
    943: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 66;
        o_index_for_a1 <= 296;
        o_index_for_a2 <= 408;
        o_index_for_a3 <= 669;
        o_index_for_a4 <= 702;
        o_index_for_a5 <= 992; 
    end
    944: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 67;
        o_index_for_a1 <= 297;
        o_index_for_a2 <= 409;
        o_index_for_a3 <= 670;
        o_index_for_a4 <= 703;
        o_index_for_a5 <= 993; 
    end
    945: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 68;
        o_index_for_a1 <= 298;
        o_index_for_a2 <= 410;
        o_index_for_a3 <= 671;
        o_index_for_a4 <= 704;
        o_index_for_a5 <= 994; 
    end
    946: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 69;
        o_index_for_a1 <= 299;
        o_index_for_a2 <= 411;
        o_index_for_a3 <= 576;
        o_index_for_a4 <= 705;
        o_index_for_a5 <= 995; 
    end
    947: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 70;
        o_index_for_a1 <= 300;
        o_index_for_a2 <= 412;
        o_index_for_a3 <= 577;
        o_index_for_a4 <= 706;
        o_index_for_a5 <= 996; 
    end
    948: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 71;
        o_index_for_a1 <= 301;
        o_index_for_a2 <= 413;
        o_index_for_a3 <= 578;
        o_index_for_a4 <= 707;
        o_index_for_a5 <= 997; 
    end
    949: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 72;
        o_index_for_a1 <= 302;
        o_index_for_a2 <= 414;
        o_index_for_a3 <= 579;
        o_index_for_a4 <= 708;
        o_index_for_a5 <= 998; 
    end
    950: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 73;
        o_index_for_a1 <= 303;
        o_index_for_a2 <= 415;
        o_index_for_a3 <= 580;
        o_index_for_a4 <= 709;
        o_index_for_a5 <= 999; 
    end
    951: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 74;
        o_index_for_a1 <= 304;
        o_index_for_a2 <= 416;
        o_index_for_a3 <= 581;
        o_index_for_a4 <= 710;
        o_index_for_a5 <= 1000; 
    end
    952: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 75;
        o_index_for_a1 <= 305;
        o_index_for_a2 <= 417;
        o_index_for_a3 <= 582;
        o_index_for_a4 <= 711;
        o_index_for_a5 <= 1001; 
    end
    953: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 76;
        o_index_for_a1 <= 306;
        o_index_for_a2 <= 418;
        o_index_for_a3 <= 583;
        o_index_for_a4 <= 712;
        o_index_for_a5 <= 1002; 
    end
    954: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 77;
        o_index_for_a1 <= 307;
        o_index_for_a2 <= 419;
        o_index_for_a3 <= 584;
        o_index_for_a4 <= 713;
        o_index_for_a5 <= 1003; 
    end
    955: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 78;
        o_index_for_a1 <= 308;
        o_index_for_a2 <= 420;
        o_index_for_a3 <= 585;
        o_index_for_a4 <= 714;
        o_index_for_a5 <= 1004; 
    end
    956: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 79;
        o_index_for_a1 <= 309;
        o_index_for_a2 <= 421;
        o_index_for_a3 <= 586;
        o_index_for_a4 <= 715;
        o_index_for_a5 <= 1005; 
    end
    957: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 80;
        o_index_for_a1 <= 310;
        o_index_for_a2 <= 422;
        o_index_for_a3 <= 587;
        o_index_for_a4 <= 716;
        o_index_for_a5 <= 1006; 
    end
    958: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 81;
        o_index_for_a1 <= 311;
        o_index_for_a2 <= 423;
        o_index_for_a3 <= 588;
        o_index_for_a4 <= 717;
        o_index_for_a5 <= 1007; 
    end
    959: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 82;
        o_index_for_a1 <= 312;
        o_index_for_a2 <= 424;
        o_index_for_a3 <= 589;
        o_index_for_a4 <= 718;
        o_index_for_a5 <= 1008; 
    end
    960: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 456;
        o_index_for_a1 <= 594;
        o_index_for_a2 <= 934;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    961: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 457;
        o_index_for_a1 <= 595;
        o_index_for_a2 <= 935;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    962: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 458;
        o_index_for_a1 <= 596;
        o_index_for_a2 <= 936;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    963: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 459;
        o_index_for_a1 <= 597;
        o_index_for_a2 <= 937;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    964: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 460;
        o_index_for_a1 <= 598;
        o_index_for_a2 <= 938;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    965: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 461;
        o_index_for_a1 <= 599;
        o_index_for_a2 <= 939;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    966: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 462;
        o_index_for_a1 <= 600;
        o_index_for_a2 <= 940;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    967: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 463;
        o_index_for_a1 <= 601;
        o_index_for_a2 <= 941;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    968: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 464;
        o_index_for_a1 <= 602;
        o_index_for_a2 <= 942;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    969: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 465;
        o_index_for_a1 <= 603;
        o_index_for_a2 <= 943;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    970: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 466;
        o_index_for_a1 <= 604;
        o_index_for_a2 <= 944;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    971: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 467;
        o_index_for_a1 <= 605;
        o_index_for_a2 <= 945;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    972: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 468;
        o_index_for_a1 <= 606;
        o_index_for_a2 <= 946;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    973: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 469;
        o_index_for_a1 <= 607;
        o_index_for_a2 <= 947;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    974: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 470;
        o_index_for_a1 <= 608;
        o_index_for_a2 <= 948;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    975: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 471;
        o_index_for_a1 <= 609;
        o_index_for_a2 <= 949;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    976: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 472;
        o_index_for_a1 <= 610;
        o_index_for_a2 <= 950;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    977: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 473;
        o_index_for_a1 <= 611;
        o_index_for_a2 <= 951;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    978: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 474;
        o_index_for_a1 <= 612;
        o_index_for_a2 <= 952;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    979: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 475;
        o_index_for_a1 <= 613;
        o_index_for_a2 <= 953;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    980: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 476;
        o_index_for_a1 <= 614;
        o_index_for_a2 <= 954;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    981: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 477;
        o_index_for_a1 <= 615;
        o_index_for_a2 <= 955;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    982: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 478;
        o_index_for_a1 <= 616;
        o_index_for_a2 <= 956;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    983: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 479;
        o_index_for_a1 <= 617;
        o_index_for_a2 <= 957;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    984: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 384;
        o_index_for_a1 <= 618;
        o_index_for_a2 <= 958;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    985: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 385;
        o_index_for_a1 <= 619;
        o_index_for_a2 <= 959;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    986: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 386;
        o_index_for_a1 <= 620;
        o_index_for_a2 <= 864;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    987: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 387;
        o_index_for_a1 <= 621;
        o_index_for_a2 <= 865;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    988: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 388;
        o_index_for_a1 <= 622;
        o_index_for_a2 <= 866;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    989: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 389;
        o_index_for_a1 <= 623;
        o_index_for_a2 <= 867;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    990: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 390;
        o_index_for_a1 <= 624;
        o_index_for_a2 <= 868;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    991: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 391;
        o_index_for_a1 <= 625;
        o_index_for_a2 <= 869;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    992: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 392;
        o_index_for_a1 <= 626;
        o_index_for_a2 <= 870;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    993: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 393;
        o_index_for_a1 <= 627;
        o_index_for_a2 <= 871;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    994: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 394;
        o_index_for_a1 <= 628;
        o_index_for_a2 <= 872;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    995: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 395;
        o_index_for_a1 <= 629;
        o_index_for_a2 <= 873;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    996: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 396;
        o_index_for_a1 <= 630;
        o_index_for_a2 <= 874;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    997: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 397;
        o_index_for_a1 <= 631;
        o_index_for_a2 <= 875;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    998: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 398;
        o_index_for_a1 <= 632;
        o_index_for_a2 <= 876;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    999: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 399;
        o_index_for_a1 <= 633;
        o_index_for_a2 <= 877;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1000: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 400;
        o_index_for_a1 <= 634;
        o_index_for_a2 <= 878;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1001: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 401;
        o_index_for_a1 <= 635;
        o_index_for_a2 <= 879;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1002: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 402;
        o_index_for_a1 <= 636;
        o_index_for_a2 <= 880;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1003: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 403;
        o_index_for_a1 <= 637;
        o_index_for_a2 <= 881;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1004: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 404;
        o_index_for_a1 <= 638;
        o_index_for_a2 <= 882;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1005: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 405;
        o_index_for_a1 <= 639;
        o_index_for_a2 <= 883;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1006: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 406;
        o_index_for_a1 <= 640;
        o_index_for_a2 <= 884;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1007: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 407;
        o_index_for_a1 <= 641;
        o_index_for_a2 <= 885;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1008: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 408;
        o_index_for_a1 <= 642;
        o_index_for_a2 <= 886;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1009: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 409;
        o_index_for_a1 <= 643;
        o_index_for_a2 <= 887;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1010: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 410;
        o_index_for_a1 <= 644;
        o_index_for_a2 <= 888;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1011: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 411;
        o_index_for_a1 <= 645;
        o_index_for_a2 <= 889;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1012: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 412;
        o_index_for_a1 <= 646;
        o_index_for_a2 <= 890;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1013: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 413;
        o_index_for_a1 <= 647;
        o_index_for_a2 <= 891;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1014: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 414;
        o_index_for_a1 <= 648;
        o_index_for_a2 <= 892;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1015: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 415;
        o_index_for_a1 <= 649;
        o_index_for_a2 <= 893;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1016: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 416;
        o_index_for_a1 <= 650;
        o_index_for_a2 <= 894;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1017: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 417;
        o_index_for_a1 <= 651;
        o_index_for_a2 <= 895;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1018: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 418;
        o_index_for_a1 <= 652;
        o_index_for_a2 <= 896;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1019: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 419;
        o_index_for_a1 <= 653;
        o_index_for_a2 <= 897;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1020: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 420;
        o_index_for_a1 <= 654;
        o_index_for_a2 <= 898;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1021: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 421;
        o_index_for_a1 <= 655;
        o_index_for_a2 <= 899;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1022: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 422;
        o_index_for_a1 <= 656;
        o_index_for_a2 <= 900;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1023: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 423;
        o_index_for_a1 <= 657;
        o_index_for_a2 <= 901;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1024: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 424;
        o_index_for_a1 <= 658;
        o_index_for_a2 <= 902;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1025: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 425;
        o_index_for_a1 <= 659;
        o_index_for_a2 <= 903;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1026: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 426;
        o_index_for_a1 <= 660;
        o_index_for_a2 <= 904;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1027: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 427;
        o_index_for_a1 <= 661;
        o_index_for_a2 <= 905;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1028: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 428;
        o_index_for_a1 <= 662;
        o_index_for_a2 <= 906;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1029: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 429;
        o_index_for_a1 <= 663;
        o_index_for_a2 <= 907;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1030: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 430;
        o_index_for_a1 <= 664;
        o_index_for_a2 <= 908;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1031: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 431;
        o_index_for_a1 <= 665;
        o_index_for_a2 <= 909;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1032: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 432;
        o_index_for_a1 <= 666;
        o_index_for_a2 <= 910;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1033: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 433;
        o_index_for_a1 <= 667;
        o_index_for_a2 <= 911;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1034: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 434;
        o_index_for_a1 <= 668;
        o_index_for_a2 <= 912;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1035: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 435;
        o_index_for_a1 <= 669;
        o_index_for_a2 <= 913;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1036: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 436;
        o_index_for_a1 <= 670;
        o_index_for_a2 <= 914;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1037: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 437;
        o_index_for_a1 <= 671;
        o_index_for_a2 <= 915;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1038: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 438;
        o_index_for_a1 <= 576;
        o_index_for_a2 <= 916;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1039: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 439;
        o_index_for_a1 <= 577;
        o_index_for_a2 <= 917;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1040: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 440;
        o_index_for_a1 <= 578;
        o_index_for_a2 <= 918;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1041: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 441;
        o_index_for_a1 <= 579;
        o_index_for_a2 <= 919;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1042: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 442;
        o_index_for_a1 <= 580;
        o_index_for_a2 <= 920;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1043: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 443;
        o_index_for_a1 <= 581;
        o_index_for_a2 <= 921;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1044: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 444;
        o_index_for_a1 <= 582;
        o_index_for_a2 <= 922;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1045: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 445;
        o_index_for_a1 <= 583;
        o_index_for_a2 <= 923;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1046: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 446;
        o_index_for_a1 <= 584;
        o_index_for_a2 <= 924;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1047: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 447;
        o_index_for_a1 <= 585;
        o_index_for_a2 <= 925;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1048: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 448;
        o_index_for_a1 <= 586;
        o_index_for_a2 <= 926;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1049: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 449;
        o_index_for_a1 <= 587;
        o_index_for_a2 <= 927;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1050: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 450;
        o_index_for_a1 <= 588;
        o_index_for_a2 <= 928;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1051: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 451;
        o_index_for_a1 <= 589;
        o_index_for_a2 <= 929;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1052: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 452;
        o_index_for_a1 <= 590;
        o_index_for_a2 <= 930;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1053: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 453;
        o_index_for_a1 <= 591;
        o_index_for_a2 <= 931;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1054: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 454;
        o_index_for_a1 <= 592;
        o_index_for_a2 <= 932;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1055: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 3;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 455;
        o_index_for_a1 <= 593;
        o_index_for_a2 <= 933;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1056: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 108;
        o_index_for_a1 <= 192;
        o_index_for_a2 <= 559;
        o_index_for_a3 <= 819;
        o_index_for_a4 <= 936;
        o_index_for_a5 <= 1082; 
    end
    1057: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 109;
        o_index_for_a1 <= 193;
        o_index_for_a2 <= 560;
        o_index_for_a3 <= 820;
        o_index_for_a4 <= 937;
        o_index_for_a5 <= 1083; 
    end
    1058: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 110;
        o_index_for_a1 <= 194;
        o_index_for_a2 <= 561;
        o_index_for_a3 <= 821;
        o_index_for_a4 <= 938;
        o_index_for_a5 <= 1084; 
    end
    1059: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 111;
        o_index_for_a1 <= 195;
        o_index_for_a2 <= 562;
        o_index_for_a3 <= 822;
        o_index_for_a4 <= 939;
        o_index_for_a5 <= 1085; 
    end
    1060: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 112;
        o_index_for_a1 <= 196;
        o_index_for_a2 <= 563;
        o_index_for_a3 <= 823;
        o_index_for_a4 <= 940;
        o_index_for_a5 <= 1086; 
    end
    1061: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 113;
        o_index_for_a1 <= 197;
        o_index_for_a2 <= 564;
        o_index_for_a3 <= 824;
        o_index_for_a4 <= 941;
        o_index_for_a5 <= 1087; 
    end
    1062: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 114;
        o_index_for_a1 <= 198;
        o_index_for_a2 <= 565;
        o_index_for_a3 <= 825;
        o_index_for_a4 <= 942;
        o_index_for_a5 <= 1088; 
    end
    1063: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 115;
        o_index_for_a1 <= 199;
        o_index_for_a2 <= 566;
        o_index_for_a3 <= 826;
        o_index_for_a4 <= 943;
        o_index_for_a5 <= 1089; 
    end
    1064: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 116;
        o_index_for_a1 <= 200;
        o_index_for_a2 <= 567;
        o_index_for_a3 <= 827;
        o_index_for_a4 <= 944;
        o_index_for_a5 <= 1090; 
    end
    1065: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 117;
        o_index_for_a1 <= 201;
        o_index_for_a2 <= 568;
        o_index_for_a3 <= 828;
        o_index_for_a4 <= 945;
        o_index_for_a5 <= 1091; 
    end
    1066: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 118;
        o_index_for_a1 <= 202;
        o_index_for_a2 <= 569;
        o_index_for_a3 <= 829;
        o_index_for_a4 <= 946;
        o_index_for_a5 <= 1092; 
    end
    1067: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 119;
        o_index_for_a1 <= 203;
        o_index_for_a2 <= 570;
        o_index_for_a3 <= 830;
        o_index_for_a4 <= 947;
        o_index_for_a5 <= 1093; 
    end
    1068: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 120;
        o_index_for_a1 <= 204;
        o_index_for_a2 <= 571;
        o_index_for_a3 <= 831;
        o_index_for_a4 <= 948;
        o_index_for_a5 <= 1094; 
    end
    1069: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 121;
        o_index_for_a1 <= 205;
        o_index_for_a2 <= 572;
        o_index_for_a3 <= 832;
        o_index_for_a4 <= 949;
        o_index_for_a5 <= 1095; 
    end
    1070: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 122;
        o_index_for_a1 <= 206;
        o_index_for_a2 <= 573;
        o_index_for_a3 <= 833;
        o_index_for_a4 <= 950;
        o_index_for_a5 <= 1096; 
    end
    1071: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 123;
        o_index_for_a1 <= 207;
        o_index_for_a2 <= 574;
        o_index_for_a3 <= 834;
        o_index_for_a4 <= 951;
        o_index_for_a5 <= 1097; 
    end
    1072: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 124;
        o_index_for_a1 <= 208;
        o_index_for_a2 <= 575;
        o_index_for_a3 <= 835;
        o_index_for_a4 <= 952;
        o_index_for_a5 <= 1098; 
    end
    1073: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 125;
        o_index_for_a1 <= 209;
        o_index_for_a2 <= 480;
        o_index_for_a3 <= 836;
        o_index_for_a4 <= 953;
        o_index_for_a5 <= 1099; 
    end
    1074: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 126;
        o_index_for_a1 <= 210;
        o_index_for_a2 <= 481;
        o_index_for_a3 <= 837;
        o_index_for_a4 <= 954;
        o_index_for_a5 <= 1100; 
    end
    1075: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 127;
        o_index_for_a1 <= 211;
        o_index_for_a2 <= 482;
        o_index_for_a3 <= 838;
        o_index_for_a4 <= 955;
        o_index_for_a5 <= 1101; 
    end
    1076: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 128;
        o_index_for_a1 <= 212;
        o_index_for_a2 <= 483;
        o_index_for_a3 <= 839;
        o_index_for_a4 <= 956;
        o_index_for_a5 <= 1102; 
    end
    1077: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 129;
        o_index_for_a1 <= 213;
        o_index_for_a2 <= 484;
        o_index_for_a3 <= 840;
        o_index_for_a4 <= 957;
        o_index_for_a5 <= 1103; 
    end
    1078: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 130;
        o_index_for_a1 <= 214;
        o_index_for_a2 <= 485;
        o_index_for_a3 <= 841;
        o_index_for_a4 <= 958;
        o_index_for_a5 <= 1104; 
    end
    1079: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 131;
        o_index_for_a1 <= 215;
        o_index_for_a2 <= 486;
        o_index_for_a3 <= 842;
        o_index_for_a4 <= 959;
        o_index_for_a5 <= 1105; 
    end
    1080: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 132;
        o_index_for_a1 <= 216;
        o_index_for_a2 <= 487;
        o_index_for_a3 <= 843;
        o_index_for_a4 <= 864;
        o_index_for_a5 <= 1106; 
    end
    1081: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 133;
        o_index_for_a1 <= 217;
        o_index_for_a2 <= 488;
        o_index_for_a3 <= 844;
        o_index_for_a4 <= 865;
        o_index_for_a5 <= 1107; 
    end
    1082: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 134;
        o_index_for_a1 <= 218;
        o_index_for_a2 <= 489;
        o_index_for_a3 <= 845;
        o_index_for_a4 <= 866;
        o_index_for_a5 <= 1108; 
    end
    1083: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 135;
        o_index_for_a1 <= 219;
        o_index_for_a2 <= 490;
        o_index_for_a3 <= 846;
        o_index_for_a4 <= 867;
        o_index_for_a5 <= 1109; 
    end
    1084: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 136;
        o_index_for_a1 <= 220;
        o_index_for_a2 <= 491;
        o_index_for_a3 <= 847;
        o_index_for_a4 <= 868;
        o_index_for_a5 <= 1110; 
    end
    1085: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 137;
        o_index_for_a1 <= 221;
        o_index_for_a2 <= 492;
        o_index_for_a3 <= 848;
        o_index_for_a4 <= 869;
        o_index_for_a5 <= 1111; 
    end
    1086: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 138;
        o_index_for_a1 <= 222;
        o_index_for_a2 <= 493;
        o_index_for_a3 <= 849;
        o_index_for_a4 <= 870;
        o_index_for_a5 <= 1112; 
    end
    1087: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 139;
        o_index_for_a1 <= 223;
        o_index_for_a2 <= 494;
        o_index_for_a3 <= 850;
        o_index_for_a4 <= 871;
        o_index_for_a5 <= 1113; 
    end
    1088: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 140;
        o_index_for_a1 <= 224;
        o_index_for_a2 <= 495;
        o_index_for_a3 <= 851;
        o_index_for_a4 <= 872;
        o_index_for_a5 <= 1114; 
    end
    1089: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 141;
        o_index_for_a1 <= 225;
        o_index_for_a2 <= 496;
        o_index_for_a3 <= 852;
        o_index_for_a4 <= 873;
        o_index_for_a5 <= 1115; 
    end
    1090: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 142;
        o_index_for_a1 <= 226;
        o_index_for_a2 <= 497;
        o_index_for_a3 <= 853;
        o_index_for_a4 <= 874;
        o_index_for_a5 <= 1116; 
    end
    1091: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 143;
        o_index_for_a1 <= 227;
        o_index_for_a2 <= 498;
        o_index_for_a3 <= 854;
        o_index_for_a4 <= 875;
        o_index_for_a5 <= 1117; 
    end
    1092: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 144;
        o_index_for_a1 <= 228;
        o_index_for_a2 <= 499;
        o_index_for_a3 <= 855;
        o_index_for_a4 <= 876;
        o_index_for_a5 <= 1118; 
    end
    1093: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 145;
        o_index_for_a1 <= 229;
        o_index_for_a2 <= 500;
        o_index_for_a3 <= 856;
        o_index_for_a4 <= 877;
        o_index_for_a5 <= 1119; 
    end
    1094: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 146;
        o_index_for_a1 <= 230;
        o_index_for_a2 <= 501;
        o_index_for_a3 <= 857;
        o_index_for_a4 <= 878;
        o_index_for_a5 <= 1120; 
    end
    1095: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 147;
        o_index_for_a1 <= 231;
        o_index_for_a2 <= 502;
        o_index_for_a3 <= 858;
        o_index_for_a4 <= 879;
        o_index_for_a5 <= 1121; 
    end
    1096: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 148;
        o_index_for_a1 <= 232;
        o_index_for_a2 <= 503;
        o_index_for_a3 <= 859;
        o_index_for_a4 <= 880;
        o_index_for_a5 <= 1122; 
    end
    1097: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 149;
        o_index_for_a1 <= 233;
        o_index_for_a2 <= 504;
        o_index_for_a3 <= 860;
        o_index_for_a4 <= 881;
        o_index_for_a5 <= 1123; 
    end
    1098: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 150;
        o_index_for_a1 <= 234;
        o_index_for_a2 <= 505;
        o_index_for_a3 <= 861;
        o_index_for_a4 <= 882;
        o_index_for_a5 <= 1124; 
    end
    1099: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 151;
        o_index_for_a1 <= 235;
        o_index_for_a2 <= 506;
        o_index_for_a3 <= 862;
        o_index_for_a4 <= 883;
        o_index_for_a5 <= 1125; 
    end
    1100: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 152;
        o_index_for_a1 <= 236;
        o_index_for_a2 <= 507;
        o_index_for_a3 <= 863;
        o_index_for_a4 <= 884;
        o_index_for_a5 <= 1126; 
    end
    1101: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 153;
        o_index_for_a1 <= 237;
        o_index_for_a2 <= 508;
        o_index_for_a3 <= 768;
        o_index_for_a4 <= 885;
        o_index_for_a5 <= 1127; 
    end
    1102: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 154;
        o_index_for_a1 <= 238;
        o_index_for_a2 <= 509;
        o_index_for_a3 <= 769;
        o_index_for_a4 <= 886;
        o_index_for_a5 <= 1128; 
    end
    1103: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 155;
        o_index_for_a1 <= 239;
        o_index_for_a2 <= 510;
        o_index_for_a3 <= 770;
        o_index_for_a4 <= 887;
        o_index_for_a5 <= 1129; 
    end
    1104: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 156;
        o_index_for_a1 <= 240;
        o_index_for_a2 <= 511;
        o_index_for_a3 <= 771;
        o_index_for_a4 <= 888;
        o_index_for_a5 <= 1130; 
    end
    1105: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 157;
        o_index_for_a1 <= 241;
        o_index_for_a2 <= 512;
        o_index_for_a3 <= 772;
        o_index_for_a4 <= 889;
        o_index_for_a5 <= 1131; 
    end
    1106: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 158;
        o_index_for_a1 <= 242;
        o_index_for_a2 <= 513;
        o_index_for_a3 <= 773;
        o_index_for_a4 <= 890;
        o_index_for_a5 <= 1132; 
    end
    1107: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 159;
        o_index_for_a1 <= 243;
        o_index_for_a2 <= 514;
        o_index_for_a3 <= 774;
        o_index_for_a4 <= 891;
        o_index_for_a5 <= 1133; 
    end
    1108: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 160;
        o_index_for_a1 <= 244;
        o_index_for_a2 <= 515;
        o_index_for_a3 <= 775;
        o_index_for_a4 <= 892;
        o_index_for_a5 <= 1134; 
    end
    1109: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 161;
        o_index_for_a1 <= 245;
        o_index_for_a2 <= 516;
        o_index_for_a3 <= 776;
        o_index_for_a4 <= 893;
        o_index_for_a5 <= 1135; 
    end
    1110: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 162;
        o_index_for_a1 <= 246;
        o_index_for_a2 <= 517;
        o_index_for_a3 <= 777;
        o_index_for_a4 <= 894;
        o_index_for_a5 <= 1136; 
    end
    1111: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 163;
        o_index_for_a1 <= 247;
        o_index_for_a2 <= 518;
        o_index_for_a3 <= 778;
        o_index_for_a4 <= 895;
        o_index_for_a5 <= 1137; 
    end
    1112: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 164;
        o_index_for_a1 <= 248;
        o_index_for_a2 <= 519;
        o_index_for_a3 <= 779;
        o_index_for_a4 <= 896;
        o_index_for_a5 <= 1138; 
    end
    1113: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 165;
        o_index_for_a1 <= 249;
        o_index_for_a2 <= 520;
        o_index_for_a3 <= 780;
        o_index_for_a4 <= 897;
        o_index_for_a5 <= 1139; 
    end
    1114: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 166;
        o_index_for_a1 <= 250;
        o_index_for_a2 <= 521;
        o_index_for_a3 <= 781;
        o_index_for_a4 <= 898;
        o_index_for_a5 <= 1140; 
    end
    1115: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 167;
        o_index_for_a1 <= 251;
        o_index_for_a2 <= 522;
        o_index_for_a3 <= 782;
        o_index_for_a4 <= 899;
        o_index_for_a5 <= 1141; 
    end
    1116: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 168;
        o_index_for_a1 <= 252;
        o_index_for_a2 <= 523;
        o_index_for_a3 <= 783;
        o_index_for_a4 <= 900;
        o_index_for_a5 <= 1142; 
    end
    1117: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 169;
        o_index_for_a1 <= 253;
        o_index_for_a2 <= 524;
        o_index_for_a3 <= 784;
        o_index_for_a4 <= 901;
        o_index_for_a5 <= 1143; 
    end
    1118: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 170;
        o_index_for_a1 <= 254;
        o_index_for_a2 <= 525;
        o_index_for_a3 <= 785;
        o_index_for_a4 <= 902;
        o_index_for_a5 <= 1144; 
    end
    1119: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 171;
        o_index_for_a1 <= 255;
        o_index_for_a2 <= 526;
        o_index_for_a3 <= 786;
        o_index_for_a4 <= 903;
        o_index_for_a5 <= 1145; 
    end
    1120: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 172;
        o_index_for_a1 <= 256;
        o_index_for_a2 <= 527;
        o_index_for_a3 <= 787;
        o_index_for_a4 <= 904;
        o_index_for_a5 <= 1146; 
    end
    1121: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 173;
        o_index_for_a1 <= 257;
        o_index_for_a2 <= 528;
        o_index_for_a3 <= 788;
        o_index_for_a4 <= 905;
        o_index_for_a5 <= 1147; 
    end
    1122: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 174;
        o_index_for_a1 <= 258;
        o_index_for_a2 <= 529;
        o_index_for_a3 <= 789;
        o_index_for_a4 <= 906;
        o_index_for_a5 <= 1148; 
    end
    1123: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 175;
        o_index_for_a1 <= 259;
        o_index_for_a2 <= 530;
        o_index_for_a3 <= 790;
        o_index_for_a4 <= 907;
        o_index_for_a5 <= 1149; 
    end
    1124: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 176;
        o_index_for_a1 <= 260;
        o_index_for_a2 <= 531;
        o_index_for_a3 <= 791;
        o_index_for_a4 <= 908;
        o_index_for_a5 <= 1150; 
    end
    1125: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 177;
        o_index_for_a1 <= 261;
        o_index_for_a2 <= 532;
        o_index_for_a3 <= 792;
        o_index_for_a4 <= 909;
        o_index_for_a5 <= 1151; 
    end
    1126: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 178;
        o_index_for_a1 <= 262;
        o_index_for_a2 <= 533;
        o_index_for_a3 <= 793;
        o_index_for_a4 <= 910;
        o_index_for_a5 <= 1056; 
    end
    1127: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 179;
        o_index_for_a1 <= 263;
        o_index_for_a2 <= 534;
        o_index_for_a3 <= 794;
        o_index_for_a4 <= 911;
        o_index_for_a5 <= 1057; 
    end
    1128: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 180;
        o_index_for_a1 <= 264;
        o_index_for_a2 <= 535;
        o_index_for_a3 <= 795;
        o_index_for_a4 <= 912;
        o_index_for_a5 <= 1058; 
    end
    1129: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 181;
        o_index_for_a1 <= 265;
        o_index_for_a2 <= 536;
        o_index_for_a3 <= 796;
        o_index_for_a4 <= 913;
        o_index_for_a5 <= 1059; 
    end
    1130: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 182;
        o_index_for_a1 <= 266;
        o_index_for_a2 <= 537;
        o_index_for_a3 <= 797;
        o_index_for_a4 <= 914;
        o_index_for_a5 <= 1060; 
    end
    1131: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 183;
        o_index_for_a1 <= 267;
        o_index_for_a2 <= 538;
        o_index_for_a3 <= 798;
        o_index_for_a4 <= 915;
        o_index_for_a5 <= 1061; 
    end
    1132: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 184;
        o_index_for_a1 <= 268;
        o_index_for_a2 <= 539;
        o_index_for_a3 <= 799;
        o_index_for_a4 <= 916;
        o_index_for_a5 <= 1062; 
    end
    1133: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 185;
        o_index_for_a1 <= 269;
        o_index_for_a2 <= 540;
        o_index_for_a3 <= 800;
        o_index_for_a4 <= 917;
        o_index_for_a5 <= 1063; 
    end
    1134: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 186;
        o_index_for_a1 <= 270;
        o_index_for_a2 <= 541;
        o_index_for_a3 <= 801;
        o_index_for_a4 <= 918;
        o_index_for_a5 <= 1064; 
    end
    1135: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 187;
        o_index_for_a1 <= 271;
        o_index_for_a2 <= 542;
        o_index_for_a3 <= 802;
        o_index_for_a4 <= 919;
        o_index_for_a5 <= 1065; 
    end
    1136: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 188;
        o_index_for_a1 <= 272;
        o_index_for_a2 <= 543;
        o_index_for_a3 <= 803;
        o_index_for_a4 <= 920;
        o_index_for_a5 <= 1066; 
    end
    1137: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 189;
        o_index_for_a1 <= 273;
        o_index_for_a2 <= 544;
        o_index_for_a3 <= 804;
        o_index_for_a4 <= 921;
        o_index_for_a5 <= 1067; 
    end
    1138: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 190;
        o_index_for_a1 <= 274;
        o_index_for_a2 <= 545;
        o_index_for_a3 <= 805;
        o_index_for_a4 <= 922;
        o_index_for_a5 <= 1068; 
    end
    1139: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 191;
        o_index_for_a1 <= 275;
        o_index_for_a2 <= 546;
        o_index_for_a3 <= 806;
        o_index_for_a4 <= 923;
        o_index_for_a5 <= 1069; 
    end
    1140: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 96;
        o_index_for_a1 <= 276;
        o_index_for_a2 <= 547;
        o_index_for_a3 <= 807;
        o_index_for_a4 <= 924;
        o_index_for_a5 <= 1070; 
    end
    1141: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 97;
        o_index_for_a1 <= 277;
        o_index_for_a2 <= 548;
        o_index_for_a3 <= 808;
        o_index_for_a4 <= 925;
        o_index_for_a5 <= 1071; 
    end
    1142: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 98;
        o_index_for_a1 <= 278;
        o_index_for_a2 <= 549;
        o_index_for_a3 <= 809;
        o_index_for_a4 <= 926;
        o_index_for_a5 <= 1072; 
    end
    1143: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 99;
        o_index_for_a1 <= 279;
        o_index_for_a2 <= 550;
        o_index_for_a3 <= 810;
        o_index_for_a4 <= 927;
        o_index_for_a5 <= 1073; 
    end
    1144: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 100;
        o_index_for_a1 <= 280;
        o_index_for_a2 <= 551;
        o_index_for_a3 <= 811;
        o_index_for_a4 <= 928;
        o_index_for_a5 <= 1074; 
    end
    1145: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 101;
        o_index_for_a1 <= 281;
        o_index_for_a2 <= 552;
        o_index_for_a3 <= 812;
        o_index_for_a4 <= 929;
        o_index_for_a5 <= 1075; 
    end
    1146: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 102;
        o_index_for_a1 <= 282;
        o_index_for_a2 <= 553;
        o_index_for_a3 <= 813;
        o_index_for_a4 <= 930;
        o_index_for_a5 <= 1076; 
    end
    1147: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 103;
        o_index_for_a1 <= 283;
        o_index_for_a2 <= 554;
        o_index_for_a3 <= 814;
        o_index_for_a4 <= 931;
        o_index_for_a5 <= 1077; 
    end
    1148: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 104;
        o_index_for_a1 <= 284;
        o_index_for_a2 <= 555;
        o_index_for_a3 <= 815;
        o_index_for_a4 <= 932;
        o_index_for_a5 <= 1078; 
    end
    1149: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 105;
        o_index_for_a1 <= 285;
        o_index_for_a2 <= 556;
        o_index_for_a3 <= 816;
        o_index_for_a4 <= 933;
        o_index_for_a5 <= 1079; 
    end
    1150: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 106;
        o_index_for_a1 <= 286;
        o_index_for_a2 <= 557;
        o_index_for_a3 <= 817;
        o_index_for_a4 <= 934;
        o_index_for_a5 <= 1080; 
    end
    1151: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 3; 
        o_index_for_a0 <= 107;
        o_index_for_a1 <= 287;
        o_index_for_a2 <= 558;
        o_index_for_a3 <= 818;
        o_index_for_a4 <= 935;
        o_index_for_a5 <= 1081; 
    end
    1152: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 7;
        o_index_for_a1 <= 480;
        o_index_for_a2 <= 1063;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1153: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 8;
        o_index_for_a1 <= 481;
        o_index_for_a2 <= 1064;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1154: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 9;
        o_index_for_a1 <= 482;
        o_index_for_a2 <= 1065;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1155: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 10;
        o_index_for_a1 <= 483;
        o_index_for_a2 <= 1066;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1156: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 11;
        o_index_for_a1 <= 484;
        o_index_for_a2 <= 1067;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1157: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 12;
        o_index_for_a1 <= 485;
        o_index_for_a2 <= 1068;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1158: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 13;
        o_index_for_a1 <= 486;
        o_index_for_a2 <= 1069;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1159: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 14;
        o_index_for_a1 <= 487;
        o_index_for_a2 <= 1070;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1160: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 15;
        o_index_for_a1 <= 488;
        o_index_for_a2 <= 1071;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1161: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 16;
        o_index_for_a1 <= 489;
        o_index_for_a2 <= 1072;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1162: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 17;
        o_index_for_a1 <= 490;
        o_index_for_a2 <= 1073;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1163: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 18;
        o_index_for_a1 <= 491;
        o_index_for_a2 <= 1074;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1164: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 19;
        o_index_for_a1 <= 492;
        o_index_for_a2 <= 1075;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1165: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 20;
        o_index_for_a1 <= 493;
        o_index_for_a2 <= 1076;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1166: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 21;
        o_index_for_a1 <= 494;
        o_index_for_a2 <= 1077;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1167: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 22;
        o_index_for_a1 <= 495;
        o_index_for_a2 <= 1078;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1168: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 23;
        o_index_for_a1 <= 496;
        o_index_for_a2 <= 1079;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1169: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 24;
        o_index_for_a1 <= 497;
        o_index_for_a2 <= 1080;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1170: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 25;
        o_index_for_a1 <= 498;
        o_index_for_a2 <= 1081;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1171: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 26;
        o_index_for_a1 <= 499;
        o_index_for_a2 <= 1082;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1172: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 27;
        o_index_for_a1 <= 500;
        o_index_for_a2 <= 1083;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1173: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 28;
        o_index_for_a1 <= 501;
        o_index_for_a2 <= 1084;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1174: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 29;
        o_index_for_a1 <= 502;
        o_index_for_a2 <= 1085;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1175: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 30;
        o_index_for_a1 <= 503;
        o_index_for_a2 <= 1086;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1176: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 31;
        o_index_for_a1 <= 504;
        o_index_for_a2 <= 1087;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1177: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 32;
        o_index_for_a1 <= 505;
        o_index_for_a2 <= 1088;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1178: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 33;
        o_index_for_a1 <= 506;
        o_index_for_a2 <= 1089;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1179: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 34;
        o_index_for_a1 <= 507;
        o_index_for_a2 <= 1090;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1180: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 35;
        o_index_for_a1 <= 508;
        o_index_for_a2 <= 1091;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1181: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 36;
        o_index_for_a1 <= 509;
        o_index_for_a2 <= 1092;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1182: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 37;
        o_index_for_a1 <= 510;
        o_index_for_a2 <= 1093;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1183: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 38;
        o_index_for_a1 <= 511;
        o_index_for_a2 <= 1094;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1184: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 39;
        o_index_for_a1 <= 512;
        o_index_for_a2 <= 1095;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1185: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 40;
        o_index_for_a1 <= 513;
        o_index_for_a2 <= 1096;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1186: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 41;
        o_index_for_a1 <= 514;
        o_index_for_a2 <= 1097;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1187: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 42;
        o_index_for_a1 <= 515;
        o_index_for_a2 <= 1098;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1188: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 43;
        o_index_for_a1 <= 516;
        o_index_for_a2 <= 1099;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1189: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 44;
        o_index_for_a1 <= 517;
        o_index_for_a2 <= 1100;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1190: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 45;
        o_index_for_a1 <= 518;
        o_index_for_a2 <= 1101;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1191: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 46;
        o_index_for_a1 <= 519;
        o_index_for_a2 <= 1102;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1192: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 47;
        o_index_for_a1 <= 520;
        o_index_for_a2 <= 1103;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1193: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 48;
        o_index_for_a1 <= 521;
        o_index_for_a2 <= 1104;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1194: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 49;
        o_index_for_a1 <= 522;
        o_index_for_a2 <= 1105;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1195: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 50;
        o_index_for_a1 <= 523;
        o_index_for_a2 <= 1106;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1196: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 51;
        o_index_for_a1 <= 524;
        o_index_for_a2 <= 1107;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1197: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 52;
        o_index_for_a1 <= 525;
        o_index_for_a2 <= 1108;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1198: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 53;
        o_index_for_a1 <= 526;
        o_index_for_a2 <= 1109;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1199: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 54;
        o_index_for_a1 <= 527;
        o_index_for_a2 <= 1110;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1200: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 55;
        o_index_for_a1 <= 528;
        o_index_for_a2 <= 1111;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1201: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 56;
        o_index_for_a1 <= 529;
        o_index_for_a2 <= 1112;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1202: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 57;
        o_index_for_a1 <= 530;
        o_index_for_a2 <= 1113;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1203: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 58;
        o_index_for_a1 <= 531;
        o_index_for_a2 <= 1114;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1204: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 59;
        o_index_for_a1 <= 532;
        o_index_for_a2 <= 1115;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1205: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 60;
        o_index_for_a1 <= 533;
        o_index_for_a2 <= 1116;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1206: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 61;
        o_index_for_a1 <= 534;
        o_index_for_a2 <= 1117;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1207: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 62;
        o_index_for_a1 <= 535;
        o_index_for_a2 <= 1118;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1208: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 63;
        o_index_for_a1 <= 536;
        o_index_for_a2 <= 1119;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1209: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 64;
        o_index_for_a1 <= 537;
        o_index_for_a2 <= 1120;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1210: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 65;
        o_index_for_a1 <= 538;
        o_index_for_a2 <= 1121;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1211: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 66;
        o_index_for_a1 <= 539;
        o_index_for_a2 <= 1122;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1212: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 67;
        o_index_for_a1 <= 540;
        o_index_for_a2 <= 1123;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1213: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 68;
        o_index_for_a1 <= 541;
        o_index_for_a2 <= 1124;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1214: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 69;
        o_index_for_a1 <= 542;
        o_index_for_a2 <= 1125;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1215: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 70;
        o_index_for_a1 <= 543;
        o_index_for_a2 <= 1126;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1216: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 71;
        o_index_for_a1 <= 544;
        o_index_for_a2 <= 1127;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1217: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 72;
        o_index_for_a1 <= 545;
        o_index_for_a2 <= 1128;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1218: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 73;
        o_index_for_a1 <= 546;
        o_index_for_a2 <= 1129;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1219: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 74;
        o_index_for_a1 <= 547;
        o_index_for_a2 <= 1130;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1220: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 75;
        o_index_for_a1 <= 548;
        o_index_for_a2 <= 1131;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1221: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 76;
        o_index_for_a1 <= 549;
        o_index_for_a2 <= 1132;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1222: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 77;
        o_index_for_a1 <= 550;
        o_index_for_a2 <= 1133;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1223: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 78;
        o_index_for_a1 <= 551;
        o_index_for_a2 <= 1134;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1224: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 79;
        o_index_for_a1 <= 552;
        o_index_for_a2 <= 1135;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1225: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 80;
        o_index_for_a1 <= 553;
        o_index_for_a2 <= 1136;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1226: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 81;
        o_index_for_a1 <= 554;
        o_index_for_a2 <= 1137;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1227: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 82;
        o_index_for_a1 <= 555;
        o_index_for_a2 <= 1138;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1228: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 83;
        o_index_for_a1 <= 556;
        o_index_for_a2 <= 1139;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1229: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 84;
        o_index_for_a1 <= 557;
        o_index_for_a2 <= 1140;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1230: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 85;
        o_index_for_a1 <= 558;
        o_index_for_a2 <= 1141;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1231: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 86;
        o_index_for_a1 <= 559;
        o_index_for_a2 <= 1142;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1232: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 87;
        o_index_for_a1 <= 560;
        o_index_for_a2 <= 1143;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1233: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 88;
        o_index_for_a1 <= 561;
        o_index_for_a2 <= 1144;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1234: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 89;
        o_index_for_a1 <= 562;
        o_index_for_a2 <= 1145;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1235: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 90;
        o_index_for_a1 <= 563;
        o_index_for_a2 <= 1146;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1236: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 91;
        o_index_for_a1 <= 564;
        o_index_for_a2 <= 1147;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1237: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 92;
        o_index_for_a1 <= 565;
        o_index_for_a2 <= 1148;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1238: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 93;
        o_index_for_a1 <= 566;
        o_index_for_a2 <= 1149;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1239: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 94;
        o_index_for_a1 <= 567;
        o_index_for_a2 <= 1150;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1240: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 95;
        o_index_for_a1 <= 568;
        o_index_for_a2 <= 1151;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1241: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 0;
        o_index_for_a1 <= 569;
        o_index_for_a2 <= 1056;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1242: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1;
        o_index_for_a1 <= 570;
        o_index_for_a2 <= 1057;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1243: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 2;
        o_index_for_a1 <= 571;
        o_index_for_a2 <= 1058;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1244: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 3;
        o_index_for_a1 <= 572;
        o_index_for_a2 <= 1059;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1245: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 4;
        o_index_for_a1 <= 573;
        o_index_for_a2 <= 1060;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1246: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 5;
        o_index_for_a1 <= 574;
        o_index_for_a2 <= 1061;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1247: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 4;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 6;
        o_index_for_a1 <= 575;
        o_index_for_a2 <= 1062;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1248: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 0;
        o_index_for_a1 <= 96;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1249: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1;
        o_index_for_a1 <= 97;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1250: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 2;
        o_index_for_a1 <= 98;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1251: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 3;
        o_index_for_a1 <= 99;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1252: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 4;
        o_index_for_a1 <= 100;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1253: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 5;
        o_index_for_a1 <= 101;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1254: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 6;
        o_index_for_a1 <= 102;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1255: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 7;
        o_index_for_a1 <= 103;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1256: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 8;
        o_index_for_a1 <= 104;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1257: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 9;
        o_index_for_a1 <= 105;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1258: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 10;
        o_index_for_a1 <= 106;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1259: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 11;
        o_index_for_a1 <= 107;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1260: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 12;
        o_index_for_a1 <= 108;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1261: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 13;
        o_index_for_a1 <= 109;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1262: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 14;
        o_index_for_a1 <= 110;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1263: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 15;
        o_index_for_a1 <= 111;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1264: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 16;
        o_index_for_a1 <= 112;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1265: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 17;
        o_index_for_a1 <= 113;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1266: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 18;
        o_index_for_a1 <= 114;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1267: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 19;
        o_index_for_a1 <= 115;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1268: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 20;
        o_index_for_a1 <= 116;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1269: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 21;
        o_index_for_a1 <= 117;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1270: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 22;
        o_index_for_a1 <= 118;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1271: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 23;
        o_index_for_a1 <= 119;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1272: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 24;
        o_index_for_a1 <= 120;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1273: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 25;
        o_index_for_a1 <= 121;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1274: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 26;
        o_index_for_a1 <= 122;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1275: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 27;
        o_index_for_a1 <= 123;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1276: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 28;
        o_index_for_a1 <= 124;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1277: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 29;
        o_index_for_a1 <= 125;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1278: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 30;
        o_index_for_a1 <= 126;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1279: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 31;
        o_index_for_a1 <= 127;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1280: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 32;
        o_index_for_a1 <= 128;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1281: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 33;
        o_index_for_a1 <= 129;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1282: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 34;
        o_index_for_a1 <= 130;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1283: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 35;
        o_index_for_a1 <= 131;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1284: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 36;
        o_index_for_a1 <= 132;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1285: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 37;
        o_index_for_a1 <= 133;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1286: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 38;
        o_index_for_a1 <= 134;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1287: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 39;
        o_index_for_a1 <= 135;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1288: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 40;
        o_index_for_a1 <= 136;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1289: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 41;
        o_index_for_a1 <= 137;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1290: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 42;
        o_index_for_a1 <= 138;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1291: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 43;
        o_index_for_a1 <= 139;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1292: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 44;
        o_index_for_a1 <= 140;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1293: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 45;
        o_index_for_a1 <= 141;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1294: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 46;
        o_index_for_a1 <= 142;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1295: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 47;
        o_index_for_a1 <= 143;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1296: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 48;
        o_index_for_a1 <= 144;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1297: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 49;
        o_index_for_a1 <= 145;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1298: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 50;
        o_index_for_a1 <= 146;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1299: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 51;
        o_index_for_a1 <= 147;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1300: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 52;
        o_index_for_a1 <= 148;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1301: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 53;
        o_index_for_a1 <= 149;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1302: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 54;
        o_index_for_a1 <= 150;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1303: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 55;
        o_index_for_a1 <= 151;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1304: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 56;
        o_index_for_a1 <= 152;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1305: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 57;
        o_index_for_a1 <= 153;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1306: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 58;
        o_index_for_a1 <= 154;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1307: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 59;
        o_index_for_a1 <= 155;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1308: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 60;
        o_index_for_a1 <= 156;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1309: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 61;
        o_index_for_a1 <= 157;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1310: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 62;
        o_index_for_a1 <= 158;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1311: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 63;
        o_index_for_a1 <= 159;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1312: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 64;
        o_index_for_a1 <= 160;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1313: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 65;
        o_index_for_a1 <= 161;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1314: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 66;
        o_index_for_a1 <= 162;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1315: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 67;
        o_index_for_a1 <= 163;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1316: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 68;
        o_index_for_a1 <= 164;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1317: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 69;
        o_index_for_a1 <= 165;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1318: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 70;
        o_index_for_a1 <= 166;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1319: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 71;
        o_index_for_a1 <= 167;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1320: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 72;
        o_index_for_a1 <= 168;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1321: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 73;
        o_index_for_a1 <= 169;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1322: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 74;
        o_index_for_a1 <= 170;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1323: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 75;
        o_index_for_a1 <= 171;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1324: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 76;
        o_index_for_a1 <= 172;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1325: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 77;
        o_index_for_a1 <= 173;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1326: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 78;
        o_index_for_a1 <= 174;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1327: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 79;
        o_index_for_a1 <= 175;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1328: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 80;
        o_index_for_a1 <= 176;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1329: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 81;
        o_index_for_a1 <= 177;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1330: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 82;
        o_index_for_a1 <= 178;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1331: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 83;
        o_index_for_a1 <= 179;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1332: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 84;
        o_index_for_a1 <= 180;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1333: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 85;
        o_index_for_a1 <= 181;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1334: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 86;
        o_index_for_a1 <= 182;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1335: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 87;
        o_index_for_a1 <= 183;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1336: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 88;
        o_index_for_a1 <= 184;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1337: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 89;
        o_index_for_a1 <= 185;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1338: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 90;
        o_index_for_a1 <= 186;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1339: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 91;
        o_index_for_a1 <= 187;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1340: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 92;
        o_index_for_a1 <= 188;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1341: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 93;
        o_index_for_a1 <= 189;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1342: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 94;
        o_index_for_a1 <= 190;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1343: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 95;
        o_index_for_a1 <= 191;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1344: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 96;
        o_index_for_a1 <= 192;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1345: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 97;
        o_index_for_a1 <= 193;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1346: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 98;
        o_index_for_a1 <= 194;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1347: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 99;
        o_index_for_a1 <= 195;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1348: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 100;
        o_index_for_a1 <= 196;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1349: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 101;
        o_index_for_a1 <= 197;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1350: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 102;
        o_index_for_a1 <= 198;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1351: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 103;
        o_index_for_a1 <= 199;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1352: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 104;
        o_index_for_a1 <= 200;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1353: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 105;
        o_index_for_a1 <= 201;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1354: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 106;
        o_index_for_a1 <= 202;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1355: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 107;
        o_index_for_a1 <= 203;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1356: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 108;
        o_index_for_a1 <= 204;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1357: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 109;
        o_index_for_a1 <= 205;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1358: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 110;
        o_index_for_a1 <= 206;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1359: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 111;
        o_index_for_a1 <= 207;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1360: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 112;
        o_index_for_a1 <= 208;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1361: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 113;
        o_index_for_a1 <= 209;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1362: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 114;
        o_index_for_a1 <= 210;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1363: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 115;
        o_index_for_a1 <= 211;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1364: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 116;
        o_index_for_a1 <= 212;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1365: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 117;
        o_index_for_a1 <= 213;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1366: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 118;
        o_index_for_a1 <= 214;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1367: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 119;
        o_index_for_a1 <= 215;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1368: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 120;
        o_index_for_a1 <= 216;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1369: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 121;
        o_index_for_a1 <= 217;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1370: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 122;
        o_index_for_a1 <= 218;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1371: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 123;
        o_index_for_a1 <= 219;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1372: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 124;
        o_index_for_a1 <= 220;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1373: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 125;
        o_index_for_a1 <= 221;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1374: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 126;
        o_index_for_a1 <= 222;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1375: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 127;
        o_index_for_a1 <= 223;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1376: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 128;
        o_index_for_a1 <= 224;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1377: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 129;
        o_index_for_a1 <= 225;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1378: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 130;
        o_index_for_a1 <= 226;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1379: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 131;
        o_index_for_a1 <= 227;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1380: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 132;
        o_index_for_a1 <= 228;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1381: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 133;
        o_index_for_a1 <= 229;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1382: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 134;
        o_index_for_a1 <= 230;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1383: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 135;
        o_index_for_a1 <= 231;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1384: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 136;
        o_index_for_a1 <= 232;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1385: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 137;
        o_index_for_a1 <= 233;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1386: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 138;
        o_index_for_a1 <= 234;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1387: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 139;
        o_index_for_a1 <= 235;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1388: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 140;
        o_index_for_a1 <= 236;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1389: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 141;
        o_index_for_a1 <= 237;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1390: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 142;
        o_index_for_a1 <= 238;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1391: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 143;
        o_index_for_a1 <= 239;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1392: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 144;
        o_index_for_a1 <= 240;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1393: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 145;
        o_index_for_a1 <= 241;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1394: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 146;
        o_index_for_a1 <= 242;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1395: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 147;
        o_index_for_a1 <= 243;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1396: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 148;
        o_index_for_a1 <= 244;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1397: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 149;
        o_index_for_a1 <= 245;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1398: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 150;
        o_index_for_a1 <= 246;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1399: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 151;
        o_index_for_a1 <= 247;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1400: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 152;
        o_index_for_a1 <= 248;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1401: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 153;
        o_index_for_a1 <= 249;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1402: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 154;
        o_index_for_a1 <= 250;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1403: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 155;
        o_index_for_a1 <= 251;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1404: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 156;
        o_index_for_a1 <= 252;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1405: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 157;
        o_index_for_a1 <= 253;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1406: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 158;
        o_index_for_a1 <= 254;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1407: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 159;
        o_index_for_a1 <= 255;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1408: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 160;
        o_index_for_a1 <= 256;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1409: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 161;
        o_index_for_a1 <= 257;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1410: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 162;
        o_index_for_a1 <= 258;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1411: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 163;
        o_index_for_a1 <= 259;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1412: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 164;
        o_index_for_a1 <= 260;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1413: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 165;
        o_index_for_a1 <= 261;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1414: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 166;
        o_index_for_a1 <= 262;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1415: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 167;
        o_index_for_a1 <= 263;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1416: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 168;
        o_index_for_a1 <= 264;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1417: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 169;
        o_index_for_a1 <= 265;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1418: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 170;
        o_index_for_a1 <= 266;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1419: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 171;
        o_index_for_a1 <= 267;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1420: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 172;
        o_index_for_a1 <= 268;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1421: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 173;
        o_index_for_a1 <= 269;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1422: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 174;
        o_index_for_a1 <= 270;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1423: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 175;
        o_index_for_a1 <= 271;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1424: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 176;
        o_index_for_a1 <= 272;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1425: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 177;
        o_index_for_a1 <= 273;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1426: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 178;
        o_index_for_a1 <= 274;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1427: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 179;
        o_index_for_a1 <= 275;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1428: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 180;
        o_index_for_a1 <= 276;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1429: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 181;
        o_index_for_a1 <= 277;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1430: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 182;
        o_index_for_a1 <= 278;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1431: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 183;
        o_index_for_a1 <= 279;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1432: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 184;
        o_index_for_a1 <= 280;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1433: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 185;
        o_index_for_a1 <= 281;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1434: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 186;
        o_index_for_a1 <= 282;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1435: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 187;
        o_index_for_a1 <= 283;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1436: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 188;
        o_index_for_a1 <= 284;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1437: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 189;
        o_index_for_a1 <= 285;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1438: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 190;
        o_index_for_a1 <= 286;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1439: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 191;
        o_index_for_a1 <= 287;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1440: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 192;
        o_index_for_a1 <= 288;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1441: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 193;
        o_index_for_a1 <= 289;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1442: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 194;
        o_index_for_a1 <= 290;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1443: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 195;
        o_index_for_a1 <= 291;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1444: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 196;
        o_index_for_a1 <= 292;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1445: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 197;
        o_index_for_a1 <= 293;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1446: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 198;
        o_index_for_a1 <= 294;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1447: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 199;
        o_index_for_a1 <= 295;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1448: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 200;
        o_index_for_a1 <= 296;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1449: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 201;
        o_index_for_a1 <= 297;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1450: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 202;
        o_index_for_a1 <= 298;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1451: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 203;
        o_index_for_a1 <= 299;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1452: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 204;
        o_index_for_a1 <= 300;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1453: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 205;
        o_index_for_a1 <= 301;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1454: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 206;
        o_index_for_a1 <= 302;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1455: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 207;
        o_index_for_a1 <= 303;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1456: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 208;
        o_index_for_a1 <= 304;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1457: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 209;
        o_index_for_a1 <= 305;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1458: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 210;
        o_index_for_a1 <= 306;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1459: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 211;
        o_index_for_a1 <= 307;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1460: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 212;
        o_index_for_a1 <= 308;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1461: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 213;
        o_index_for_a1 <= 309;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1462: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 214;
        o_index_for_a1 <= 310;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1463: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 215;
        o_index_for_a1 <= 311;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1464: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 216;
        o_index_for_a1 <= 312;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1465: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 217;
        o_index_for_a1 <= 313;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1466: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 218;
        o_index_for_a1 <= 314;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1467: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 219;
        o_index_for_a1 <= 315;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1468: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 220;
        o_index_for_a1 <= 316;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1469: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 221;
        o_index_for_a1 <= 317;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1470: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 222;
        o_index_for_a1 <= 318;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1471: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 223;
        o_index_for_a1 <= 319;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1472: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 224;
        o_index_for_a1 <= 320;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1473: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 225;
        o_index_for_a1 <= 321;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1474: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 226;
        o_index_for_a1 <= 322;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1475: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 227;
        o_index_for_a1 <= 323;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1476: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 228;
        o_index_for_a1 <= 324;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1477: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 229;
        o_index_for_a1 <= 325;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1478: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 230;
        o_index_for_a1 <= 326;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1479: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 231;
        o_index_for_a1 <= 327;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1480: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 232;
        o_index_for_a1 <= 328;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1481: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 233;
        o_index_for_a1 <= 329;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1482: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 234;
        o_index_for_a1 <= 330;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1483: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 235;
        o_index_for_a1 <= 331;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1484: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 236;
        o_index_for_a1 <= 332;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1485: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 237;
        o_index_for_a1 <= 333;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1486: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 238;
        o_index_for_a1 <= 334;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1487: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 239;
        o_index_for_a1 <= 335;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1488: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 240;
        o_index_for_a1 <= 336;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1489: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 241;
        o_index_for_a1 <= 337;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1490: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 242;
        o_index_for_a1 <= 338;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1491: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 243;
        o_index_for_a1 <= 339;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1492: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 244;
        o_index_for_a1 <= 340;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1493: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 245;
        o_index_for_a1 <= 341;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1494: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 246;
        o_index_for_a1 <= 342;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1495: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 247;
        o_index_for_a1 <= 343;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1496: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 248;
        o_index_for_a1 <= 344;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1497: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 249;
        o_index_for_a1 <= 345;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1498: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 250;
        o_index_for_a1 <= 346;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1499: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 251;
        o_index_for_a1 <= 347;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1500: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 252;
        o_index_for_a1 <= 348;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1501: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 253;
        o_index_for_a1 <= 349;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1502: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 254;
        o_index_for_a1 <= 350;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1503: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 255;
        o_index_for_a1 <= 351;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1504: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 256;
        o_index_for_a1 <= 352;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1505: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 257;
        o_index_for_a1 <= 353;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1506: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 258;
        o_index_for_a1 <= 354;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1507: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 259;
        o_index_for_a1 <= 355;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1508: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 260;
        o_index_for_a1 <= 356;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1509: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 261;
        o_index_for_a1 <= 357;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1510: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 262;
        o_index_for_a1 <= 358;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1511: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 263;
        o_index_for_a1 <= 359;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1512: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 264;
        o_index_for_a1 <= 360;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1513: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 265;
        o_index_for_a1 <= 361;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1514: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 266;
        o_index_for_a1 <= 362;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1515: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 267;
        o_index_for_a1 <= 363;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1516: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 268;
        o_index_for_a1 <= 364;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1517: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 269;
        o_index_for_a1 <= 365;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1518: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 270;
        o_index_for_a1 <= 366;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1519: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 271;
        o_index_for_a1 <= 367;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1520: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 272;
        o_index_for_a1 <= 368;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1521: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 273;
        o_index_for_a1 <= 369;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1522: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 274;
        o_index_for_a1 <= 370;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1523: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 275;
        o_index_for_a1 <= 371;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1524: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 276;
        o_index_for_a1 <= 372;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1525: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 277;
        o_index_for_a1 <= 373;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1526: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 278;
        o_index_for_a1 <= 374;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1527: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 279;
        o_index_for_a1 <= 375;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1528: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 280;
        o_index_for_a1 <= 376;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1529: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 281;
        o_index_for_a1 <= 377;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1530: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 282;
        o_index_for_a1 <= 378;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1531: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 283;
        o_index_for_a1 <= 379;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1532: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 284;
        o_index_for_a1 <= 380;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1533: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 285;
        o_index_for_a1 <= 381;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1534: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 286;
        o_index_for_a1 <= 382;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1535: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 287;
        o_index_for_a1 <= 383;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1536: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 288;
        o_index_for_a1 <= 384;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1537: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 289;
        o_index_for_a1 <= 385;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1538: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 290;
        o_index_for_a1 <= 386;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1539: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 291;
        o_index_for_a1 <= 387;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1540: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 292;
        o_index_for_a1 <= 388;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1541: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 293;
        o_index_for_a1 <= 389;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1542: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 294;
        o_index_for_a1 <= 390;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1543: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 295;
        o_index_for_a1 <= 391;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1544: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 296;
        o_index_for_a1 <= 392;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1545: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 297;
        o_index_for_a1 <= 393;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1546: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 298;
        o_index_for_a1 <= 394;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1547: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 299;
        o_index_for_a1 <= 395;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1548: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 300;
        o_index_for_a1 <= 396;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1549: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 301;
        o_index_for_a1 <= 397;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1550: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 302;
        o_index_for_a1 <= 398;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1551: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 303;
        o_index_for_a1 <= 399;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1552: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 304;
        o_index_for_a1 <= 400;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1553: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 305;
        o_index_for_a1 <= 401;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1554: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 306;
        o_index_for_a1 <= 402;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1555: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 307;
        o_index_for_a1 <= 403;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1556: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 308;
        o_index_for_a1 <= 404;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1557: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 309;
        o_index_for_a1 <= 405;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1558: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 310;
        o_index_for_a1 <= 406;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1559: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 311;
        o_index_for_a1 <= 407;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1560: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 312;
        o_index_for_a1 <= 408;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1561: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 313;
        o_index_for_a1 <= 409;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1562: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 314;
        o_index_for_a1 <= 410;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1563: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 315;
        o_index_for_a1 <= 411;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1564: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 316;
        o_index_for_a1 <= 412;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1565: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 317;
        o_index_for_a1 <= 413;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1566: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 318;
        o_index_for_a1 <= 414;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1567: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 319;
        o_index_for_a1 <= 415;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1568: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 320;
        o_index_for_a1 <= 416;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1569: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 321;
        o_index_for_a1 <= 417;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1570: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 322;
        o_index_for_a1 <= 418;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1571: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 323;
        o_index_for_a1 <= 419;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1572: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 324;
        o_index_for_a1 <= 420;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1573: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 325;
        o_index_for_a1 <= 421;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1574: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 326;
        o_index_for_a1 <= 422;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1575: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 327;
        o_index_for_a1 <= 423;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1576: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 328;
        o_index_for_a1 <= 424;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1577: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 329;
        o_index_for_a1 <= 425;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1578: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 330;
        o_index_for_a1 <= 426;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1579: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 331;
        o_index_for_a1 <= 427;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1580: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 332;
        o_index_for_a1 <= 428;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1581: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 333;
        o_index_for_a1 <= 429;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1582: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 334;
        o_index_for_a1 <= 430;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1583: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 335;
        o_index_for_a1 <= 431;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1584: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 336;
        o_index_for_a1 <= 432;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1585: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 337;
        o_index_for_a1 <= 433;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1586: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 338;
        o_index_for_a1 <= 434;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1587: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 339;
        o_index_for_a1 <= 435;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1588: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 340;
        o_index_for_a1 <= 436;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1589: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 341;
        o_index_for_a1 <= 437;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1590: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 342;
        o_index_for_a1 <= 438;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1591: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 343;
        o_index_for_a1 <= 439;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1592: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 344;
        o_index_for_a1 <= 440;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1593: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 345;
        o_index_for_a1 <= 441;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1594: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 346;
        o_index_for_a1 <= 442;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1595: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 347;
        o_index_for_a1 <= 443;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1596: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 348;
        o_index_for_a1 <= 444;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1597: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 349;
        o_index_for_a1 <= 445;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1598: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 350;
        o_index_for_a1 <= 446;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1599: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 351;
        o_index_for_a1 <= 447;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1600: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 352;
        o_index_for_a1 <= 448;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1601: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 353;
        o_index_for_a1 <= 449;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1602: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 354;
        o_index_for_a1 <= 450;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1603: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 355;
        o_index_for_a1 <= 451;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1604: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 356;
        o_index_for_a1 <= 452;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1605: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 357;
        o_index_for_a1 <= 453;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1606: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 358;
        o_index_for_a1 <= 454;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1607: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 359;
        o_index_for_a1 <= 455;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1608: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 360;
        o_index_for_a1 <= 456;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1609: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 361;
        o_index_for_a1 <= 457;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1610: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 362;
        o_index_for_a1 <= 458;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1611: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 363;
        o_index_for_a1 <= 459;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1612: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 364;
        o_index_for_a1 <= 460;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1613: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 365;
        o_index_for_a1 <= 461;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1614: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 366;
        o_index_for_a1 <= 462;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1615: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 367;
        o_index_for_a1 <= 463;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1616: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 368;
        o_index_for_a1 <= 464;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1617: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 369;
        o_index_for_a1 <= 465;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1618: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 370;
        o_index_for_a1 <= 466;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1619: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 371;
        o_index_for_a1 <= 467;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1620: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 372;
        o_index_for_a1 <= 468;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1621: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 373;
        o_index_for_a1 <= 469;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1622: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 374;
        o_index_for_a1 <= 470;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1623: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 375;
        o_index_for_a1 <= 471;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1624: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 376;
        o_index_for_a1 <= 472;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1625: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 377;
        o_index_for_a1 <= 473;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1626: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 378;
        o_index_for_a1 <= 474;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1627: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 379;
        o_index_for_a1 <= 475;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1628: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 380;
        o_index_for_a1 <= 476;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1629: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 381;
        o_index_for_a1 <= 477;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1630: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 382;
        o_index_for_a1 <= 478;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1631: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 383;
        o_index_for_a1 <= 479;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1632: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 384;
        o_index_for_a1 <= 480;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1633: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 385;
        o_index_for_a1 <= 481;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1634: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 386;
        o_index_for_a1 <= 482;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1635: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 387;
        o_index_for_a1 <= 483;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1636: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 388;
        o_index_for_a1 <= 484;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1637: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 389;
        o_index_for_a1 <= 485;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1638: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 390;
        o_index_for_a1 <= 486;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1639: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 391;
        o_index_for_a1 <= 487;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1640: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 392;
        o_index_for_a1 <= 488;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1641: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 393;
        o_index_for_a1 <= 489;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1642: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 394;
        o_index_for_a1 <= 490;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1643: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 395;
        o_index_for_a1 <= 491;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1644: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 396;
        o_index_for_a1 <= 492;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1645: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 397;
        o_index_for_a1 <= 493;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1646: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 398;
        o_index_for_a1 <= 494;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1647: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 399;
        o_index_for_a1 <= 495;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1648: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 400;
        o_index_for_a1 <= 496;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1649: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 401;
        o_index_for_a1 <= 497;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1650: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 402;
        o_index_for_a1 <= 498;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1651: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 403;
        o_index_for_a1 <= 499;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1652: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 404;
        o_index_for_a1 <= 500;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1653: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 405;
        o_index_for_a1 <= 501;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1654: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 406;
        o_index_for_a1 <= 502;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1655: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 407;
        o_index_for_a1 <= 503;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1656: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 408;
        o_index_for_a1 <= 504;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1657: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 409;
        o_index_for_a1 <= 505;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1658: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 410;
        o_index_for_a1 <= 506;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1659: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 411;
        o_index_for_a1 <= 507;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1660: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 412;
        o_index_for_a1 <= 508;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1661: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 413;
        o_index_for_a1 <= 509;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1662: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 414;
        o_index_for_a1 <= 510;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1663: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 415;
        o_index_for_a1 <= 511;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1664: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 416;
        o_index_for_a1 <= 512;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1665: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 417;
        o_index_for_a1 <= 513;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1666: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 418;
        o_index_for_a1 <= 514;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1667: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 419;
        o_index_for_a1 <= 515;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1668: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 420;
        o_index_for_a1 <= 516;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1669: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 421;
        o_index_for_a1 <= 517;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1670: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 422;
        o_index_for_a1 <= 518;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1671: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 423;
        o_index_for_a1 <= 519;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1672: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 424;
        o_index_for_a1 <= 520;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1673: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 425;
        o_index_for_a1 <= 521;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1674: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 426;
        o_index_for_a1 <= 522;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1675: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 427;
        o_index_for_a1 <= 523;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1676: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 428;
        o_index_for_a1 <= 524;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1677: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 429;
        o_index_for_a1 <= 525;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1678: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 430;
        o_index_for_a1 <= 526;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1679: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 431;
        o_index_for_a1 <= 527;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1680: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 432;
        o_index_for_a1 <= 528;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1681: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 433;
        o_index_for_a1 <= 529;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1682: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 434;
        o_index_for_a1 <= 530;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1683: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 435;
        o_index_for_a1 <= 531;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1684: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 436;
        o_index_for_a1 <= 532;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1685: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 437;
        o_index_for_a1 <= 533;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1686: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 438;
        o_index_for_a1 <= 534;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1687: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 439;
        o_index_for_a1 <= 535;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1688: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 440;
        o_index_for_a1 <= 536;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1689: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 441;
        o_index_for_a1 <= 537;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1690: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 442;
        o_index_for_a1 <= 538;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1691: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 443;
        o_index_for_a1 <= 539;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1692: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 444;
        o_index_for_a1 <= 540;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1693: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 445;
        o_index_for_a1 <= 541;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1694: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 446;
        o_index_for_a1 <= 542;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1695: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 447;
        o_index_for_a1 <= 543;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1696: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 448;
        o_index_for_a1 <= 544;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1697: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 449;
        o_index_for_a1 <= 545;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1698: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 450;
        o_index_for_a1 <= 546;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1699: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 451;
        o_index_for_a1 <= 547;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1700: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 452;
        o_index_for_a1 <= 548;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1701: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 453;
        o_index_for_a1 <= 549;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1702: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 454;
        o_index_for_a1 <= 550;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1703: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 455;
        o_index_for_a1 <= 551;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1704: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 456;
        o_index_for_a1 <= 552;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1705: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 457;
        o_index_for_a1 <= 553;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1706: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 458;
        o_index_for_a1 <= 554;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1707: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 459;
        o_index_for_a1 <= 555;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1708: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 460;
        o_index_for_a1 <= 556;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1709: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 461;
        o_index_for_a1 <= 557;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1710: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 462;
        o_index_for_a1 <= 558;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1711: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 463;
        o_index_for_a1 <= 559;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1712: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 464;
        o_index_for_a1 <= 560;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1713: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 465;
        o_index_for_a1 <= 561;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1714: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 466;
        o_index_for_a1 <= 562;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1715: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 467;
        o_index_for_a1 <= 563;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1716: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 468;
        o_index_for_a1 <= 564;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1717: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 469;
        o_index_for_a1 <= 565;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1718: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 470;
        o_index_for_a1 <= 566;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1719: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 471;
        o_index_for_a1 <= 567;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1720: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 472;
        o_index_for_a1 <= 568;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1721: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 473;
        o_index_for_a1 <= 569;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1722: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 474;
        o_index_for_a1 <= 570;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1723: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 475;
        o_index_for_a1 <= 571;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1724: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 476;
        o_index_for_a1 <= 572;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1725: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 477;
        o_index_for_a1 <= 573;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1726: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 478;
        o_index_for_a1 <= 574;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1727: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 479;
        o_index_for_a1 <= 575;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1728: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 480;
        o_index_for_a1 <= 576;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1729: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 481;
        o_index_for_a1 <= 577;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1730: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 482;
        o_index_for_a1 <= 578;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1731: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 483;
        o_index_for_a1 <= 579;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1732: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 484;
        o_index_for_a1 <= 580;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1733: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 485;
        o_index_for_a1 <= 581;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1734: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 486;
        o_index_for_a1 <= 582;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1735: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 487;
        o_index_for_a1 <= 583;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1736: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 488;
        o_index_for_a1 <= 584;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1737: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 489;
        o_index_for_a1 <= 585;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1738: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 490;
        o_index_for_a1 <= 586;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1739: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 491;
        o_index_for_a1 <= 587;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1740: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 492;
        o_index_for_a1 <= 588;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1741: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 493;
        o_index_for_a1 <= 589;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1742: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 494;
        o_index_for_a1 <= 590;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1743: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 495;
        o_index_for_a1 <= 591;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1744: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 496;
        o_index_for_a1 <= 592;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1745: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 497;
        o_index_for_a1 <= 593;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1746: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 498;
        o_index_for_a1 <= 594;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1747: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 499;
        o_index_for_a1 <= 595;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1748: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 500;
        o_index_for_a1 <= 596;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1749: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 501;
        o_index_for_a1 <= 597;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1750: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 502;
        o_index_for_a1 <= 598;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1751: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 503;
        o_index_for_a1 <= 599;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1752: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 504;
        o_index_for_a1 <= 600;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1753: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 505;
        o_index_for_a1 <= 601;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1754: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 506;
        o_index_for_a1 <= 602;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1755: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 507;
        o_index_for_a1 <= 603;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1756: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 508;
        o_index_for_a1 <= 604;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1757: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 509;
        o_index_for_a1 <= 605;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1758: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 510;
        o_index_for_a1 <= 606;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1759: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 511;
        o_index_for_a1 <= 607;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1760: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 512;
        o_index_for_a1 <= 608;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1761: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 513;
        o_index_for_a1 <= 609;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1762: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 514;
        o_index_for_a1 <= 610;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1763: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 515;
        o_index_for_a1 <= 611;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1764: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 516;
        o_index_for_a1 <= 612;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1765: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 517;
        o_index_for_a1 <= 613;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1766: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 518;
        o_index_for_a1 <= 614;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1767: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 519;
        o_index_for_a1 <= 615;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1768: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 520;
        o_index_for_a1 <= 616;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1769: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 521;
        o_index_for_a1 <= 617;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1770: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 522;
        o_index_for_a1 <= 618;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1771: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 523;
        o_index_for_a1 <= 619;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1772: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 524;
        o_index_for_a1 <= 620;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1773: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 525;
        o_index_for_a1 <= 621;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1774: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 526;
        o_index_for_a1 <= 622;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1775: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 527;
        o_index_for_a1 <= 623;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1776: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 528;
        o_index_for_a1 <= 624;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1777: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 529;
        o_index_for_a1 <= 625;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1778: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 530;
        o_index_for_a1 <= 626;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1779: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 531;
        o_index_for_a1 <= 627;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1780: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 532;
        o_index_for_a1 <= 628;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1781: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 533;
        o_index_for_a1 <= 629;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1782: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 534;
        o_index_for_a1 <= 630;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1783: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 535;
        o_index_for_a1 <= 631;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1784: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 536;
        o_index_for_a1 <= 632;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1785: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 537;
        o_index_for_a1 <= 633;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1786: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 538;
        o_index_for_a1 <= 634;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1787: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 539;
        o_index_for_a1 <= 635;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1788: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 540;
        o_index_for_a1 <= 636;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1789: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 541;
        o_index_for_a1 <= 637;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1790: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 542;
        o_index_for_a1 <= 638;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1791: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 543;
        o_index_for_a1 <= 639;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1792: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 544;
        o_index_for_a1 <= 640;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1793: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 545;
        o_index_for_a1 <= 641;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1794: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 546;
        o_index_for_a1 <= 642;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1795: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 547;
        o_index_for_a1 <= 643;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1796: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 548;
        o_index_for_a1 <= 644;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1797: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 549;
        o_index_for_a1 <= 645;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1798: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 550;
        o_index_for_a1 <= 646;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1799: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 551;
        o_index_for_a1 <= 647;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1800: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 552;
        o_index_for_a1 <= 648;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1801: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 553;
        o_index_for_a1 <= 649;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1802: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 554;
        o_index_for_a1 <= 650;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1803: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 555;
        o_index_for_a1 <= 651;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1804: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 556;
        o_index_for_a1 <= 652;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1805: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 557;
        o_index_for_a1 <= 653;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1806: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 558;
        o_index_for_a1 <= 654;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1807: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 559;
        o_index_for_a1 <= 655;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1808: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 560;
        o_index_for_a1 <= 656;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1809: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 561;
        o_index_for_a1 <= 657;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1810: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 562;
        o_index_for_a1 <= 658;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1811: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 563;
        o_index_for_a1 <= 659;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1812: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 564;
        o_index_for_a1 <= 660;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1813: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 565;
        o_index_for_a1 <= 661;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1814: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 566;
        o_index_for_a1 <= 662;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1815: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 567;
        o_index_for_a1 <= 663;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1816: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 568;
        o_index_for_a1 <= 664;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1817: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 569;
        o_index_for_a1 <= 665;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1818: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 570;
        o_index_for_a1 <= 666;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1819: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 571;
        o_index_for_a1 <= 667;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1820: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 572;
        o_index_for_a1 <= 668;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1821: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 573;
        o_index_for_a1 <= 669;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1822: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 574;
        o_index_for_a1 <= 670;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1823: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 575;
        o_index_for_a1 <= 671;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1824: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 576;
        o_index_for_a1 <= 672;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1825: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 577;
        o_index_for_a1 <= 673;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1826: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 578;
        o_index_for_a1 <= 674;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1827: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 579;
        o_index_for_a1 <= 675;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1828: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 580;
        o_index_for_a1 <= 676;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1829: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 581;
        o_index_for_a1 <= 677;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1830: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 582;
        o_index_for_a1 <= 678;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1831: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 583;
        o_index_for_a1 <= 679;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1832: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 584;
        o_index_for_a1 <= 680;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1833: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 585;
        o_index_for_a1 <= 681;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1834: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 586;
        o_index_for_a1 <= 682;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1835: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 587;
        o_index_for_a1 <= 683;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1836: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 588;
        o_index_for_a1 <= 684;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1837: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 589;
        o_index_for_a1 <= 685;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1838: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 590;
        o_index_for_a1 <= 686;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1839: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 591;
        o_index_for_a1 <= 687;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1840: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 592;
        o_index_for_a1 <= 688;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1841: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 593;
        o_index_for_a1 <= 689;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1842: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 594;
        o_index_for_a1 <= 690;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1843: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 595;
        o_index_for_a1 <= 691;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1844: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 596;
        o_index_for_a1 <= 692;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1845: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 597;
        o_index_for_a1 <= 693;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1846: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 598;
        o_index_for_a1 <= 694;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1847: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 599;
        o_index_for_a1 <= 695;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1848: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 600;
        o_index_for_a1 <= 696;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1849: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 601;
        o_index_for_a1 <= 697;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1850: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 602;
        o_index_for_a1 <= 698;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1851: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 603;
        o_index_for_a1 <= 699;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1852: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 604;
        o_index_for_a1 <= 700;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1853: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 605;
        o_index_for_a1 <= 701;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1854: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 606;
        o_index_for_a1 <= 702;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1855: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 607;
        o_index_for_a1 <= 703;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1856: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 608;
        o_index_for_a1 <= 704;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1857: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 609;
        o_index_for_a1 <= 705;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1858: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 610;
        o_index_for_a1 <= 706;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1859: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 611;
        o_index_for_a1 <= 707;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1860: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 612;
        o_index_for_a1 <= 708;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1861: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 613;
        o_index_for_a1 <= 709;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1862: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 614;
        o_index_for_a1 <= 710;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1863: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 615;
        o_index_for_a1 <= 711;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1864: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 616;
        o_index_for_a1 <= 712;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1865: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 617;
        o_index_for_a1 <= 713;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1866: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 618;
        o_index_for_a1 <= 714;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1867: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 619;
        o_index_for_a1 <= 715;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1868: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 620;
        o_index_for_a1 <= 716;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1869: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 621;
        o_index_for_a1 <= 717;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1870: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 622;
        o_index_for_a1 <= 718;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1871: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 623;
        o_index_for_a1 <= 719;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1872: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 624;
        o_index_for_a1 <= 720;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1873: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 625;
        o_index_for_a1 <= 721;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1874: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 626;
        o_index_for_a1 <= 722;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1875: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 627;
        o_index_for_a1 <= 723;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1876: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 628;
        o_index_for_a1 <= 724;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1877: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 629;
        o_index_for_a1 <= 725;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1878: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 630;
        o_index_for_a1 <= 726;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1879: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 631;
        o_index_for_a1 <= 727;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1880: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 632;
        o_index_for_a1 <= 728;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1881: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 633;
        o_index_for_a1 <= 729;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1882: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 634;
        o_index_for_a1 <= 730;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1883: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 635;
        o_index_for_a1 <= 731;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1884: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 636;
        o_index_for_a1 <= 732;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1885: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 637;
        o_index_for_a1 <= 733;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1886: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 638;
        o_index_for_a1 <= 734;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1887: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 639;
        o_index_for_a1 <= 735;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1888: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 640;
        o_index_for_a1 <= 736;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1889: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 641;
        o_index_for_a1 <= 737;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1890: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 642;
        o_index_for_a1 <= 738;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1891: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 643;
        o_index_for_a1 <= 739;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1892: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 644;
        o_index_for_a1 <= 740;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1893: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 645;
        o_index_for_a1 <= 741;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1894: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 646;
        o_index_for_a1 <= 742;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1895: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 647;
        o_index_for_a1 <= 743;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1896: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 648;
        o_index_for_a1 <= 744;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1897: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 649;
        o_index_for_a1 <= 745;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1898: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 650;
        o_index_for_a1 <= 746;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1899: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 651;
        o_index_for_a1 <= 747;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1900: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 652;
        o_index_for_a1 <= 748;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1901: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 653;
        o_index_for_a1 <= 749;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1902: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 654;
        o_index_for_a1 <= 750;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1903: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 655;
        o_index_for_a1 <= 751;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1904: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 656;
        o_index_for_a1 <= 752;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1905: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 657;
        o_index_for_a1 <= 753;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1906: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 658;
        o_index_for_a1 <= 754;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1907: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 659;
        o_index_for_a1 <= 755;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1908: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 660;
        o_index_for_a1 <= 756;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1909: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 661;
        o_index_for_a1 <= 757;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1910: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 662;
        o_index_for_a1 <= 758;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1911: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 663;
        o_index_for_a1 <= 759;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1912: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 664;
        o_index_for_a1 <= 760;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1913: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 665;
        o_index_for_a1 <= 761;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1914: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 666;
        o_index_for_a1 <= 762;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1915: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 667;
        o_index_for_a1 <= 763;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1916: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 668;
        o_index_for_a1 <= 764;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1917: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 669;
        o_index_for_a1 <= 765;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1918: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 670;
        o_index_for_a1 <= 766;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1919: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 671;
        o_index_for_a1 <= 767;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1920: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 672;
        o_index_for_a1 <= 768;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1921: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 673;
        o_index_for_a1 <= 769;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1922: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 674;
        o_index_for_a1 <= 770;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1923: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 675;
        o_index_for_a1 <= 771;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1924: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 676;
        o_index_for_a1 <= 772;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1925: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 677;
        o_index_for_a1 <= 773;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1926: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 678;
        o_index_for_a1 <= 774;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1927: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 679;
        o_index_for_a1 <= 775;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1928: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 680;
        o_index_for_a1 <= 776;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1929: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 681;
        o_index_for_a1 <= 777;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1930: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 682;
        o_index_for_a1 <= 778;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1931: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 683;
        o_index_for_a1 <= 779;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1932: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 684;
        o_index_for_a1 <= 780;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1933: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 685;
        o_index_for_a1 <= 781;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1934: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 686;
        o_index_for_a1 <= 782;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1935: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 687;
        o_index_for_a1 <= 783;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1936: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 688;
        o_index_for_a1 <= 784;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1937: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 689;
        o_index_for_a1 <= 785;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1938: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 690;
        o_index_for_a1 <= 786;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1939: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 691;
        o_index_for_a1 <= 787;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1940: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 692;
        o_index_for_a1 <= 788;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1941: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 693;
        o_index_for_a1 <= 789;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1942: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 694;
        o_index_for_a1 <= 790;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1943: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 695;
        o_index_for_a1 <= 791;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1944: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 696;
        o_index_for_a1 <= 792;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1945: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 697;
        o_index_for_a1 <= 793;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1946: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 698;
        o_index_for_a1 <= 794;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1947: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 699;
        o_index_for_a1 <= 795;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1948: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 700;
        o_index_for_a1 <= 796;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1949: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 701;
        o_index_for_a1 <= 797;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1950: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 702;
        o_index_for_a1 <= 798;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1951: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 703;
        o_index_for_a1 <= 799;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1952: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 704;
        o_index_for_a1 <= 800;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1953: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 705;
        o_index_for_a1 <= 801;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1954: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 706;
        o_index_for_a1 <= 802;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1955: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 707;
        o_index_for_a1 <= 803;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1956: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 708;
        o_index_for_a1 <= 804;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1957: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 709;
        o_index_for_a1 <= 805;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1958: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 710;
        o_index_for_a1 <= 806;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1959: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 711;
        o_index_for_a1 <= 807;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1960: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 712;
        o_index_for_a1 <= 808;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1961: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 713;
        o_index_for_a1 <= 809;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1962: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 714;
        o_index_for_a1 <= 810;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1963: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 715;
        o_index_for_a1 <= 811;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1964: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 716;
        o_index_for_a1 <= 812;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1965: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 717;
        o_index_for_a1 <= 813;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1966: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 718;
        o_index_for_a1 <= 814;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1967: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 719;
        o_index_for_a1 <= 815;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1968: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 720;
        o_index_for_a1 <= 816;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1969: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 721;
        o_index_for_a1 <= 817;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1970: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 722;
        o_index_for_a1 <= 818;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1971: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 723;
        o_index_for_a1 <= 819;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1972: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 724;
        o_index_for_a1 <= 820;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1973: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 725;
        o_index_for_a1 <= 821;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1974: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 726;
        o_index_for_a1 <= 822;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1975: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 727;
        o_index_for_a1 <= 823;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1976: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 728;
        o_index_for_a1 <= 824;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1977: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 729;
        o_index_for_a1 <= 825;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1978: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 730;
        o_index_for_a1 <= 826;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1979: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 731;
        o_index_for_a1 <= 827;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1980: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 732;
        o_index_for_a1 <= 828;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1981: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 733;
        o_index_for_a1 <= 829;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1982: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 734;
        o_index_for_a1 <= 830;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1983: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 735;
        o_index_for_a1 <= 831;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1984: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 736;
        o_index_for_a1 <= 832;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1985: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 737;
        o_index_for_a1 <= 833;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1986: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 738;
        o_index_for_a1 <= 834;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1987: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 739;
        o_index_for_a1 <= 835;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1988: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 740;
        o_index_for_a1 <= 836;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1989: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 741;
        o_index_for_a1 <= 837;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1990: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 742;
        o_index_for_a1 <= 838;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1991: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 743;
        o_index_for_a1 <= 839;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1992: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 744;
        o_index_for_a1 <= 840;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1993: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 745;
        o_index_for_a1 <= 841;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1994: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 746;
        o_index_for_a1 <= 842;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1995: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 747;
        o_index_for_a1 <= 843;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1996: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 748;
        o_index_for_a1 <= 844;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1997: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 749;
        o_index_for_a1 <= 845;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1998: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 750;
        o_index_for_a1 <= 846;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    1999: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 751;
        o_index_for_a1 <= 847;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2000: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 752;
        o_index_for_a1 <= 848;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2001: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 753;
        o_index_for_a1 <= 849;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2002: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 754;
        o_index_for_a1 <= 850;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2003: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 755;
        o_index_for_a1 <= 851;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2004: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 756;
        o_index_for_a1 <= 852;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2005: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 757;
        o_index_for_a1 <= 853;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2006: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 758;
        o_index_for_a1 <= 854;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2007: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 759;
        o_index_for_a1 <= 855;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2008: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 760;
        o_index_for_a1 <= 856;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2009: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 761;
        o_index_for_a1 <= 857;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2010: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 762;
        o_index_for_a1 <= 858;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2011: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 763;
        o_index_for_a1 <= 859;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2012: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 764;
        o_index_for_a1 <= 860;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2013: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 765;
        o_index_for_a1 <= 861;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2014: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 766;
        o_index_for_a1 <= 862;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2015: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 767;
        o_index_for_a1 <= 863;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2016: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 768;
        o_index_for_a1 <= 864;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2017: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 769;
        o_index_for_a1 <= 865;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2018: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 770;
        o_index_for_a1 <= 866;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2019: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 771;
        o_index_for_a1 <= 867;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2020: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 772;
        o_index_for_a1 <= 868;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2021: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 773;
        o_index_for_a1 <= 869;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2022: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 774;
        o_index_for_a1 <= 870;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2023: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 775;
        o_index_for_a1 <= 871;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2024: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 776;
        o_index_for_a1 <= 872;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2025: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 777;
        o_index_for_a1 <= 873;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2026: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 778;
        o_index_for_a1 <= 874;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2027: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 779;
        o_index_for_a1 <= 875;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2028: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 780;
        o_index_for_a1 <= 876;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2029: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 781;
        o_index_for_a1 <= 877;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2030: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 782;
        o_index_for_a1 <= 878;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2031: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 783;
        o_index_for_a1 <= 879;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2032: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 784;
        o_index_for_a1 <= 880;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2033: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 785;
        o_index_for_a1 <= 881;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2034: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 786;
        o_index_for_a1 <= 882;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2035: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 787;
        o_index_for_a1 <= 883;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2036: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 788;
        o_index_for_a1 <= 884;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2037: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 789;
        o_index_for_a1 <= 885;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2038: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 790;
        o_index_for_a1 <= 886;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2039: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 791;
        o_index_for_a1 <= 887;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2040: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 792;
        o_index_for_a1 <= 888;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2041: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 793;
        o_index_for_a1 <= 889;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2042: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 794;
        o_index_for_a1 <= 890;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2043: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 795;
        o_index_for_a1 <= 891;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2044: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 796;
        o_index_for_a1 <= 892;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2045: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 797;
        o_index_for_a1 <= 893;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2046: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 798;
        o_index_for_a1 <= 894;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2047: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 799;
        o_index_for_a1 <= 895;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2048: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 800;
        o_index_for_a1 <= 896;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2049: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 801;
        o_index_for_a1 <= 897;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2050: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 802;
        o_index_for_a1 <= 898;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2051: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 803;
        o_index_for_a1 <= 899;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2052: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 804;
        o_index_for_a1 <= 900;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2053: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 805;
        o_index_for_a1 <= 901;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2054: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 806;
        o_index_for_a1 <= 902;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2055: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 807;
        o_index_for_a1 <= 903;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2056: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 808;
        o_index_for_a1 <= 904;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2057: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 809;
        o_index_for_a1 <= 905;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2058: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 810;
        o_index_for_a1 <= 906;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2059: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 811;
        o_index_for_a1 <= 907;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2060: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 812;
        o_index_for_a1 <= 908;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2061: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 813;
        o_index_for_a1 <= 909;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2062: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 814;
        o_index_for_a1 <= 910;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2063: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 815;
        o_index_for_a1 <= 911;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2064: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 816;
        o_index_for_a1 <= 912;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2065: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 817;
        o_index_for_a1 <= 913;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2066: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 818;
        o_index_for_a1 <= 914;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2067: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 819;
        o_index_for_a1 <= 915;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2068: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 820;
        o_index_for_a1 <= 916;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2069: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 821;
        o_index_for_a1 <= 917;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2070: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 822;
        o_index_for_a1 <= 918;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2071: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 823;
        o_index_for_a1 <= 919;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2072: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 824;
        o_index_for_a1 <= 920;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2073: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 825;
        o_index_for_a1 <= 921;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2074: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 826;
        o_index_for_a1 <= 922;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2075: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 827;
        o_index_for_a1 <= 923;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2076: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 828;
        o_index_for_a1 <= 924;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2077: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 829;
        o_index_for_a1 <= 925;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2078: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 830;
        o_index_for_a1 <= 926;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2079: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 831;
        o_index_for_a1 <= 927;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2080: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 832;
        o_index_for_a1 <= 928;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2081: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 833;
        o_index_for_a1 <= 929;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2082: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 834;
        o_index_for_a1 <= 930;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2083: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 835;
        o_index_for_a1 <= 931;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2084: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 836;
        o_index_for_a1 <= 932;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2085: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 837;
        o_index_for_a1 <= 933;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2086: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 838;
        o_index_for_a1 <= 934;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2087: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 839;
        o_index_for_a1 <= 935;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2088: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 840;
        o_index_for_a1 <= 936;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2089: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 841;
        o_index_for_a1 <= 937;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2090: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 842;
        o_index_for_a1 <= 938;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2091: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 843;
        o_index_for_a1 <= 939;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2092: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 844;
        o_index_for_a1 <= 940;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2093: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 845;
        o_index_for_a1 <= 941;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2094: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 846;
        o_index_for_a1 <= 942;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2095: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 847;
        o_index_for_a1 <= 943;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2096: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 848;
        o_index_for_a1 <= 944;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2097: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 849;
        o_index_for_a1 <= 945;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2098: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 850;
        o_index_for_a1 <= 946;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2099: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 851;
        o_index_for_a1 <= 947;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2100: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 852;
        o_index_for_a1 <= 948;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2101: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 853;
        o_index_for_a1 <= 949;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2102: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 854;
        o_index_for_a1 <= 950;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2103: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 855;
        o_index_for_a1 <= 951;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2104: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 856;
        o_index_for_a1 <= 952;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2105: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 857;
        o_index_for_a1 <= 953;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2106: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 858;
        o_index_for_a1 <= 954;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2107: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 859;
        o_index_for_a1 <= 955;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2108: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 860;
        o_index_for_a1 <= 956;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2109: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 861;
        o_index_for_a1 <= 957;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2110: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 862;
        o_index_for_a1 <= 958;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2111: begin
        o_branch_for_a0 <= 6;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 863;
        o_index_for_a1 <= 959;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2112: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 864;
        o_index_for_a1 <= 960;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2113: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 865;
        o_index_for_a1 <= 961;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2114: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 866;
        o_index_for_a1 <= 962;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2115: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 867;
        o_index_for_a1 <= 963;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2116: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 868;
        o_index_for_a1 <= 964;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2117: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 869;
        o_index_for_a1 <= 965;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2118: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 870;
        o_index_for_a1 <= 966;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2119: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 871;
        o_index_for_a1 <= 967;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2120: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 872;
        o_index_for_a1 <= 968;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2121: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 873;
        o_index_for_a1 <= 969;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2122: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 874;
        o_index_for_a1 <= 970;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2123: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 875;
        o_index_for_a1 <= 971;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2124: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 876;
        o_index_for_a1 <= 972;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2125: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 877;
        o_index_for_a1 <= 973;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2126: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 878;
        o_index_for_a1 <= 974;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2127: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 879;
        o_index_for_a1 <= 975;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2128: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 880;
        o_index_for_a1 <= 976;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2129: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 881;
        o_index_for_a1 <= 977;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2130: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 882;
        o_index_for_a1 <= 978;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2131: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 883;
        o_index_for_a1 <= 979;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2132: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 884;
        o_index_for_a1 <= 980;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2133: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 885;
        o_index_for_a1 <= 981;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2134: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 886;
        o_index_for_a1 <= 982;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2135: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 887;
        o_index_for_a1 <= 983;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2136: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 888;
        o_index_for_a1 <= 984;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2137: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 889;
        o_index_for_a1 <= 985;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2138: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 890;
        o_index_for_a1 <= 986;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2139: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 891;
        o_index_for_a1 <= 987;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2140: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 892;
        o_index_for_a1 <= 988;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2141: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 893;
        o_index_for_a1 <= 989;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2142: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 894;
        o_index_for_a1 <= 990;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2143: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 895;
        o_index_for_a1 <= 991;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2144: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 896;
        o_index_for_a1 <= 992;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2145: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 897;
        o_index_for_a1 <= 993;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2146: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 898;
        o_index_for_a1 <= 994;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2147: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 899;
        o_index_for_a1 <= 995;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2148: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 900;
        o_index_for_a1 <= 996;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2149: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 901;
        o_index_for_a1 <= 997;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2150: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 902;
        o_index_for_a1 <= 998;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2151: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 903;
        o_index_for_a1 <= 999;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2152: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 904;
        o_index_for_a1 <= 1000;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2153: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 905;
        o_index_for_a1 <= 1001;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2154: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 906;
        o_index_for_a1 <= 1002;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2155: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 907;
        o_index_for_a1 <= 1003;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2156: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 908;
        o_index_for_a1 <= 1004;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2157: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 909;
        o_index_for_a1 <= 1005;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2158: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 910;
        o_index_for_a1 <= 1006;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2159: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 911;
        o_index_for_a1 <= 1007;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2160: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 912;
        o_index_for_a1 <= 1008;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2161: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 913;
        o_index_for_a1 <= 1009;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2162: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 914;
        o_index_for_a1 <= 1010;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2163: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 915;
        o_index_for_a1 <= 1011;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2164: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 916;
        o_index_for_a1 <= 1012;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2165: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 917;
        o_index_for_a1 <= 1013;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2166: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 918;
        o_index_for_a1 <= 1014;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2167: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 919;
        o_index_for_a1 <= 1015;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2168: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 920;
        o_index_for_a1 <= 1016;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2169: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 921;
        o_index_for_a1 <= 1017;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2170: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 922;
        o_index_for_a1 <= 1018;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2171: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 923;
        o_index_for_a1 <= 1019;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2172: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 924;
        o_index_for_a1 <= 1020;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2173: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 925;
        o_index_for_a1 <= 1021;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2174: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 926;
        o_index_for_a1 <= 1022;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2175: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 927;
        o_index_for_a1 <= 1023;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2176: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 928;
        o_index_for_a1 <= 1024;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2177: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 929;
        o_index_for_a1 <= 1025;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2178: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 930;
        o_index_for_a1 <= 1026;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2179: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 931;
        o_index_for_a1 <= 1027;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2180: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 932;
        o_index_for_a1 <= 1028;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2181: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 933;
        o_index_for_a1 <= 1029;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2182: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 934;
        o_index_for_a1 <= 1030;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2183: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 935;
        o_index_for_a1 <= 1031;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2184: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 936;
        o_index_for_a1 <= 1032;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2185: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 937;
        o_index_for_a1 <= 1033;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2186: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 938;
        o_index_for_a1 <= 1034;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2187: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 939;
        o_index_for_a1 <= 1035;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2188: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 940;
        o_index_for_a1 <= 1036;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2189: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 941;
        o_index_for_a1 <= 1037;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2190: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 942;
        o_index_for_a1 <= 1038;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2191: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 943;
        o_index_for_a1 <= 1039;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2192: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 944;
        o_index_for_a1 <= 1040;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2193: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 945;
        o_index_for_a1 <= 1041;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2194: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 946;
        o_index_for_a1 <= 1042;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2195: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 947;
        o_index_for_a1 <= 1043;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2196: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 948;
        o_index_for_a1 <= 1044;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2197: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 949;
        o_index_for_a1 <= 1045;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2198: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 950;
        o_index_for_a1 <= 1046;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2199: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 951;
        o_index_for_a1 <= 1047;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2200: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 952;
        o_index_for_a1 <= 1048;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2201: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 953;
        o_index_for_a1 <= 1049;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2202: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 954;
        o_index_for_a1 <= 1050;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2203: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 955;
        o_index_for_a1 <= 1051;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2204: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 956;
        o_index_for_a1 <= 1052;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2205: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 957;
        o_index_for_a1 <= 1053;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2206: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 958;
        o_index_for_a1 <= 1054;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2207: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 959;
        o_index_for_a1 <= 1055;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2208: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 960;
        o_index_for_a1 <= 1056;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2209: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 961;
        o_index_for_a1 <= 1057;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2210: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 962;
        o_index_for_a1 <= 1058;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2211: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 963;
        o_index_for_a1 <= 1059;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2212: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 964;
        o_index_for_a1 <= 1060;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2213: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 965;
        o_index_for_a1 <= 1061;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2214: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 966;
        o_index_for_a1 <= 1062;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2215: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 967;
        o_index_for_a1 <= 1063;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2216: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 968;
        o_index_for_a1 <= 1064;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2217: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 969;
        o_index_for_a1 <= 1065;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2218: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 970;
        o_index_for_a1 <= 1066;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2219: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 971;
        o_index_for_a1 <= 1067;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2220: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 972;
        o_index_for_a1 <= 1068;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2221: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 973;
        o_index_for_a1 <= 1069;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2222: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 974;
        o_index_for_a1 <= 1070;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2223: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 975;
        o_index_for_a1 <= 1071;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2224: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 976;
        o_index_for_a1 <= 1072;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2225: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 977;
        o_index_for_a1 <= 1073;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2226: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 978;
        o_index_for_a1 <= 1074;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2227: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 979;
        o_index_for_a1 <= 1075;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2228: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 980;
        o_index_for_a1 <= 1076;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2229: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 981;
        o_index_for_a1 <= 1077;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2230: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 982;
        o_index_for_a1 <= 1078;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2231: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 983;
        o_index_for_a1 <= 1079;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2232: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 984;
        o_index_for_a1 <= 1080;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2233: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 985;
        o_index_for_a1 <= 1081;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2234: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 986;
        o_index_for_a1 <= 1082;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2235: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 987;
        o_index_for_a1 <= 1083;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2236: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 988;
        o_index_for_a1 <= 1084;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2237: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 989;
        o_index_for_a1 <= 1085;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2238: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 990;
        o_index_for_a1 <= 1086;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2239: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 991;
        o_index_for_a1 <= 1087;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2240: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 992;
        o_index_for_a1 <= 1088;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2241: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 993;
        o_index_for_a1 <= 1089;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2242: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 994;
        o_index_for_a1 <= 1090;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2243: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 995;
        o_index_for_a1 <= 1091;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2244: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 996;
        o_index_for_a1 <= 1092;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2245: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 997;
        o_index_for_a1 <= 1093;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2246: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 998;
        o_index_for_a1 <= 1094;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2247: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 999;
        o_index_for_a1 <= 1095;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2248: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1000;
        o_index_for_a1 <= 1096;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2249: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1001;
        o_index_for_a1 <= 1097;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2250: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1002;
        o_index_for_a1 <= 1098;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2251: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1003;
        o_index_for_a1 <= 1099;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2252: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1004;
        o_index_for_a1 <= 1100;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2253: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1005;
        o_index_for_a1 <= 1101;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2254: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1006;
        o_index_for_a1 <= 1102;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2255: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1007;
        o_index_for_a1 <= 1103;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2256: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1008;
        o_index_for_a1 <= 1104;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2257: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1009;
        o_index_for_a1 <= 1105;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2258: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1010;
        o_index_for_a1 <= 1106;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2259: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1011;
        o_index_for_a1 <= 1107;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2260: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1012;
        o_index_for_a1 <= 1108;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2261: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1013;
        o_index_for_a1 <= 1109;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2262: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1014;
        o_index_for_a1 <= 1110;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2263: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1015;
        o_index_for_a1 <= 1111;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2264: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1016;
        o_index_for_a1 <= 1112;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2265: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1017;
        o_index_for_a1 <= 1113;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2266: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1018;
        o_index_for_a1 <= 1114;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2267: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1019;
        o_index_for_a1 <= 1115;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2268: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1020;
        o_index_for_a1 <= 1116;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2269: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1021;
        o_index_for_a1 <= 1117;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2270: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1022;
        o_index_for_a1 <= 1118;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2271: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1023;
        o_index_for_a1 <= 1119;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2272: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1024;
        o_index_for_a1 <= 1120;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2273: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1025;
        o_index_for_a1 <= 1121;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2274: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1026;
        o_index_for_a1 <= 1122;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2275: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1027;
        o_index_for_a1 <= 1123;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2276: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1028;
        o_index_for_a1 <= 1124;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2277: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1029;
        o_index_for_a1 <= 1125;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2278: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1030;
        o_index_for_a1 <= 1126;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2279: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1031;
        o_index_for_a1 <= 1127;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2280: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1032;
        o_index_for_a1 <= 1128;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2281: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1033;
        o_index_for_a1 <= 1129;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2282: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1034;
        o_index_for_a1 <= 1130;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2283: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1035;
        o_index_for_a1 <= 1131;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2284: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1036;
        o_index_for_a1 <= 1132;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2285: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1037;
        o_index_for_a1 <= 1133;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2286: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1038;
        o_index_for_a1 <= 1134;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2287: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1039;
        o_index_for_a1 <= 1135;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2288: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1040;
        o_index_for_a1 <= 1136;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2289: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1041;
        o_index_for_a1 <= 1137;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2290: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1042;
        o_index_for_a1 <= 1138;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2291: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1043;
        o_index_for_a1 <= 1139;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2292: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1044;
        o_index_for_a1 <= 1140;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2293: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1045;
        o_index_for_a1 <= 1141;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2294: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1046;
        o_index_for_a1 <= 1142;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2295: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1047;
        o_index_for_a1 <= 1143;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2296: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1048;
        o_index_for_a1 <= 1144;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2297: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1049;
        o_index_for_a1 <= 1145;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2298: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1050;
        o_index_for_a1 <= 1146;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2299: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1051;
        o_index_for_a1 <= 1147;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2300: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1052;
        o_index_for_a1 <= 1148;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2301: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1053;
        o_index_for_a1 <= 1149;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2302: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1054;
        o_index_for_a1 <= 1150;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    2303: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 7;
        o_branch_for_a3 <= 7;
        o_branch_for_a4 <= 7;
        o_branch_for_a5 <= 7; 
        o_index_for_a0 <= 1055;
        o_index_for_a1 <= 1151;
        o_index_for_a2 <= 1152;
        o_index_for_a3 <= 1152;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1152; 
    end
    default: begin // This case is for simulation purposes only.
        o_branch_for_a0 <= 'x;
        o_branch_for_a1 <= 'x;
        o_branch_for_a2 <= 'x;
        o_branch_for_a3 <= 'x;
        o_branch_for_a4 <= 'x;
        o_branch_for_a5 <= 'x; 
        o_index_for_a0 <= 'x;
        o_index_for_a1 <= 'x;
        o_index_for_a2 <= 'x;
        o_index_for_a3 <= 'x;
        o_index_for_a4 <= 'x;
        o_index_for_a5 <= 'x; 
    end
    endcase
end

endmodule: ldpc_column_to_row_rom

`default_nettype wire
