// Generated from template at 01/31/2017
`timescale 10ps / 10ps

`default_nettype none

module ldpc_row_to_column_rom #(
	parameter integer INPUT_LENGTH = 2304,
    parameter integer EXPANSION_FACTOR = 96
) (
    input  wire logic                                   i_valid,
    output      logic [$clog2(24*EXPANSION_FACTOR)-1:0] o_index_for_a0,
    output      logic [$clog2(24*EXPANSION_FACTOR)-1:0] o_index_for_a1,
    output      logic [$clog2(24*EXPANSION_FACTOR)-1:0] o_index_for_a2,
    output      logic [$clog2(24*EXPANSION_FACTOR)-1:0] o_index_for_a3,
    output      logic [$clog2(24*EXPANSION_FACTOR)-1:0] o_index_for_a4,
    output      logic [$clog2(24*EXPANSION_FACTOR)-1:0] o_index_for_a5,
    output      logic [$clog2(24*EXPANSION_FACTOR)-1:0] o_index_for_a6, 
    output      logic [$clog2(8)-1:0]                   o_branch_for_a0,
    output      logic [$clog2(8)-1:0]                   o_branch_for_a1,
    output      logic [$clog2(8)-1:0]                   o_branch_for_a2,
    output      logic [$clog2(8)-1:0]                   o_branch_for_a3,
    output      logic [$clog2(8)-1:0]                   o_branch_for_a4,
    output      logic [$clog2(8)-1:0]                   o_branch_for_a5,
    output      logic [$clog2(8)-1:0]                   o_branch_for_a6,
    input  wire logic                                   i_clock,
	input  wire logic                                   i_reset
);

logic [$clog2(INPUT_LENGTH)-1:0] count;

always_ff @(posedge i_clock) begin
    if (i_reset == 1'b1) begin
        count <= 0;
    end else if (i_valid) begin
        if (count == INPUT_LENGTH-1) begin
            count <= 0;
        end else begin
            count <= count + 1;
        end
    end

    case (count)
    0: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 98;
        o_index_for_a1 <= 215;
        o_index_for_a2 <= 809;
        o_index_for_a3 <= 877;
        o_index_for_a4 <= 1241;
        o_index_for_a5 <= 1248; 
        o_index_for_a6 <= 2304; 
    end
    1: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 99;
        o_index_for_a1 <= 216;
        o_index_for_a2 <= 810;
        o_index_for_a3 <= 878;
        o_index_for_a4 <= 1242;
        o_index_for_a5 <= 1249; 
        o_index_for_a6 <= 2304; 
    end
    2: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 100;
        o_index_for_a1 <= 217;
        o_index_for_a2 <= 811;
        o_index_for_a3 <= 879;
        o_index_for_a4 <= 1243;
        o_index_for_a5 <= 1250; 
        o_index_for_a6 <= 2304; 
    end
    3: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 101;
        o_index_for_a1 <= 218;
        o_index_for_a2 <= 812;
        o_index_for_a3 <= 880;
        o_index_for_a4 <= 1244;
        o_index_for_a5 <= 1251; 
        o_index_for_a6 <= 2304; 
    end
    4: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 102;
        o_index_for_a1 <= 219;
        o_index_for_a2 <= 813;
        o_index_for_a3 <= 881;
        o_index_for_a4 <= 1245;
        o_index_for_a5 <= 1252; 
        o_index_for_a6 <= 2304; 
    end
    5: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 103;
        o_index_for_a1 <= 220;
        o_index_for_a2 <= 814;
        o_index_for_a3 <= 882;
        o_index_for_a4 <= 1246;
        o_index_for_a5 <= 1253; 
        o_index_for_a6 <= 2304; 
    end
    6: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 104;
        o_index_for_a1 <= 221;
        o_index_for_a2 <= 815;
        o_index_for_a3 <= 883;
        o_index_for_a4 <= 1247;
        o_index_for_a5 <= 1254; 
        o_index_for_a6 <= 2304; 
    end
    7: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 105;
        o_index_for_a1 <= 222;
        o_index_for_a2 <= 816;
        o_index_for_a3 <= 884;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1255; 
        o_index_for_a6 <= 2304; 
    end
    8: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 106;
        o_index_for_a1 <= 223;
        o_index_for_a2 <= 817;
        o_index_for_a3 <= 885;
        o_index_for_a4 <= 1153;
        o_index_for_a5 <= 1256; 
        o_index_for_a6 <= 2304; 
    end
    9: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 107;
        o_index_for_a1 <= 224;
        o_index_for_a2 <= 818;
        o_index_for_a3 <= 886;
        o_index_for_a4 <= 1154;
        o_index_for_a5 <= 1257; 
        o_index_for_a6 <= 2304; 
    end
    10: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 108;
        o_index_for_a1 <= 225;
        o_index_for_a2 <= 819;
        o_index_for_a3 <= 887;
        o_index_for_a4 <= 1155;
        o_index_for_a5 <= 1258; 
        o_index_for_a6 <= 2304; 
    end
    11: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 109;
        o_index_for_a1 <= 226;
        o_index_for_a2 <= 820;
        o_index_for_a3 <= 888;
        o_index_for_a4 <= 1156;
        o_index_for_a5 <= 1259; 
        o_index_for_a6 <= 2304; 
    end
    12: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 110;
        o_index_for_a1 <= 227;
        o_index_for_a2 <= 821;
        o_index_for_a3 <= 889;
        o_index_for_a4 <= 1157;
        o_index_for_a5 <= 1260; 
        o_index_for_a6 <= 2304; 
    end
    13: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 111;
        o_index_for_a1 <= 228;
        o_index_for_a2 <= 822;
        o_index_for_a3 <= 890;
        o_index_for_a4 <= 1158;
        o_index_for_a5 <= 1261; 
        o_index_for_a6 <= 2304; 
    end
    14: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 112;
        o_index_for_a1 <= 229;
        o_index_for_a2 <= 823;
        o_index_for_a3 <= 891;
        o_index_for_a4 <= 1159;
        o_index_for_a5 <= 1262; 
        o_index_for_a6 <= 2304; 
    end
    15: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 113;
        o_index_for_a1 <= 230;
        o_index_for_a2 <= 824;
        o_index_for_a3 <= 892;
        o_index_for_a4 <= 1160;
        o_index_for_a5 <= 1263; 
        o_index_for_a6 <= 2304; 
    end
    16: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 114;
        o_index_for_a1 <= 231;
        o_index_for_a2 <= 825;
        o_index_for_a3 <= 893;
        o_index_for_a4 <= 1161;
        o_index_for_a5 <= 1264; 
        o_index_for_a6 <= 2304; 
    end
    17: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 115;
        o_index_for_a1 <= 232;
        o_index_for_a2 <= 826;
        o_index_for_a3 <= 894;
        o_index_for_a4 <= 1162;
        o_index_for_a5 <= 1265; 
        o_index_for_a6 <= 2304; 
    end
    18: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 116;
        o_index_for_a1 <= 233;
        o_index_for_a2 <= 827;
        o_index_for_a3 <= 895;
        o_index_for_a4 <= 1163;
        o_index_for_a5 <= 1266; 
        o_index_for_a6 <= 2304; 
    end
    19: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 117;
        o_index_for_a1 <= 234;
        o_index_for_a2 <= 828;
        o_index_for_a3 <= 896;
        o_index_for_a4 <= 1164;
        o_index_for_a5 <= 1267; 
        o_index_for_a6 <= 2304; 
    end
    20: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 118;
        o_index_for_a1 <= 235;
        o_index_for_a2 <= 829;
        o_index_for_a3 <= 897;
        o_index_for_a4 <= 1165;
        o_index_for_a5 <= 1268; 
        o_index_for_a6 <= 2304; 
    end
    21: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 119;
        o_index_for_a1 <= 236;
        o_index_for_a2 <= 830;
        o_index_for_a3 <= 898;
        o_index_for_a4 <= 1166;
        o_index_for_a5 <= 1269; 
        o_index_for_a6 <= 2304; 
    end
    22: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 120;
        o_index_for_a1 <= 237;
        o_index_for_a2 <= 831;
        o_index_for_a3 <= 899;
        o_index_for_a4 <= 1167;
        o_index_for_a5 <= 1270; 
        o_index_for_a6 <= 2304; 
    end
    23: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 121;
        o_index_for_a1 <= 238;
        o_index_for_a2 <= 832;
        o_index_for_a3 <= 900;
        o_index_for_a4 <= 1168;
        o_index_for_a5 <= 1271; 
        o_index_for_a6 <= 2304; 
    end
    24: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 122;
        o_index_for_a1 <= 239;
        o_index_for_a2 <= 833;
        o_index_for_a3 <= 901;
        o_index_for_a4 <= 1169;
        o_index_for_a5 <= 1272; 
        o_index_for_a6 <= 2304; 
    end
    25: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 123;
        o_index_for_a1 <= 240;
        o_index_for_a2 <= 834;
        o_index_for_a3 <= 902;
        o_index_for_a4 <= 1170;
        o_index_for_a5 <= 1273; 
        o_index_for_a6 <= 2304; 
    end
    26: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 124;
        o_index_for_a1 <= 241;
        o_index_for_a2 <= 835;
        o_index_for_a3 <= 903;
        o_index_for_a4 <= 1171;
        o_index_for_a5 <= 1274; 
        o_index_for_a6 <= 2304; 
    end
    27: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 125;
        o_index_for_a1 <= 242;
        o_index_for_a2 <= 836;
        o_index_for_a3 <= 904;
        o_index_for_a4 <= 1172;
        o_index_for_a5 <= 1275; 
        o_index_for_a6 <= 2304; 
    end
    28: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 126;
        o_index_for_a1 <= 243;
        o_index_for_a2 <= 837;
        o_index_for_a3 <= 905;
        o_index_for_a4 <= 1173;
        o_index_for_a5 <= 1276; 
        o_index_for_a6 <= 2304; 
    end
    29: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 127;
        o_index_for_a1 <= 244;
        o_index_for_a2 <= 838;
        o_index_for_a3 <= 906;
        o_index_for_a4 <= 1174;
        o_index_for_a5 <= 1277; 
        o_index_for_a6 <= 2304; 
    end
    30: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 128;
        o_index_for_a1 <= 245;
        o_index_for_a2 <= 839;
        o_index_for_a3 <= 907;
        o_index_for_a4 <= 1175;
        o_index_for_a5 <= 1278; 
        o_index_for_a6 <= 2304; 
    end
    31: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 129;
        o_index_for_a1 <= 246;
        o_index_for_a2 <= 840;
        o_index_for_a3 <= 908;
        o_index_for_a4 <= 1176;
        o_index_for_a5 <= 1279; 
        o_index_for_a6 <= 2304; 
    end
    32: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 130;
        o_index_for_a1 <= 247;
        o_index_for_a2 <= 841;
        o_index_for_a3 <= 909;
        o_index_for_a4 <= 1177;
        o_index_for_a5 <= 1280; 
        o_index_for_a6 <= 2304; 
    end
    33: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 131;
        o_index_for_a1 <= 248;
        o_index_for_a2 <= 842;
        o_index_for_a3 <= 910;
        o_index_for_a4 <= 1178;
        o_index_for_a5 <= 1281; 
        o_index_for_a6 <= 2304; 
    end
    34: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 132;
        o_index_for_a1 <= 249;
        o_index_for_a2 <= 843;
        o_index_for_a3 <= 911;
        o_index_for_a4 <= 1179;
        o_index_for_a5 <= 1282; 
        o_index_for_a6 <= 2304; 
    end
    35: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 133;
        o_index_for_a1 <= 250;
        o_index_for_a2 <= 844;
        o_index_for_a3 <= 912;
        o_index_for_a4 <= 1180;
        o_index_for_a5 <= 1283; 
        o_index_for_a6 <= 2304; 
    end
    36: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 134;
        o_index_for_a1 <= 251;
        o_index_for_a2 <= 845;
        o_index_for_a3 <= 913;
        o_index_for_a4 <= 1181;
        o_index_for_a5 <= 1284; 
        o_index_for_a6 <= 2304; 
    end
    37: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 135;
        o_index_for_a1 <= 252;
        o_index_for_a2 <= 846;
        o_index_for_a3 <= 914;
        o_index_for_a4 <= 1182;
        o_index_for_a5 <= 1285; 
        o_index_for_a6 <= 2304; 
    end
    38: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 136;
        o_index_for_a1 <= 253;
        o_index_for_a2 <= 847;
        o_index_for_a3 <= 915;
        o_index_for_a4 <= 1183;
        o_index_for_a5 <= 1286; 
        o_index_for_a6 <= 2304; 
    end
    39: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 137;
        o_index_for_a1 <= 254;
        o_index_for_a2 <= 848;
        o_index_for_a3 <= 916;
        o_index_for_a4 <= 1184;
        o_index_for_a5 <= 1287; 
        o_index_for_a6 <= 2304; 
    end
    40: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 138;
        o_index_for_a1 <= 255;
        o_index_for_a2 <= 849;
        o_index_for_a3 <= 917;
        o_index_for_a4 <= 1185;
        o_index_for_a5 <= 1288; 
        o_index_for_a6 <= 2304; 
    end
    41: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 139;
        o_index_for_a1 <= 256;
        o_index_for_a2 <= 850;
        o_index_for_a3 <= 918;
        o_index_for_a4 <= 1186;
        o_index_for_a5 <= 1289; 
        o_index_for_a6 <= 2304; 
    end
    42: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 140;
        o_index_for_a1 <= 257;
        o_index_for_a2 <= 851;
        o_index_for_a3 <= 919;
        o_index_for_a4 <= 1187;
        o_index_for_a5 <= 1290; 
        o_index_for_a6 <= 2304; 
    end
    43: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 141;
        o_index_for_a1 <= 258;
        o_index_for_a2 <= 852;
        o_index_for_a3 <= 920;
        o_index_for_a4 <= 1188;
        o_index_for_a5 <= 1291; 
        o_index_for_a6 <= 2304; 
    end
    44: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 142;
        o_index_for_a1 <= 259;
        o_index_for_a2 <= 853;
        o_index_for_a3 <= 921;
        o_index_for_a4 <= 1189;
        o_index_for_a5 <= 1292; 
        o_index_for_a6 <= 2304; 
    end
    45: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 143;
        o_index_for_a1 <= 260;
        o_index_for_a2 <= 854;
        o_index_for_a3 <= 922;
        o_index_for_a4 <= 1190;
        o_index_for_a5 <= 1293; 
        o_index_for_a6 <= 2304; 
    end
    46: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 144;
        o_index_for_a1 <= 261;
        o_index_for_a2 <= 855;
        o_index_for_a3 <= 923;
        o_index_for_a4 <= 1191;
        o_index_for_a5 <= 1294; 
        o_index_for_a6 <= 2304; 
    end
    47: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 145;
        o_index_for_a1 <= 262;
        o_index_for_a2 <= 856;
        o_index_for_a3 <= 924;
        o_index_for_a4 <= 1192;
        o_index_for_a5 <= 1295; 
        o_index_for_a6 <= 2304; 
    end
    48: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 146;
        o_index_for_a1 <= 263;
        o_index_for_a2 <= 857;
        o_index_for_a3 <= 925;
        o_index_for_a4 <= 1193;
        o_index_for_a5 <= 1296; 
        o_index_for_a6 <= 2304; 
    end
    49: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 147;
        o_index_for_a1 <= 264;
        o_index_for_a2 <= 858;
        o_index_for_a3 <= 926;
        o_index_for_a4 <= 1194;
        o_index_for_a5 <= 1297; 
        o_index_for_a6 <= 2304; 
    end
    50: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 148;
        o_index_for_a1 <= 265;
        o_index_for_a2 <= 859;
        o_index_for_a3 <= 927;
        o_index_for_a4 <= 1195;
        o_index_for_a5 <= 1298; 
        o_index_for_a6 <= 2304; 
    end
    51: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 149;
        o_index_for_a1 <= 266;
        o_index_for_a2 <= 860;
        o_index_for_a3 <= 928;
        o_index_for_a4 <= 1196;
        o_index_for_a5 <= 1299; 
        o_index_for_a6 <= 2304; 
    end
    52: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 150;
        o_index_for_a1 <= 267;
        o_index_for_a2 <= 861;
        o_index_for_a3 <= 929;
        o_index_for_a4 <= 1197;
        o_index_for_a5 <= 1300; 
        o_index_for_a6 <= 2304; 
    end
    53: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 151;
        o_index_for_a1 <= 268;
        o_index_for_a2 <= 862;
        o_index_for_a3 <= 930;
        o_index_for_a4 <= 1198;
        o_index_for_a5 <= 1301; 
        o_index_for_a6 <= 2304; 
    end
    54: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 152;
        o_index_for_a1 <= 269;
        o_index_for_a2 <= 863;
        o_index_for_a3 <= 931;
        o_index_for_a4 <= 1199;
        o_index_for_a5 <= 1302; 
        o_index_for_a6 <= 2304; 
    end
    55: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 153;
        o_index_for_a1 <= 270;
        o_index_for_a2 <= 768;
        o_index_for_a3 <= 932;
        o_index_for_a4 <= 1200;
        o_index_for_a5 <= 1303; 
        o_index_for_a6 <= 2304; 
    end
    56: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 154;
        o_index_for_a1 <= 271;
        o_index_for_a2 <= 769;
        o_index_for_a3 <= 933;
        o_index_for_a4 <= 1201;
        o_index_for_a5 <= 1304; 
        o_index_for_a6 <= 2304; 
    end
    57: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 155;
        o_index_for_a1 <= 272;
        o_index_for_a2 <= 770;
        o_index_for_a3 <= 934;
        o_index_for_a4 <= 1202;
        o_index_for_a5 <= 1305; 
        o_index_for_a6 <= 2304; 
    end
    58: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 156;
        o_index_for_a1 <= 273;
        o_index_for_a2 <= 771;
        o_index_for_a3 <= 935;
        o_index_for_a4 <= 1203;
        o_index_for_a5 <= 1306; 
        o_index_for_a6 <= 2304; 
    end
    59: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 157;
        o_index_for_a1 <= 274;
        o_index_for_a2 <= 772;
        o_index_for_a3 <= 936;
        o_index_for_a4 <= 1204;
        o_index_for_a5 <= 1307; 
        o_index_for_a6 <= 2304; 
    end
    60: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 158;
        o_index_for_a1 <= 275;
        o_index_for_a2 <= 773;
        o_index_for_a3 <= 937;
        o_index_for_a4 <= 1205;
        o_index_for_a5 <= 1308; 
        o_index_for_a6 <= 2304; 
    end
    61: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 159;
        o_index_for_a1 <= 276;
        o_index_for_a2 <= 774;
        o_index_for_a3 <= 938;
        o_index_for_a4 <= 1206;
        o_index_for_a5 <= 1309; 
        o_index_for_a6 <= 2304; 
    end
    62: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 160;
        o_index_for_a1 <= 277;
        o_index_for_a2 <= 775;
        o_index_for_a3 <= 939;
        o_index_for_a4 <= 1207;
        o_index_for_a5 <= 1310; 
        o_index_for_a6 <= 2304; 
    end
    63: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 161;
        o_index_for_a1 <= 278;
        o_index_for_a2 <= 776;
        o_index_for_a3 <= 940;
        o_index_for_a4 <= 1208;
        o_index_for_a5 <= 1311; 
        o_index_for_a6 <= 2304; 
    end
    64: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 162;
        o_index_for_a1 <= 279;
        o_index_for_a2 <= 777;
        o_index_for_a3 <= 941;
        o_index_for_a4 <= 1209;
        o_index_for_a5 <= 1312; 
        o_index_for_a6 <= 2304; 
    end
    65: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 163;
        o_index_for_a1 <= 280;
        o_index_for_a2 <= 778;
        o_index_for_a3 <= 942;
        o_index_for_a4 <= 1210;
        o_index_for_a5 <= 1313; 
        o_index_for_a6 <= 2304; 
    end
    66: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 164;
        o_index_for_a1 <= 281;
        o_index_for_a2 <= 779;
        o_index_for_a3 <= 943;
        o_index_for_a4 <= 1211;
        o_index_for_a5 <= 1314; 
        o_index_for_a6 <= 2304; 
    end
    67: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 165;
        o_index_for_a1 <= 282;
        o_index_for_a2 <= 780;
        o_index_for_a3 <= 944;
        o_index_for_a4 <= 1212;
        o_index_for_a5 <= 1315; 
        o_index_for_a6 <= 2304; 
    end
    68: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 166;
        o_index_for_a1 <= 283;
        o_index_for_a2 <= 781;
        o_index_for_a3 <= 945;
        o_index_for_a4 <= 1213;
        o_index_for_a5 <= 1316; 
        o_index_for_a6 <= 2304; 
    end
    69: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 167;
        o_index_for_a1 <= 284;
        o_index_for_a2 <= 782;
        o_index_for_a3 <= 946;
        o_index_for_a4 <= 1214;
        o_index_for_a5 <= 1317; 
        o_index_for_a6 <= 2304; 
    end
    70: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 168;
        o_index_for_a1 <= 285;
        o_index_for_a2 <= 783;
        o_index_for_a3 <= 947;
        o_index_for_a4 <= 1215;
        o_index_for_a5 <= 1318; 
        o_index_for_a6 <= 2304; 
    end
    71: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 169;
        o_index_for_a1 <= 286;
        o_index_for_a2 <= 784;
        o_index_for_a3 <= 948;
        o_index_for_a4 <= 1216;
        o_index_for_a5 <= 1319; 
        o_index_for_a6 <= 2304; 
    end
    72: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 170;
        o_index_for_a1 <= 287;
        o_index_for_a2 <= 785;
        o_index_for_a3 <= 949;
        o_index_for_a4 <= 1217;
        o_index_for_a5 <= 1320; 
        o_index_for_a6 <= 2304; 
    end
    73: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 171;
        o_index_for_a1 <= 192;
        o_index_for_a2 <= 786;
        o_index_for_a3 <= 950;
        o_index_for_a4 <= 1218;
        o_index_for_a5 <= 1321; 
        o_index_for_a6 <= 2304; 
    end
    74: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 172;
        o_index_for_a1 <= 193;
        o_index_for_a2 <= 787;
        o_index_for_a3 <= 951;
        o_index_for_a4 <= 1219;
        o_index_for_a5 <= 1322; 
        o_index_for_a6 <= 2304; 
    end
    75: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 173;
        o_index_for_a1 <= 194;
        o_index_for_a2 <= 788;
        o_index_for_a3 <= 952;
        o_index_for_a4 <= 1220;
        o_index_for_a5 <= 1323; 
        o_index_for_a6 <= 2304; 
    end
    76: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 174;
        o_index_for_a1 <= 195;
        o_index_for_a2 <= 789;
        o_index_for_a3 <= 953;
        o_index_for_a4 <= 1221;
        o_index_for_a5 <= 1324; 
        o_index_for_a6 <= 2304; 
    end
    77: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 175;
        o_index_for_a1 <= 196;
        o_index_for_a2 <= 790;
        o_index_for_a3 <= 954;
        o_index_for_a4 <= 1222;
        o_index_for_a5 <= 1325; 
        o_index_for_a6 <= 2304; 
    end
    78: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 176;
        o_index_for_a1 <= 197;
        o_index_for_a2 <= 791;
        o_index_for_a3 <= 955;
        o_index_for_a4 <= 1223;
        o_index_for_a5 <= 1326; 
        o_index_for_a6 <= 2304; 
    end
    79: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 177;
        o_index_for_a1 <= 198;
        o_index_for_a2 <= 792;
        o_index_for_a3 <= 956;
        o_index_for_a4 <= 1224;
        o_index_for_a5 <= 1327; 
        o_index_for_a6 <= 2304; 
    end
    80: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 178;
        o_index_for_a1 <= 199;
        o_index_for_a2 <= 793;
        o_index_for_a3 <= 957;
        o_index_for_a4 <= 1225;
        o_index_for_a5 <= 1328; 
        o_index_for_a6 <= 2304; 
    end
    81: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 179;
        o_index_for_a1 <= 200;
        o_index_for_a2 <= 794;
        o_index_for_a3 <= 958;
        o_index_for_a4 <= 1226;
        o_index_for_a5 <= 1329; 
        o_index_for_a6 <= 2304; 
    end
    82: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 180;
        o_index_for_a1 <= 201;
        o_index_for_a2 <= 795;
        o_index_for_a3 <= 959;
        o_index_for_a4 <= 1227;
        o_index_for_a5 <= 1330; 
        o_index_for_a6 <= 2304; 
    end
    83: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 181;
        o_index_for_a1 <= 202;
        o_index_for_a2 <= 796;
        o_index_for_a3 <= 864;
        o_index_for_a4 <= 1228;
        o_index_for_a5 <= 1331; 
        o_index_for_a6 <= 2304; 
    end
    84: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 182;
        o_index_for_a1 <= 203;
        o_index_for_a2 <= 797;
        o_index_for_a3 <= 865;
        o_index_for_a4 <= 1229;
        o_index_for_a5 <= 1332; 
        o_index_for_a6 <= 2304; 
    end
    85: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 183;
        o_index_for_a1 <= 204;
        o_index_for_a2 <= 798;
        o_index_for_a3 <= 866;
        o_index_for_a4 <= 1230;
        o_index_for_a5 <= 1333; 
        o_index_for_a6 <= 2304; 
    end
    86: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 184;
        o_index_for_a1 <= 205;
        o_index_for_a2 <= 799;
        o_index_for_a3 <= 867;
        o_index_for_a4 <= 1231;
        o_index_for_a5 <= 1334; 
        o_index_for_a6 <= 2304; 
    end
    87: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 185;
        o_index_for_a1 <= 206;
        o_index_for_a2 <= 800;
        o_index_for_a3 <= 868;
        o_index_for_a4 <= 1232;
        o_index_for_a5 <= 1335; 
        o_index_for_a6 <= 2304; 
    end
    88: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 186;
        o_index_for_a1 <= 207;
        o_index_for_a2 <= 801;
        o_index_for_a3 <= 869;
        o_index_for_a4 <= 1233;
        o_index_for_a5 <= 1336; 
        o_index_for_a6 <= 2304; 
    end
    89: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 187;
        o_index_for_a1 <= 208;
        o_index_for_a2 <= 802;
        o_index_for_a3 <= 870;
        o_index_for_a4 <= 1234;
        o_index_for_a5 <= 1337; 
        o_index_for_a6 <= 2304; 
    end
    90: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 188;
        o_index_for_a1 <= 209;
        o_index_for_a2 <= 803;
        o_index_for_a3 <= 871;
        o_index_for_a4 <= 1235;
        o_index_for_a5 <= 1338; 
        o_index_for_a6 <= 2304; 
    end
    91: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 189;
        o_index_for_a1 <= 210;
        o_index_for_a2 <= 804;
        o_index_for_a3 <= 872;
        o_index_for_a4 <= 1236;
        o_index_for_a5 <= 1339; 
        o_index_for_a6 <= 2304; 
    end
    92: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 190;
        o_index_for_a1 <= 211;
        o_index_for_a2 <= 805;
        o_index_for_a3 <= 873;
        o_index_for_a4 <= 1237;
        o_index_for_a5 <= 1340; 
        o_index_for_a6 <= 2304; 
    end
    93: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 191;
        o_index_for_a1 <= 212;
        o_index_for_a2 <= 806;
        o_index_for_a3 <= 874;
        o_index_for_a4 <= 1238;
        o_index_for_a5 <= 1341; 
        o_index_for_a6 <= 2304; 
    end
    94: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 96;
        o_index_for_a1 <= 213;
        o_index_for_a2 <= 807;
        o_index_for_a3 <= 875;
        o_index_for_a4 <= 1239;
        o_index_for_a5 <= 1342; 
        o_index_for_a6 <= 2304; 
    end
    95: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 97;
        o_index_for_a1 <= 214;
        o_index_for_a2 <= 808;
        o_index_for_a3 <= 876;
        o_index_for_a4 <= 1240;
        o_index_for_a5 <= 1343; 
        o_index_for_a6 <= 2304; 
    end
    96: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 165;
        o_index_for_a1 <= 554;
        o_index_for_a2 <= 593;
        o_index_for_a3 <= 759;
        o_index_for_a4 <= 1140;
        o_index_for_a5 <= 1248; 
        o_index_for_a6 <= 1344; 
    end
    97: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 166;
        o_index_for_a1 <= 555;
        o_index_for_a2 <= 594;
        o_index_for_a3 <= 760;
        o_index_for_a4 <= 1141;
        o_index_for_a5 <= 1249; 
        o_index_for_a6 <= 1345; 
    end
    98: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 167;
        o_index_for_a1 <= 556;
        o_index_for_a2 <= 595;
        o_index_for_a3 <= 761;
        o_index_for_a4 <= 1142;
        o_index_for_a5 <= 1250; 
        o_index_for_a6 <= 1346; 
    end
    99: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 168;
        o_index_for_a1 <= 557;
        o_index_for_a2 <= 596;
        o_index_for_a3 <= 762;
        o_index_for_a4 <= 1143;
        o_index_for_a5 <= 1251; 
        o_index_for_a6 <= 1347; 
    end
    100: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 169;
        o_index_for_a1 <= 558;
        o_index_for_a2 <= 597;
        o_index_for_a3 <= 763;
        o_index_for_a4 <= 1144;
        o_index_for_a5 <= 1252; 
        o_index_for_a6 <= 1348; 
    end
    101: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 170;
        o_index_for_a1 <= 559;
        o_index_for_a2 <= 598;
        o_index_for_a3 <= 764;
        o_index_for_a4 <= 1145;
        o_index_for_a5 <= 1253; 
        o_index_for_a6 <= 1349; 
    end
    102: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 171;
        o_index_for_a1 <= 560;
        o_index_for_a2 <= 599;
        o_index_for_a3 <= 765;
        o_index_for_a4 <= 1146;
        o_index_for_a5 <= 1254; 
        o_index_for_a6 <= 1350; 
    end
    103: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 172;
        o_index_for_a1 <= 561;
        o_index_for_a2 <= 600;
        o_index_for_a3 <= 766;
        o_index_for_a4 <= 1147;
        o_index_for_a5 <= 1255; 
        o_index_for_a6 <= 1351; 
    end
    104: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 173;
        o_index_for_a1 <= 562;
        o_index_for_a2 <= 601;
        o_index_for_a3 <= 767;
        o_index_for_a4 <= 1148;
        o_index_for_a5 <= 1256; 
        o_index_for_a6 <= 1352; 
    end
    105: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 174;
        o_index_for_a1 <= 563;
        o_index_for_a2 <= 602;
        o_index_for_a3 <= 672;
        o_index_for_a4 <= 1149;
        o_index_for_a5 <= 1257; 
        o_index_for_a6 <= 1353; 
    end
    106: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 175;
        o_index_for_a1 <= 564;
        o_index_for_a2 <= 603;
        o_index_for_a3 <= 673;
        o_index_for_a4 <= 1150;
        o_index_for_a5 <= 1258; 
        o_index_for_a6 <= 1354; 
    end
    107: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 176;
        o_index_for_a1 <= 565;
        o_index_for_a2 <= 604;
        o_index_for_a3 <= 674;
        o_index_for_a4 <= 1151;
        o_index_for_a5 <= 1259; 
        o_index_for_a6 <= 1355; 
    end
    108: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 177;
        o_index_for_a1 <= 566;
        o_index_for_a2 <= 605;
        o_index_for_a3 <= 675;
        o_index_for_a4 <= 1056;
        o_index_for_a5 <= 1260; 
        o_index_for_a6 <= 1356; 
    end
    109: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 178;
        o_index_for_a1 <= 567;
        o_index_for_a2 <= 606;
        o_index_for_a3 <= 676;
        o_index_for_a4 <= 1057;
        o_index_for_a5 <= 1261; 
        o_index_for_a6 <= 1357; 
    end
    110: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 179;
        o_index_for_a1 <= 568;
        o_index_for_a2 <= 607;
        o_index_for_a3 <= 677;
        o_index_for_a4 <= 1058;
        o_index_for_a5 <= 1262; 
        o_index_for_a6 <= 1358; 
    end
    111: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 180;
        o_index_for_a1 <= 569;
        o_index_for_a2 <= 608;
        o_index_for_a3 <= 678;
        o_index_for_a4 <= 1059;
        o_index_for_a5 <= 1263; 
        o_index_for_a6 <= 1359; 
    end
    112: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 181;
        o_index_for_a1 <= 570;
        o_index_for_a2 <= 609;
        o_index_for_a3 <= 679;
        o_index_for_a4 <= 1060;
        o_index_for_a5 <= 1264; 
        o_index_for_a6 <= 1360; 
    end
    113: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 182;
        o_index_for_a1 <= 571;
        o_index_for_a2 <= 610;
        o_index_for_a3 <= 680;
        o_index_for_a4 <= 1061;
        o_index_for_a5 <= 1265; 
        o_index_for_a6 <= 1361; 
    end
    114: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 183;
        o_index_for_a1 <= 572;
        o_index_for_a2 <= 611;
        o_index_for_a3 <= 681;
        o_index_for_a4 <= 1062;
        o_index_for_a5 <= 1266; 
        o_index_for_a6 <= 1362; 
    end
    115: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 184;
        o_index_for_a1 <= 573;
        o_index_for_a2 <= 612;
        o_index_for_a3 <= 682;
        o_index_for_a4 <= 1063;
        o_index_for_a5 <= 1267; 
        o_index_for_a6 <= 1363; 
    end
    116: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 185;
        o_index_for_a1 <= 574;
        o_index_for_a2 <= 613;
        o_index_for_a3 <= 683;
        o_index_for_a4 <= 1064;
        o_index_for_a5 <= 1268; 
        o_index_for_a6 <= 1364; 
    end
    117: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 186;
        o_index_for_a1 <= 575;
        o_index_for_a2 <= 614;
        o_index_for_a3 <= 684;
        o_index_for_a4 <= 1065;
        o_index_for_a5 <= 1269; 
        o_index_for_a6 <= 1365; 
    end
    118: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 187;
        o_index_for_a1 <= 480;
        o_index_for_a2 <= 615;
        o_index_for_a3 <= 685;
        o_index_for_a4 <= 1066;
        o_index_for_a5 <= 1270; 
        o_index_for_a6 <= 1366; 
    end
    119: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 188;
        o_index_for_a1 <= 481;
        o_index_for_a2 <= 616;
        o_index_for_a3 <= 686;
        o_index_for_a4 <= 1067;
        o_index_for_a5 <= 1271; 
        o_index_for_a6 <= 1367; 
    end
    120: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 189;
        o_index_for_a1 <= 482;
        o_index_for_a2 <= 617;
        o_index_for_a3 <= 687;
        o_index_for_a4 <= 1068;
        o_index_for_a5 <= 1272; 
        o_index_for_a6 <= 1368; 
    end
    121: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 190;
        o_index_for_a1 <= 483;
        o_index_for_a2 <= 618;
        o_index_for_a3 <= 688;
        o_index_for_a4 <= 1069;
        o_index_for_a5 <= 1273; 
        o_index_for_a6 <= 1369; 
    end
    122: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 191;
        o_index_for_a1 <= 484;
        o_index_for_a2 <= 619;
        o_index_for_a3 <= 689;
        o_index_for_a4 <= 1070;
        o_index_for_a5 <= 1274; 
        o_index_for_a6 <= 1370; 
    end
    123: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 96;
        o_index_for_a1 <= 485;
        o_index_for_a2 <= 620;
        o_index_for_a3 <= 690;
        o_index_for_a4 <= 1071;
        o_index_for_a5 <= 1275; 
        o_index_for_a6 <= 1371; 
    end
    124: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 97;
        o_index_for_a1 <= 486;
        o_index_for_a2 <= 621;
        o_index_for_a3 <= 691;
        o_index_for_a4 <= 1072;
        o_index_for_a5 <= 1276; 
        o_index_for_a6 <= 1372; 
    end
    125: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 98;
        o_index_for_a1 <= 487;
        o_index_for_a2 <= 622;
        o_index_for_a3 <= 692;
        o_index_for_a4 <= 1073;
        o_index_for_a5 <= 1277; 
        o_index_for_a6 <= 1373; 
    end
    126: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 99;
        o_index_for_a1 <= 488;
        o_index_for_a2 <= 623;
        o_index_for_a3 <= 693;
        o_index_for_a4 <= 1074;
        o_index_for_a5 <= 1278; 
        o_index_for_a6 <= 1374; 
    end
    127: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 100;
        o_index_for_a1 <= 489;
        o_index_for_a2 <= 624;
        o_index_for_a3 <= 694;
        o_index_for_a4 <= 1075;
        o_index_for_a5 <= 1279; 
        o_index_for_a6 <= 1375; 
    end
    128: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 101;
        o_index_for_a1 <= 490;
        o_index_for_a2 <= 625;
        o_index_for_a3 <= 695;
        o_index_for_a4 <= 1076;
        o_index_for_a5 <= 1280; 
        o_index_for_a6 <= 1376; 
    end
    129: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 102;
        o_index_for_a1 <= 491;
        o_index_for_a2 <= 626;
        o_index_for_a3 <= 696;
        o_index_for_a4 <= 1077;
        o_index_for_a5 <= 1281; 
        o_index_for_a6 <= 1377; 
    end
    130: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 103;
        o_index_for_a1 <= 492;
        o_index_for_a2 <= 627;
        o_index_for_a3 <= 697;
        o_index_for_a4 <= 1078;
        o_index_for_a5 <= 1282; 
        o_index_for_a6 <= 1378; 
    end
    131: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 104;
        o_index_for_a1 <= 493;
        o_index_for_a2 <= 628;
        o_index_for_a3 <= 698;
        o_index_for_a4 <= 1079;
        o_index_for_a5 <= 1283; 
        o_index_for_a6 <= 1379; 
    end
    132: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 105;
        o_index_for_a1 <= 494;
        o_index_for_a2 <= 629;
        o_index_for_a3 <= 699;
        o_index_for_a4 <= 1080;
        o_index_for_a5 <= 1284; 
        o_index_for_a6 <= 1380; 
    end
    133: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 106;
        o_index_for_a1 <= 495;
        o_index_for_a2 <= 630;
        o_index_for_a3 <= 700;
        o_index_for_a4 <= 1081;
        o_index_for_a5 <= 1285; 
        o_index_for_a6 <= 1381; 
    end
    134: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 107;
        o_index_for_a1 <= 496;
        o_index_for_a2 <= 631;
        o_index_for_a3 <= 701;
        o_index_for_a4 <= 1082;
        o_index_for_a5 <= 1286; 
        o_index_for_a6 <= 1382; 
    end
    135: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 108;
        o_index_for_a1 <= 497;
        o_index_for_a2 <= 632;
        o_index_for_a3 <= 702;
        o_index_for_a4 <= 1083;
        o_index_for_a5 <= 1287; 
        o_index_for_a6 <= 1383; 
    end
    136: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 109;
        o_index_for_a1 <= 498;
        o_index_for_a2 <= 633;
        o_index_for_a3 <= 703;
        o_index_for_a4 <= 1084;
        o_index_for_a5 <= 1288; 
        o_index_for_a6 <= 1384; 
    end
    137: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 110;
        o_index_for_a1 <= 499;
        o_index_for_a2 <= 634;
        o_index_for_a3 <= 704;
        o_index_for_a4 <= 1085;
        o_index_for_a5 <= 1289; 
        o_index_for_a6 <= 1385; 
    end
    138: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 111;
        o_index_for_a1 <= 500;
        o_index_for_a2 <= 635;
        o_index_for_a3 <= 705;
        o_index_for_a4 <= 1086;
        o_index_for_a5 <= 1290; 
        o_index_for_a6 <= 1386; 
    end
    139: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 112;
        o_index_for_a1 <= 501;
        o_index_for_a2 <= 636;
        o_index_for_a3 <= 706;
        o_index_for_a4 <= 1087;
        o_index_for_a5 <= 1291; 
        o_index_for_a6 <= 1387; 
    end
    140: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 113;
        o_index_for_a1 <= 502;
        o_index_for_a2 <= 637;
        o_index_for_a3 <= 707;
        o_index_for_a4 <= 1088;
        o_index_for_a5 <= 1292; 
        o_index_for_a6 <= 1388; 
    end
    141: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 114;
        o_index_for_a1 <= 503;
        o_index_for_a2 <= 638;
        o_index_for_a3 <= 708;
        o_index_for_a4 <= 1089;
        o_index_for_a5 <= 1293; 
        o_index_for_a6 <= 1389; 
    end
    142: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 115;
        o_index_for_a1 <= 504;
        o_index_for_a2 <= 639;
        o_index_for_a3 <= 709;
        o_index_for_a4 <= 1090;
        o_index_for_a5 <= 1294; 
        o_index_for_a6 <= 1390; 
    end
    143: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 116;
        o_index_for_a1 <= 505;
        o_index_for_a2 <= 640;
        o_index_for_a3 <= 710;
        o_index_for_a4 <= 1091;
        o_index_for_a5 <= 1295; 
        o_index_for_a6 <= 1391; 
    end
    144: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 117;
        o_index_for_a1 <= 506;
        o_index_for_a2 <= 641;
        o_index_for_a3 <= 711;
        o_index_for_a4 <= 1092;
        o_index_for_a5 <= 1296; 
        o_index_for_a6 <= 1392; 
    end
    145: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 118;
        o_index_for_a1 <= 507;
        o_index_for_a2 <= 642;
        o_index_for_a3 <= 712;
        o_index_for_a4 <= 1093;
        o_index_for_a5 <= 1297; 
        o_index_for_a6 <= 1393; 
    end
    146: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 119;
        o_index_for_a1 <= 508;
        o_index_for_a2 <= 643;
        o_index_for_a3 <= 713;
        o_index_for_a4 <= 1094;
        o_index_for_a5 <= 1298; 
        o_index_for_a6 <= 1394; 
    end
    147: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 120;
        o_index_for_a1 <= 509;
        o_index_for_a2 <= 644;
        o_index_for_a3 <= 714;
        o_index_for_a4 <= 1095;
        o_index_for_a5 <= 1299; 
        o_index_for_a6 <= 1395; 
    end
    148: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 121;
        o_index_for_a1 <= 510;
        o_index_for_a2 <= 645;
        o_index_for_a3 <= 715;
        o_index_for_a4 <= 1096;
        o_index_for_a5 <= 1300; 
        o_index_for_a6 <= 1396; 
    end
    149: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 122;
        o_index_for_a1 <= 511;
        o_index_for_a2 <= 646;
        o_index_for_a3 <= 716;
        o_index_for_a4 <= 1097;
        o_index_for_a5 <= 1301; 
        o_index_for_a6 <= 1397; 
    end
    150: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 123;
        o_index_for_a1 <= 512;
        o_index_for_a2 <= 647;
        o_index_for_a3 <= 717;
        o_index_for_a4 <= 1098;
        o_index_for_a5 <= 1302; 
        o_index_for_a6 <= 1398; 
    end
    151: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 124;
        o_index_for_a1 <= 513;
        o_index_for_a2 <= 648;
        o_index_for_a3 <= 718;
        o_index_for_a4 <= 1099;
        o_index_for_a5 <= 1303; 
        o_index_for_a6 <= 1399; 
    end
    152: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 125;
        o_index_for_a1 <= 514;
        o_index_for_a2 <= 649;
        o_index_for_a3 <= 719;
        o_index_for_a4 <= 1100;
        o_index_for_a5 <= 1304; 
        o_index_for_a6 <= 1400; 
    end
    153: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 126;
        o_index_for_a1 <= 515;
        o_index_for_a2 <= 650;
        o_index_for_a3 <= 720;
        o_index_for_a4 <= 1101;
        o_index_for_a5 <= 1305; 
        o_index_for_a6 <= 1401; 
    end
    154: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 127;
        o_index_for_a1 <= 516;
        o_index_for_a2 <= 651;
        o_index_for_a3 <= 721;
        o_index_for_a4 <= 1102;
        o_index_for_a5 <= 1306; 
        o_index_for_a6 <= 1402; 
    end
    155: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 128;
        o_index_for_a1 <= 517;
        o_index_for_a2 <= 652;
        o_index_for_a3 <= 722;
        o_index_for_a4 <= 1103;
        o_index_for_a5 <= 1307; 
        o_index_for_a6 <= 1403; 
    end
    156: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 129;
        o_index_for_a1 <= 518;
        o_index_for_a2 <= 653;
        o_index_for_a3 <= 723;
        o_index_for_a4 <= 1104;
        o_index_for_a5 <= 1308; 
        o_index_for_a6 <= 1404; 
    end
    157: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 130;
        o_index_for_a1 <= 519;
        o_index_for_a2 <= 654;
        o_index_for_a3 <= 724;
        o_index_for_a4 <= 1105;
        o_index_for_a5 <= 1309; 
        o_index_for_a6 <= 1405; 
    end
    158: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 131;
        o_index_for_a1 <= 520;
        o_index_for_a2 <= 655;
        o_index_for_a3 <= 725;
        o_index_for_a4 <= 1106;
        o_index_for_a5 <= 1310; 
        o_index_for_a6 <= 1406; 
    end
    159: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 132;
        o_index_for_a1 <= 521;
        o_index_for_a2 <= 656;
        o_index_for_a3 <= 726;
        o_index_for_a4 <= 1107;
        o_index_for_a5 <= 1311; 
        o_index_for_a6 <= 1407; 
    end
    160: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 133;
        o_index_for_a1 <= 522;
        o_index_for_a2 <= 657;
        o_index_for_a3 <= 727;
        o_index_for_a4 <= 1108;
        o_index_for_a5 <= 1312; 
        o_index_for_a6 <= 1408; 
    end
    161: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 134;
        o_index_for_a1 <= 523;
        o_index_for_a2 <= 658;
        o_index_for_a3 <= 728;
        o_index_for_a4 <= 1109;
        o_index_for_a5 <= 1313; 
        o_index_for_a6 <= 1409; 
    end
    162: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 135;
        o_index_for_a1 <= 524;
        o_index_for_a2 <= 659;
        o_index_for_a3 <= 729;
        o_index_for_a4 <= 1110;
        o_index_for_a5 <= 1314; 
        o_index_for_a6 <= 1410; 
    end
    163: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 136;
        o_index_for_a1 <= 525;
        o_index_for_a2 <= 660;
        o_index_for_a3 <= 730;
        o_index_for_a4 <= 1111;
        o_index_for_a5 <= 1315; 
        o_index_for_a6 <= 1411; 
    end
    164: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 137;
        o_index_for_a1 <= 526;
        o_index_for_a2 <= 661;
        o_index_for_a3 <= 731;
        o_index_for_a4 <= 1112;
        o_index_for_a5 <= 1316; 
        o_index_for_a6 <= 1412; 
    end
    165: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 138;
        o_index_for_a1 <= 527;
        o_index_for_a2 <= 662;
        o_index_for_a3 <= 732;
        o_index_for_a4 <= 1113;
        o_index_for_a5 <= 1317; 
        o_index_for_a6 <= 1413; 
    end
    166: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 139;
        o_index_for_a1 <= 528;
        o_index_for_a2 <= 663;
        o_index_for_a3 <= 733;
        o_index_for_a4 <= 1114;
        o_index_for_a5 <= 1318; 
        o_index_for_a6 <= 1414; 
    end
    167: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 140;
        o_index_for_a1 <= 529;
        o_index_for_a2 <= 664;
        o_index_for_a3 <= 734;
        o_index_for_a4 <= 1115;
        o_index_for_a5 <= 1319; 
        o_index_for_a6 <= 1415; 
    end
    168: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 141;
        o_index_for_a1 <= 530;
        o_index_for_a2 <= 665;
        o_index_for_a3 <= 735;
        o_index_for_a4 <= 1116;
        o_index_for_a5 <= 1320; 
        o_index_for_a6 <= 1416; 
    end
    169: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 142;
        o_index_for_a1 <= 531;
        o_index_for_a2 <= 666;
        o_index_for_a3 <= 736;
        o_index_for_a4 <= 1117;
        o_index_for_a5 <= 1321; 
        o_index_for_a6 <= 1417; 
    end
    170: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 143;
        o_index_for_a1 <= 532;
        o_index_for_a2 <= 667;
        o_index_for_a3 <= 737;
        o_index_for_a4 <= 1118;
        o_index_for_a5 <= 1322; 
        o_index_for_a6 <= 1418; 
    end
    171: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 144;
        o_index_for_a1 <= 533;
        o_index_for_a2 <= 668;
        o_index_for_a3 <= 738;
        o_index_for_a4 <= 1119;
        o_index_for_a5 <= 1323; 
        o_index_for_a6 <= 1419; 
    end
    172: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 145;
        o_index_for_a1 <= 534;
        o_index_for_a2 <= 669;
        o_index_for_a3 <= 739;
        o_index_for_a4 <= 1120;
        o_index_for_a5 <= 1324; 
        o_index_for_a6 <= 1420; 
    end
    173: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 146;
        o_index_for_a1 <= 535;
        o_index_for_a2 <= 670;
        o_index_for_a3 <= 740;
        o_index_for_a4 <= 1121;
        o_index_for_a5 <= 1325; 
        o_index_for_a6 <= 1421; 
    end
    174: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 147;
        o_index_for_a1 <= 536;
        o_index_for_a2 <= 671;
        o_index_for_a3 <= 741;
        o_index_for_a4 <= 1122;
        o_index_for_a5 <= 1326; 
        o_index_for_a6 <= 1422; 
    end
    175: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 148;
        o_index_for_a1 <= 537;
        o_index_for_a2 <= 576;
        o_index_for_a3 <= 742;
        o_index_for_a4 <= 1123;
        o_index_for_a5 <= 1327; 
        o_index_for_a6 <= 1423; 
    end
    176: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 149;
        o_index_for_a1 <= 538;
        o_index_for_a2 <= 577;
        o_index_for_a3 <= 743;
        o_index_for_a4 <= 1124;
        o_index_for_a5 <= 1328; 
        o_index_for_a6 <= 1424; 
    end
    177: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 150;
        o_index_for_a1 <= 539;
        o_index_for_a2 <= 578;
        o_index_for_a3 <= 744;
        o_index_for_a4 <= 1125;
        o_index_for_a5 <= 1329; 
        o_index_for_a6 <= 1425; 
    end
    178: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 151;
        o_index_for_a1 <= 540;
        o_index_for_a2 <= 579;
        o_index_for_a3 <= 745;
        o_index_for_a4 <= 1126;
        o_index_for_a5 <= 1330; 
        o_index_for_a6 <= 1426; 
    end
    179: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 152;
        o_index_for_a1 <= 541;
        o_index_for_a2 <= 580;
        o_index_for_a3 <= 746;
        o_index_for_a4 <= 1127;
        o_index_for_a5 <= 1331; 
        o_index_for_a6 <= 1427; 
    end
    180: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 153;
        o_index_for_a1 <= 542;
        o_index_for_a2 <= 581;
        o_index_for_a3 <= 747;
        o_index_for_a4 <= 1128;
        o_index_for_a5 <= 1332; 
        o_index_for_a6 <= 1428; 
    end
    181: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 154;
        o_index_for_a1 <= 543;
        o_index_for_a2 <= 582;
        o_index_for_a3 <= 748;
        o_index_for_a4 <= 1129;
        o_index_for_a5 <= 1333; 
        o_index_for_a6 <= 1429; 
    end
    182: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 155;
        o_index_for_a1 <= 544;
        o_index_for_a2 <= 583;
        o_index_for_a3 <= 749;
        o_index_for_a4 <= 1130;
        o_index_for_a5 <= 1334; 
        o_index_for_a6 <= 1430; 
    end
    183: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 156;
        o_index_for_a1 <= 545;
        o_index_for_a2 <= 584;
        o_index_for_a3 <= 750;
        o_index_for_a4 <= 1131;
        o_index_for_a5 <= 1335; 
        o_index_for_a6 <= 1431; 
    end
    184: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 157;
        o_index_for_a1 <= 546;
        o_index_for_a2 <= 585;
        o_index_for_a3 <= 751;
        o_index_for_a4 <= 1132;
        o_index_for_a5 <= 1336; 
        o_index_for_a6 <= 1432; 
    end
    185: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 158;
        o_index_for_a1 <= 547;
        o_index_for_a2 <= 586;
        o_index_for_a3 <= 752;
        o_index_for_a4 <= 1133;
        o_index_for_a5 <= 1337; 
        o_index_for_a6 <= 1433; 
    end
    186: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 159;
        o_index_for_a1 <= 548;
        o_index_for_a2 <= 587;
        o_index_for_a3 <= 753;
        o_index_for_a4 <= 1134;
        o_index_for_a5 <= 1338; 
        o_index_for_a6 <= 1434; 
    end
    187: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 160;
        o_index_for_a1 <= 549;
        o_index_for_a2 <= 588;
        o_index_for_a3 <= 754;
        o_index_for_a4 <= 1135;
        o_index_for_a5 <= 1339; 
        o_index_for_a6 <= 1435; 
    end
    188: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 161;
        o_index_for_a1 <= 550;
        o_index_for_a2 <= 589;
        o_index_for_a3 <= 755;
        o_index_for_a4 <= 1136;
        o_index_for_a5 <= 1340; 
        o_index_for_a6 <= 1436; 
    end
    189: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 162;
        o_index_for_a1 <= 551;
        o_index_for_a2 <= 590;
        o_index_for_a3 <= 756;
        o_index_for_a4 <= 1137;
        o_index_for_a5 <= 1341; 
        o_index_for_a6 <= 1437; 
    end
    190: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 163;
        o_index_for_a1 <= 552;
        o_index_for_a2 <= 591;
        o_index_for_a3 <= 757;
        o_index_for_a4 <= 1138;
        o_index_for_a5 <= 1342; 
        o_index_for_a6 <= 1438; 
    end
    191: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 0;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 0;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 164;
        o_index_for_a1 <= 553;
        o_index_for_a2 <= 592;
        o_index_for_a3 <= 758;
        o_index_for_a4 <= 1139;
        o_index_for_a5 <= 1343; 
        o_index_for_a6 <= 1439; 
    end
    192: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 360;
        o_index_for_a1 <= 458;
        o_index_for_a2 <= 495;
        o_index_for_a3 <= 735;
        o_index_for_a4 <= 1056;
        o_index_for_a5 <= 1344; 
        o_index_for_a6 <= 1440; 
    end
    193: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 361;
        o_index_for_a1 <= 459;
        o_index_for_a2 <= 496;
        o_index_for_a3 <= 736;
        o_index_for_a4 <= 1057;
        o_index_for_a5 <= 1345; 
        o_index_for_a6 <= 1441; 
    end
    194: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 362;
        o_index_for_a1 <= 460;
        o_index_for_a2 <= 497;
        o_index_for_a3 <= 737;
        o_index_for_a4 <= 1058;
        o_index_for_a5 <= 1346; 
        o_index_for_a6 <= 1442; 
    end
    195: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 363;
        o_index_for_a1 <= 461;
        o_index_for_a2 <= 498;
        o_index_for_a3 <= 738;
        o_index_for_a4 <= 1059;
        o_index_for_a5 <= 1347; 
        o_index_for_a6 <= 1443; 
    end
    196: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 364;
        o_index_for_a1 <= 462;
        o_index_for_a2 <= 499;
        o_index_for_a3 <= 739;
        o_index_for_a4 <= 1060;
        o_index_for_a5 <= 1348; 
        o_index_for_a6 <= 1444; 
    end
    197: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 365;
        o_index_for_a1 <= 463;
        o_index_for_a2 <= 500;
        o_index_for_a3 <= 740;
        o_index_for_a4 <= 1061;
        o_index_for_a5 <= 1349; 
        o_index_for_a6 <= 1445; 
    end
    198: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 366;
        o_index_for_a1 <= 464;
        o_index_for_a2 <= 501;
        o_index_for_a3 <= 741;
        o_index_for_a4 <= 1062;
        o_index_for_a5 <= 1350; 
        o_index_for_a6 <= 1446; 
    end
    199: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 367;
        o_index_for_a1 <= 465;
        o_index_for_a2 <= 502;
        o_index_for_a3 <= 742;
        o_index_for_a4 <= 1063;
        o_index_for_a5 <= 1351; 
        o_index_for_a6 <= 1447; 
    end
    200: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 368;
        o_index_for_a1 <= 466;
        o_index_for_a2 <= 503;
        o_index_for_a3 <= 743;
        o_index_for_a4 <= 1064;
        o_index_for_a5 <= 1352; 
        o_index_for_a6 <= 1448; 
    end
    201: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 369;
        o_index_for_a1 <= 467;
        o_index_for_a2 <= 504;
        o_index_for_a3 <= 744;
        o_index_for_a4 <= 1065;
        o_index_for_a5 <= 1353; 
        o_index_for_a6 <= 1449; 
    end
    202: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 370;
        o_index_for_a1 <= 468;
        o_index_for_a2 <= 505;
        o_index_for_a3 <= 745;
        o_index_for_a4 <= 1066;
        o_index_for_a5 <= 1354; 
        o_index_for_a6 <= 1450; 
    end
    203: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 371;
        o_index_for_a1 <= 469;
        o_index_for_a2 <= 506;
        o_index_for_a3 <= 746;
        o_index_for_a4 <= 1067;
        o_index_for_a5 <= 1355; 
        o_index_for_a6 <= 1451; 
    end
    204: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 372;
        o_index_for_a1 <= 470;
        o_index_for_a2 <= 507;
        o_index_for_a3 <= 747;
        o_index_for_a4 <= 1068;
        o_index_for_a5 <= 1356; 
        o_index_for_a6 <= 1452; 
    end
    205: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 373;
        o_index_for_a1 <= 471;
        o_index_for_a2 <= 508;
        o_index_for_a3 <= 748;
        o_index_for_a4 <= 1069;
        o_index_for_a5 <= 1357; 
        o_index_for_a6 <= 1453; 
    end
    206: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 374;
        o_index_for_a1 <= 472;
        o_index_for_a2 <= 509;
        o_index_for_a3 <= 749;
        o_index_for_a4 <= 1070;
        o_index_for_a5 <= 1358; 
        o_index_for_a6 <= 1454; 
    end
    207: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 375;
        o_index_for_a1 <= 473;
        o_index_for_a2 <= 510;
        o_index_for_a3 <= 750;
        o_index_for_a4 <= 1071;
        o_index_for_a5 <= 1359; 
        o_index_for_a6 <= 1455; 
    end
    208: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 376;
        o_index_for_a1 <= 474;
        o_index_for_a2 <= 511;
        o_index_for_a3 <= 751;
        o_index_for_a4 <= 1072;
        o_index_for_a5 <= 1360; 
        o_index_for_a6 <= 1456; 
    end
    209: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 377;
        o_index_for_a1 <= 475;
        o_index_for_a2 <= 512;
        o_index_for_a3 <= 752;
        o_index_for_a4 <= 1073;
        o_index_for_a5 <= 1361; 
        o_index_for_a6 <= 1457; 
    end
    210: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 378;
        o_index_for_a1 <= 476;
        o_index_for_a2 <= 513;
        o_index_for_a3 <= 753;
        o_index_for_a4 <= 1074;
        o_index_for_a5 <= 1362; 
        o_index_for_a6 <= 1458; 
    end
    211: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 379;
        o_index_for_a1 <= 477;
        o_index_for_a2 <= 514;
        o_index_for_a3 <= 754;
        o_index_for_a4 <= 1075;
        o_index_for_a5 <= 1363; 
        o_index_for_a6 <= 1459; 
    end
    212: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 380;
        o_index_for_a1 <= 478;
        o_index_for_a2 <= 515;
        o_index_for_a3 <= 755;
        o_index_for_a4 <= 1076;
        o_index_for_a5 <= 1364; 
        o_index_for_a6 <= 1460; 
    end
    213: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 381;
        o_index_for_a1 <= 479;
        o_index_for_a2 <= 516;
        o_index_for_a3 <= 756;
        o_index_for_a4 <= 1077;
        o_index_for_a5 <= 1365; 
        o_index_for_a6 <= 1461; 
    end
    214: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 382;
        o_index_for_a1 <= 384;
        o_index_for_a2 <= 517;
        o_index_for_a3 <= 757;
        o_index_for_a4 <= 1078;
        o_index_for_a5 <= 1366; 
        o_index_for_a6 <= 1462; 
    end
    215: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 383;
        o_index_for_a1 <= 385;
        o_index_for_a2 <= 518;
        o_index_for_a3 <= 758;
        o_index_for_a4 <= 1079;
        o_index_for_a5 <= 1367; 
        o_index_for_a6 <= 1463; 
    end
    216: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 288;
        o_index_for_a1 <= 386;
        o_index_for_a2 <= 519;
        o_index_for_a3 <= 759;
        o_index_for_a4 <= 1080;
        o_index_for_a5 <= 1368; 
        o_index_for_a6 <= 1464; 
    end
    217: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 289;
        o_index_for_a1 <= 387;
        o_index_for_a2 <= 520;
        o_index_for_a3 <= 760;
        o_index_for_a4 <= 1081;
        o_index_for_a5 <= 1369; 
        o_index_for_a6 <= 1465; 
    end
    218: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 290;
        o_index_for_a1 <= 388;
        o_index_for_a2 <= 521;
        o_index_for_a3 <= 761;
        o_index_for_a4 <= 1082;
        o_index_for_a5 <= 1370; 
        o_index_for_a6 <= 1466; 
    end
    219: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 291;
        o_index_for_a1 <= 389;
        o_index_for_a2 <= 522;
        o_index_for_a3 <= 762;
        o_index_for_a4 <= 1083;
        o_index_for_a5 <= 1371; 
        o_index_for_a6 <= 1467; 
    end
    220: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 292;
        o_index_for_a1 <= 390;
        o_index_for_a2 <= 523;
        o_index_for_a3 <= 763;
        o_index_for_a4 <= 1084;
        o_index_for_a5 <= 1372; 
        o_index_for_a6 <= 1468; 
    end
    221: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 293;
        o_index_for_a1 <= 391;
        o_index_for_a2 <= 524;
        o_index_for_a3 <= 764;
        o_index_for_a4 <= 1085;
        o_index_for_a5 <= 1373; 
        o_index_for_a6 <= 1469; 
    end
    222: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 294;
        o_index_for_a1 <= 392;
        o_index_for_a2 <= 525;
        o_index_for_a3 <= 765;
        o_index_for_a4 <= 1086;
        o_index_for_a5 <= 1374; 
        o_index_for_a6 <= 1470; 
    end
    223: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 295;
        o_index_for_a1 <= 393;
        o_index_for_a2 <= 526;
        o_index_for_a3 <= 766;
        o_index_for_a4 <= 1087;
        o_index_for_a5 <= 1375; 
        o_index_for_a6 <= 1471; 
    end
    224: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 296;
        o_index_for_a1 <= 394;
        o_index_for_a2 <= 527;
        o_index_for_a3 <= 767;
        o_index_for_a4 <= 1088;
        o_index_for_a5 <= 1376; 
        o_index_for_a6 <= 1472; 
    end
    225: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 297;
        o_index_for_a1 <= 395;
        o_index_for_a2 <= 528;
        o_index_for_a3 <= 672;
        o_index_for_a4 <= 1089;
        o_index_for_a5 <= 1377; 
        o_index_for_a6 <= 1473; 
    end
    226: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 298;
        o_index_for_a1 <= 396;
        o_index_for_a2 <= 529;
        o_index_for_a3 <= 673;
        o_index_for_a4 <= 1090;
        o_index_for_a5 <= 1378; 
        o_index_for_a6 <= 1474; 
    end
    227: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 299;
        o_index_for_a1 <= 397;
        o_index_for_a2 <= 530;
        o_index_for_a3 <= 674;
        o_index_for_a4 <= 1091;
        o_index_for_a5 <= 1379; 
        o_index_for_a6 <= 1475; 
    end
    228: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 300;
        o_index_for_a1 <= 398;
        o_index_for_a2 <= 531;
        o_index_for_a3 <= 675;
        o_index_for_a4 <= 1092;
        o_index_for_a5 <= 1380; 
        o_index_for_a6 <= 1476; 
    end
    229: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 301;
        o_index_for_a1 <= 399;
        o_index_for_a2 <= 532;
        o_index_for_a3 <= 676;
        o_index_for_a4 <= 1093;
        o_index_for_a5 <= 1381; 
        o_index_for_a6 <= 1477; 
    end
    230: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 302;
        o_index_for_a1 <= 400;
        o_index_for_a2 <= 533;
        o_index_for_a3 <= 677;
        o_index_for_a4 <= 1094;
        o_index_for_a5 <= 1382; 
        o_index_for_a6 <= 1478; 
    end
    231: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 303;
        o_index_for_a1 <= 401;
        o_index_for_a2 <= 534;
        o_index_for_a3 <= 678;
        o_index_for_a4 <= 1095;
        o_index_for_a5 <= 1383; 
        o_index_for_a6 <= 1479; 
    end
    232: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 304;
        o_index_for_a1 <= 402;
        o_index_for_a2 <= 535;
        o_index_for_a3 <= 679;
        o_index_for_a4 <= 1096;
        o_index_for_a5 <= 1384; 
        o_index_for_a6 <= 1480; 
    end
    233: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 305;
        o_index_for_a1 <= 403;
        o_index_for_a2 <= 536;
        o_index_for_a3 <= 680;
        o_index_for_a4 <= 1097;
        o_index_for_a5 <= 1385; 
        o_index_for_a6 <= 1481; 
    end
    234: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 306;
        o_index_for_a1 <= 404;
        o_index_for_a2 <= 537;
        o_index_for_a3 <= 681;
        o_index_for_a4 <= 1098;
        o_index_for_a5 <= 1386; 
        o_index_for_a6 <= 1482; 
    end
    235: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 307;
        o_index_for_a1 <= 405;
        o_index_for_a2 <= 538;
        o_index_for_a3 <= 682;
        o_index_for_a4 <= 1099;
        o_index_for_a5 <= 1387; 
        o_index_for_a6 <= 1483; 
    end
    236: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 308;
        o_index_for_a1 <= 406;
        o_index_for_a2 <= 539;
        o_index_for_a3 <= 683;
        o_index_for_a4 <= 1100;
        o_index_for_a5 <= 1388; 
        o_index_for_a6 <= 1484; 
    end
    237: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 309;
        o_index_for_a1 <= 407;
        o_index_for_a2 <= 540;
        o_index_for_a3 <= 684;
        o_index_for_a4 <= 1101;
        o_index_for_a5 <= 1389; 
        o_index_for_a6 <= 1485; 
    end
    238: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 310;
        o_index_for_a1 <= 408;
        o_index_for_a2 <= 541;
        o_index_for_a3 <= 685;
        o_index_for_a4 <= 1102;
        o_index_for_a5 <= 1390; 
        o_index_for_a6 <= 1486; 
    end
    239: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 311;
        o_index_for_a1 <= 409;
        o_index_for_a2 <= 542;
        o_index_for_a3 <= 686;
        o_index_for_a4 <= 1103;
        o_index_for_a5 <= 1391; 
        o_index_for_a6 <= 1487; 
    end
    240: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 312;
        o_index_for_a1 <= 410;
        o_index_for_a2 <= 543;
        o_index_for_a3 <= 687;
        o_index_for_a4 <= 1104;
        o_index_for_a5 <= 1392; 
        o_index_for_a6 <= 1488; 
    end
    241: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 313;
        o_index_for_a1 <= 411;
        o_index_for_a2 <= 544;
        o_index_for_a3 <= 688;
        o_index_for_a4 <= 1105;
        o_index_for_a5 <= 1393; 
        o_index_for_a6 <= 1489; 
    end
    242: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 314;
        o_index_for_a1 <= 412;
        o_index_for_a2 <= 545;
        o_index_for_a3 <= 689;
        o_index_for_a4 <= 1106;
        o_index_for_a5 <= 1394; 
        o_index_for_a6 <= 1490; 
    end
    243: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 315;
        o_index_for_a1 <= 413;
        o_index_for_a2 <= 546;
        o_index_for_a3 <= 690;
        o_index_for_a4 <= 1107;
        o_index_for_a5 <= 1395; 
        o_index_for_a6 <= 1491; 
    end
    244: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 316;
        o_index_for_a1 <= 414;
        o_index_for_a2 <= 547;
        o_index_for_a3 <= 691;
        o_index_for_a4 <= 1108;
        o_index_for_a5 <= 1396; 
        o_index_for_a6 <= 1492; 
    end
    245: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 317;
        o_index_for_a1 <= 415;
        o_index_for_a2 <= 548;
        o_index_for_a3 <= 692;
        o_index_for_a4 <= 1109;
        o_index_for_a5 <= 1397; 
        o_index_for_a6 <= 1493; 
    end
    246: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 318;
        o_index_for_a1 <= 416;
        o_index_for_a2 <= 549;
        o_index_for_a3 <= 693;
        o_index_for_a4 <= 1110;
        o_index_for_a5 <= 1398; 
        o_index_for_a6 <= 1494; 
    end
    247: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 319;
        o_index_for_a1 <= 417;
        o_index_for_a2 <= 550;
        o_index_for_a3 <= 694;
        o_index_for_a4 <= 1111;
        o_index_for_a5 <= 1399; 
        o_index_for_a6 <= 1495; 
    end
    248: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 320;
        o_index_for_a1 <= 418;
        o_index_for_a2 <= 551;
        o_index_for_a3 <= 695;
        o_index_for_a4 <= 1112;
        o_index_for_a5 <= 1400; 
        o_index_for_a6 <= 1496; 
    end
    249: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 321;
        o_index_for_a1 <= 419;
        o_index_for_a2 <= 552;
        o_index_for_a3 <= 696;
        o_index_for_a4 <= 1113;
        o_index_for_a5 <= 1401; 
        o_index_for_a6 <= 1497; 
    end
    250: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 322;
        o_index_for_a1 <= 420;
        o_index_for_a2 <= 553;
        o_index_for_a3 <= 697;
        o_index_for_a4 <= 1114;
        o_index_for_a5 <= 1402; 
        o_index_for_a6 <= 1498; 
    end
    251: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 323;
        o_index_for_a1 <= 421;
        o_index_for_a2 <= 554;
        o_index_for_a3 <= 698;
        o_index_for_a4 <= 1115;
        o_index_for_a5 <= 1403; 
        o_index_for_a6 <= 1499; 
    end
    252: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 324;
        o_index_for_a1 <= 422;
        o_index_for_a2 <= 555;
        o_index_for_a3 <= 699;
        o_index_for_a4 <= 1116;
        o_index_for_a5 <= 1404; 
        o_index_for_a6 <= 1500; 
    end
    253: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 325;
        o_index_for_a1 <= 423;
        o_index_for_a2 <= 556;
        o_index_for_a3 <= 700;
        o_index_for_a4 <= 1117;
        o_index_for_a5 <= 1405; 
        o_index_for_a6 <= 1501; 
    end
    254: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 326;
        o_index_for_a1 <= 424;
        o_index_for_a2 <= 557;
        o_index_for_a3 <= 701;
        o_index_for_a4 <= 1118;
        o_index_for_a5 <= 1406; 
        o_index_for_a6 <= 1502; 
    end
    255: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 327;
        o_index_for_a1 <= 425;
        o_index_for_a2 <= 558;
        o_index_for_a3 <= 702;
        o_index_for_a4 <= 1119;
        o_index_for_a5 <= 1407; 
        o_index_for_a6 <= 1503; 
    end
    256: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 328;
        o_index_for_a1 <= 426;
        o_index_for_a2 <= 559;
        o_index_for_a3 <= 703;
        o_index_for_a4 <= 1120;
        o_index_for_a5 <= 1408; 
        o_index_for_a6 <= 1504; 
    end
    257: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 329;
        o_index_for_a1 <= 427;
        o_index_for_a2 <= 560;
        o_index_for_a3 <= 704;
        o_index_for_a4 <= 1121;
        o_index_for_a5 <= 1409; 
        o_index_for_a6 <= 1505; 
    end
    258: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 330;
        o_index_for_a1 <= 428;
        o_index_for_a2 <= 561;
        o_index_for_a3 <= 705;
        o_index_for_a4 <= 1122;
        o_index_for_a5 <= 1410; 
        o_index_for_a6 <= 1506; 
    end
    259: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 331;
        o_index_for_a1 <= 429;
        o_index_for_a2 <= 562;
        o_index_for_a3 <= 706;
        o_index_for_a4 <= 1123;
        o_index_for_a5 <= 1411; 
        o_index_for_a6 <= 1507; 
    end
    260: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 332;
        o_index_for_a1 <= 430;
        o_index_for_a2 <= 563;
        o_index_for_a3 <= 707;
        o_index_for_a4 <= 1124;
        o_index_for_a5 <= 1412; 
        o_index_for_a6 <= 1508; 
    end
    261: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 333;
        o_index_for_a1 <= 431;
        o_index_for_a2 <= 564;
        o_index_for_a3 <= 708;
        o_index_for_a4 <= 1125;
        o_index_for_a5 <= 1413; 
        o_index_for_a6 <= 1509; 
    end
    262: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 334;
        o_index_for_a1 <= 432;
        o_index_for_a2 <= 565;
        o_index_for_a3 <= 709;
        o_index_for_a4 <= 1126;
        o_index_for_a5 <= 1414; 
        o_index_for_a6 <= 1510; 
    end
    263: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 335;
        o_index_for_a1 <= 433;
        o_index_for_a2 <= 566;
        o_index_for_a3 <= 710;
        o_index_for_a4 <= 1127;
        o_index_for_a5 <= 1415; 
        o_index_for_a6 <= 1511; 
    end
    264: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 336;
        o_index_for_a1 <= 434;
        o_index_for_a2 <= 567;
        o_index_for_a3 <= 711;
        o_index_for_a4 <= 1128;
        o_index_for_a5 <= 1416; 
        o_index_for_a6 <= 1512; 
    end
    265: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 337;
        o_index_for_a1 <= 435;
        o_index_for_a2 <= 568;
        o_index_for_a3 <= 712;
        o_index_for_a4 <= 1129;
        o_index_for_a5 <= 1417; 
        o_index_for_a6 <= 1513; 
    end
    266: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 338;
        o_index_for_a1 <= 436;
        o_index_for_a2 <= 569;
        o_index_for_a3 <= 713;
        o_index_for_a4 <= 1130;
        o_index_for_a5 <= 1418; 
        o_index_for_a6 <= 1514; 
    end
    267: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 339;
        o_index_for_a1 <= 437;
        o_index_for_a2 <= 570;
        o_index_for_a3 <= 714;
        o_index_for_a4 <= 1131;
        o_index_for_a5 <= 1419; 
        o_index_for_a6 <= 1515; 
    end
    268: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 340;
        o_index_for_a1 <= 438;
        o_index_for_a2 <= 571;
        o_index_for_a3 <= 715;
        o_index_for_a4 <= 1132;
        o_index_for_a5 <= 1420; 
        o_index_for_a6 <= 1516; 
    end
    269: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 341;
        o_index_for_a1 <= 439;
        o_index_for_a2 <= 572;
        o_index_for_a3 <= 716;
        o_index_for_a4 <= 1133;
        o_index_for_a5 <= 1421; 
        o_index_for_a6 <= 1517; 
    end
    270: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 342;
        o_index_for_a1 <= 440;
        o_index_for_a2 <= 573;
        o_index_for_a3 <= 717;
        o_index_for_a4 <= 1134;
        o_index_for_a5 <= 1422; 
        o_index_for_a6 <= 1518; 
    end
    271: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 343;
        o_index_for_a1 <= 441;
        o_index_for_a2 <= 574;
        o_index_for_a3 <= 718;
        o_index_for_a4 <= 1135;
        o_index_for_a5 <= 1423; 
        o_index_for_a6 <= 1519; 
    end
    272: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 344;
        o_index_for_a1 <= 442;
        o_index_for_a2 <= 575;
        o_index_for_a3 <= 719;
        o_index_for_a4 <= 1136;
        o_index_for_a5 <= 1424; 
        o_index_for_a6 <= 1520; 
    end
    273: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 345;
        o_index_for_a1 <= 443;
        o_index_for_a2 <= 480;
        o_index_for_a3 <= 720;
        o_index_for_a4 <= 1137;
        o_index_for_a5 <= 1425; 
        o_index_for_a6 <= 1521; 
    end
    274: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 346;
        o_index_for_a1 <= 444;
        o_index_for_a2 <= 481;
        o_index_for_a3 <= 721;
        o_index_for_a4 <= 1138;
        o_index_for_a5 <= 1426; 
        o_index_for_a6 <= 1522; 
    end
    275: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 347;
        o_index_for_a1 <= 445;
        o_index_for_a2 <= 482;
        o_index_for_a3 <= 722;
        o_index_for_a4 <= 1139;
        o_index_for_a5 <= 1427; 
        o_index_for_a6 <= 1523; 
    end
    276: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 348;
        o_index_for_a1 <= 446;
        o_index_for_a2 <= 483;
        o_index_for_a3 <= 723;
        o_index_for_a4 <= 1140;
        o_index_for_a5 <= 1428; 
        o_index_for_a6 <= 1524; 
    end
    277: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 349;
        o_index_for_a1 <= 447;
        o_index_for_a2 <= 484;
        o_index_for_a3 <= 724;
        o_index_for_a4 <= 1141;
        o_index_for_a5 <= 1429; 
        o_index_for_a6 <= 1525; 
    end
    278: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 350;
        o_index_for_a1 <= 448;
        o_index_for_a2 <= 485;
        o_index_for_a3 <= 725;
        o_index_for_a4 <= 1142;
        o_index_for_a5 <= 1430; 
        o_index_for_a6 <= 1526; 
    end
    279: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 351;
        o_index_for_a1 <= 449;
        o_index_for_a2 <= 486;
        o_index_for_a3 <= 726;
        o_index_for_a4 <= 1143;
        o_index_for_a5 <= 1431; 
        o_index_for_a6 <= 1527; 
    end
    280: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 352;
        o_index_for_a1 <= 450;
        o_index_for_a2 <= 487;
        o_index_for_a3 <= 727;
        o_index_for_a4 <= 1144;
        o_index_for_a5 <= 1432; 
        o_index_for_a6 <= 1528; 
    end
    281: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 353;
        o_index_for_a1 <= 451;
        o_index_for_a2 <= 488;
        o_index_for_a3 <= 728;
        o_index_for_a4 <= 1145;
        o_index_for_a5 <= 1433; 
        o_index_for_a6 <= 1529; 
    end
    282: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 354;
        o_index_for_a1 <= 452;
        o_index_for_a2 <= 489;
        o_index_for_a3 <= 729;
        o_index_for_a4 <= 1146;
        o_index_for_a5 <= 1434; 
        o_index_for_a6 <= 1530; 
    end
    283: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 355;
        o_index_for_a1 <= 453;
        o_index_for_a2 <= 490;
        o_index_for_a3 <= 730;
        o_index_for_a4 <= 1147;
        o_index_for_a5 <= 1435; 
        o_index_for_a6 <= 1531; 
    end
    284: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 356;
        o_index_for_a1 <= 454;
        o_index_for_a2 <= 491;
        o_index_for_a3 <= 731;
        o_index_for_a4 <= 1148;
        o_index_for_a5 <= 1436; 
        o_index_for_a6 <= 1532; 
    end
    285: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 357;
        o_index_for_a1 <= 455;
        o_index_for_a2 <= 492;
        o_index_for_a3 <= 732;
        o_index_for_a4 <= 1149;
        o_index_for_a5 <= 1437; 
        o_index_for_a6 <= 1533; 
    end
    286: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 358;
        o_index_for_a1 <= 456;
        o_index_for_a2 <= 493;
        o_index_for_a3 <= 733;
        o_index_for_a4 <= 1150;
        o_index_for_a5 <= 1438; 
        o_index_for_a6 <= 1534; 
    end
    287: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 0;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 359;
        o_index_for_a1 <= 457;
        o_index_for_a2 <= 494;
        o_index_for_a3 <= 734;
        o_index_for_a4 <= 1151;
        o_index_for_a5 <= 1439; 
        o_index_for_a6 <= 1535; 
    end
    288: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 35;
        o_index_for_a1 <= 241;
        o_index_for_a2 <= 799;
        o_index_for_a3 <= 935;
        o_index_for_a4 <= 1440;
        o_index_for_a5 <= 1536; 
        o_index_for_a6 <= 2304; 
    end
    289: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 36;
        o_index_for_a1 <= 242;
        o_index_for_a2 <= 800;
        o_index_for_a3 <= 936;
        o_index_for_a4 <= 1441;
        o_index_for_a5 <= 1537; 
        o_index_for_a6 <= 2304; 
    end
    290: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 37;
        o_index_for_a1 <= 243;
        o_index_for_a2 <= 801;
        o_index_for_a3 <= 937;
        o_index_for_a4 <= 1442;
        o_index_for_a5 <= 1538; 
        o_index_for_a6 <= 2304; 
    end
    291: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 38;
        o_index_for_a1 <= 244;
        o_index_for_a2 <= 802;
        o_index_for_a3 <= 938;
        o_index_for_a4 <= 1443;
        o_index_for_a5 <= 1539; 
        o_index_for_a6 <= 2304; 
    end
    292: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 39;
        o_index_for_a1 <= 245;
        o_index_for_a2 <= 803;
        o_index_for_a3 <= 939;
        o_index_for_a4 <= 1444;
        o_index_for_a5 <= 1540; 
        o_index_for_a6 <= 2304; 
    end
    293: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 40;
        o_index_for_a1 <= 246;
        o_index_for_a2 <= 804;
        o_index_for_a3 <= 940;
        o_index_for_a4 <= 1445;
        o_index_for_a5 <= 1541; 
        o_index_for_a6 <= 2304; 
    end
    294: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 41;
        o_index_for_a1 <= 247;
        o_index_for_a2 <= 805;
        o_index_for_a3 <= 941;
        o_index_for_a4 <= 1446;
        o_index_for_a5 <= 1542; 
        o_index_for_a6 <= 2304; 
    end
    295: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 42;
        o_index_for_a1 <= 248;
        o_index_for_a2 <= 806;
        o_index_for_a3 <= 942;
        o_index_for_a4 <= 1447;
        o_index_for_a5 <= 1543; 
        o_index_for_a6 <= 2304; 
    end
    296: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 43;
        o_index_for_a1 <= 249;
        o_index_for_a2 <= 807;
        o_index_for_a3 <= 943;
        o_index_for_a4 <= 1448;
        o_index_for_a5 <= 1544; 
        o_index_for_a6 <= 2304; 
    end
    297: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 44;
        o_index_for_a1 <= 250;
        o_index_for_a2 <= 808;
        o_index_for_a3 <= 944;
        o_index_for_a4 <= 1449;
        o_index_for_a5 <= 1545; 
        o_index_for_a6 <= 2304; 
    end
    298: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 45;
        o_index_for_a1 <= 251;
        o_index_for_a2 <= 809;
        o_index_for_a3 <= 945;
        o_index_for_a4 <= 1450;
        o_index_for_a5 <= 1546; 
        o_index_for_a6 <= 2304; 
    end
    299: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 46;
        o_index_for_a1 <= 252;
        o_index_for_a2 <= 810;
        o_index_for_a3 <= 946;
        o_index_for_a4 <= 1451;
        o_index_for_a5 <= 1547; 
        o_index_for_a6 <= 2304; 
    end
    300: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 47;
        o_index_for_a1 <= 253;
        o_index_for_a2 <= 811;
        o_index_for_a3 <= 947;
        o_index_for_a4 <= 1452;
        o_index_for_a5 <= 1548; 
        o_index_for_a6 <= 2304; 
    end
    301: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 48;
        o_index_for_a1 <= 254;
        o_index_for_a2 <= 812;
        o_index_for_a3 <= 948;
        o_index_for_a4 <= 1453;
        o_index_for_a5 <= 1549; 
        o_index_for_a6 <= 2304; 
    end
    302: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 49;
        o_index_for_a1 <= 255;
        o_index_for_a2 <= 813;
        o_index_for_a3 <= 949;
        o_index_for_a4 <= 1454;
        o_index_for_a5 <= 1550; 
        o_index_for_a6 <= 2304; 
    end
    303: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 50;
        o_index_for_a1 <= 256;
        o_index_for_a2 <= 814;
        o_index_for_a3 <= 950;
        o_index_for_a4 <= 1455;
        o_index_for_a5 <= 1551; 
        o_index_for_a6 <= 2304; 
    end
    304: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 51;
        o_index_for_a1 <= 257;
        o_index_for_a2 <= 815;
        o_index_for_a3 <= 951;
        o_index_for_a4 <= 1456;
        o_index_for_a5 <= 1552; 
        o_index_for_a6 <= 2304; 
    end
    305: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 52;
        o_index_for_a1 <= 258;
        o_index_for_a2 <= 816;
        o_index_for_a3 <= 952;
        o_index_for_a4 <= 1457;
        o_index_for_a5 <= 1553; 
        o_index_for_a6 <= 2304; 
    end
    306: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 53;
        o_index_for_a1 <= 259;
        o_index_for_a2 <= 817;
        o_index_for_a3 <= 953;
        o_index_for_a4 <= 1458;
        o_index_for_a5 <= 1554; 
        o_index_for_a6 <= 2304; 
    end
    307: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 54;
        o_index_for_a1 <= 260;
        o_index_for_a2 <= 818;
        o_index_for_a3 <= 954;
        o_index_for_a4 <= 1459;
        o_index_for_a5 <= 1555; 
        o_index_for_a6 <= 2304; 
    end
    308: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 55;
        o_index_for_a1 <= 261;
        o_index_for_a2 <= 819;
        o_index_for_a3 <= 955;
        o_index_for_a4 <= 1460;
        o_index_for_a5 <= 1556; 
        o_index_for_a6 <= 2304; 
    end
    309: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 56;
        o_index_for_a1 <= 262;
        o_index_for_a2 <= 820;
        o_index_for_a3 <= 956;
        o_index_for_a4 <= 1461;
        o_index_for_a5 <= 1557; 
        o_index_for_a6 <= 2304; 
    end
    310: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 57;
        o_index_for_a1 <= 263;
        o_index_for_a2 <= 821;
        o_index_for_a3 <= 957;
        o_index_for_a4 <= 1462;
        o_index_for_a5 <= 1558; 
        o_index_for_a6 <= 2304; 
    end
    311: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 58;
        o_index_for_a1 <= 264;
        o_index_for_a2 <= 822;
        o_index_for_a3 <= 958;
        o_index_for_a4 <= 1463;
        o_index_for_a5 <= 1559; 
        o_index_for_a6 <= 2304; 
    end
    312: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 59;
        o_index_for_a1 <= 265;
        o_index_for_a2 <= 823;
        o_index_for_a3 <= 959;
        o_index_for_a4 <= 1464;
        o_index_for_a5 <= 1560; 
        o_index_for_a6 <= 2304; 
    end
    313: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 60;
        o_index_for_a1 <= 266;
        o_index_for_a2 <= 824;
        o_index_for_a3 <= 864;
        o_index_for_a4 <= 1465;
        o_index_for_a5 <= 1561; 
        o_index_for_a6 <= 2304; 
    end
    314: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 61;
        o_index_for_a1 <= 267;
        o_index_for_a2 <= 825;
        o_index_for_a3 <= 865;
        o_index_for_a4 <= 1466;
        o_index_for_a5 <= 1562; 
        o_index_for_a6 <= 2304; 
    end
    315: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 62;
        o_index_for_a1 <= 268;
        o_index_for_a2 <= 826;
        o_index_for_a3 <= 866;
        o_index_for_a4 <= 1467;
        o_index_for_a5 <= 1563; 
        o_index_for_a6 <= 2304; 
    end
    316: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 63;
        o_index_for_a1 <= 269;
        o_index_for_a2 <= 827;
        o_index_for_a3 <= 867;
        o_index_for_a4 <= 1468;
        o_index_for_a5 <= 1564; 
        o_index_for_a6 <= 2304; 
    end
    317: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 64;
        o_index_for_a1 <= 270;
        o_index_for_a2 <= 828;
        o_index_for_a3 <= 868;
        o_index_for_a4 <= 1469;
        o_index_for_a5 <= 1565; 
        o_index_for_a6 <= 2304; 
    end
    318: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 65;
        o_index_for_a1 <= 271;
        o_index_for_a2 <= 829;
        o_index_for_a3 <= 869;
        o_index_for_a4 <= 1470;
        o_index_for_a5 <= 1566; 
        o_index_for_a6 <= 2304; 
    end
    319: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 66;
        o_index_for_a1 <= 272;
        o_index_for_a2 <= 830;
        o_index_for_a3 <= 870;
        o_index_for_a4 <= 1471;
        o_index_for_a5 <= 1567; 
        o_index_for_a6 <= 2304; 
    end
    320: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 67;
        o_index_for_a1 <= 273;
        o_index_for_a2 <= 831;
        o_index_for_a3 <= 871;
        o_index_for_a4 <= 1472;
        o_index_for_a5 <= 1568; 
        o_index_for_a6 <= 2304; 
    end
    321: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 68;
        o_index_for_a1 <= 274;
        o_index_for_a2 <= 832;
        o_index_for_a3 <= 872;
        o_index_for_a4 <= 1473;
        o_index_for_a5 <= 1569; 
        o_index_for_a6 <= 2304; 
    end
    322: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 69;
        o_index_for_a1 <= 275;
        o_index_for_a2 <= 833;
        o_index_for_a3 <= 873;
        o_index_for_a4 <= 1474;
        o_index_for_a5 <= 1570; 
        o_index_for_a6 <= 2304; 
    end
    323: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 70;
        o_index_for_a1 <= 276;
        o_index_for_a2 <= 834;
        o_index_for_a3 <= 874;
        o_index_for_a4 <= 1475;
        o_index_for_a5 <= 1571; 
        o_index_for_a6 <= 2304; 
    end
    324: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 71;
        o_index_for_a1 <= 277;
        o_index_for_a2 <= 835;
        o_index_for_a3 <= 875;
        o_index_for_a4 <= 1476;
        o_index_for_a5 <= 1572; 
        o_index_for_a6 <= 2304; 
    end
    325: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 72;
        o_index_for_a1 <= 278;
        o_index_for_a2 <= 836;
        o_index_for_a3 <= 876;
        o_index_for_a4 <= 1477;
        o_index_for_a5 <= 1573; 
        o_index_for_a6 <= 2304; 
    end
    326: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 73;
        o_index_for_a1 <= 279;
        o_index_for_a2 <= 837;
        o_index_for_a3 <= 877;
        o_index_for_a4 <= 1478;
        o_index_for_a5 <= 1574; 
        o_index_for_a6 <= 2304; 
    end
    327: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 74;
        o_index_for_a1 <= 280;
        o_index_for_a2 <= 838;
        o_index_for_a3 <= 878;
        o_index_for_a4 <= 1479;
        o_index_for_a5 <= 1575; 
        o_index_for_a6 <= 2304; 
    end
    328: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 75;
        o_index_for_a1 <= 281;
        o_index_for_a2 <= 839;
        o_index_for_a3 <= 879;
        o_index_for_a4 <= 1480;
        o_index_for_a5 <= 1576; 
        o_index_for_a6 <= 2304; 
    end
    329: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 76;
        o_index_for_a1 <= 282;
        o_index_for_a2 <= 840;
        o_index_for_a3 <= 880;
        o_index_for_a4 <= 1481;
        o_index_for_a5 <= 1577; 
        o_index_for_a6 <= 2304; 
    end
    330: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 77;
        o_index_for_a1 <= 283;
        o_index_for_a2 <= 841;
        o_index_for_a3 <= 881;
        o_index_for_a4 <= 1482;
        o_index_for_a5 <= 1578; 
        o_index_for_a6 <= 2304; 
    end
    331: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 78;
        o_index_for_a1 <= 284;
        o_index_for_a2 <= 842;
        o_index_for_a3 <= 882;
        o_index_for_a4 <= 1483;
        o_index_for_a5 <= 1579; 
        o_index_for_a6 <= 2304; 
    end
    332: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 79;
        o_index_for_a1 <= 285;
        o_index_for_a2 <= 843;
        o_index_for_a3 <= 883;
        o_index_for_a4 <= 1484;
        o_index_for_a5 <= 1580; 
        o_index_for_a6 <= 2304; 
    end
    333: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 80;
        o_index_for_a1 <= 286;
        o_index_for_a2 <= 844;
        o_index_for_a3 <= 884;
        o_index_for_a4 <= 1485;
        o_index_for_a5 <= 1581; 
        o_index_for_a6 <= 2304; 
    end
    334: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 81;
        o_index_for_a1 <= 287;
        o_index_for_a2 <= 845;
        o_index_for_a3 <= 885;
        o_index_for_a4 <= 1486;
        o_index_for_a5 <= 1582; 
        o_index_for_a6 <= 2304; 
    end
    335: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 82;
        o_index_for_a1 <= 192;
        o_index_for_a2 <= 846;
        o_index_for_a3 <= 886;
        o_index_for_a4 <= 1487;
        o_index_for_a5 <= 1583; 
        o_index_for_a6 <= 2304; 
    end
    336: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 83;
        o_index_for_a1 <= 193;
        o_index_for_a2 <= 847;
        o_index_for_a3 <= 887;
        o_index_for_a4 <= 1488;
        o_index_for_a5 <= 1584; 
        o_index_for_a6 <= 2304; 
    end
    337: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 84;
        o_index_for_a1 <= 194;
        o_index_for_a2 <= 848;
        o_index_for_a3 <= 888;
        o_index_for_a4 <= 1489;
        o_index_for_a5 <= 1585; 
        o_index_for_a6 <= 2304; 
    end
    338: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 85;
        o_index_for_a1 <= 195;
        o_index_for_a2 <= 849;
        o_index_for_a3 <= 889;
        o_index_for_a4 <= 1490;
        o_index_for_a5 <= 1586; 
        o_index_for_a6 <= 2304; 
    end
    339: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 86;
        o_index_for_a1 <= 196;
        o_index_for_a2 <= 850;
        o_index_for_a3 <= 890;
        o_index_for_a4 <= 1491;
        o_index_for_a5 <= 1587; 
        o_index_for_a6 <= 2304; 
    end
    340: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 87;
        o_index_for_a1 <= 197;
        o_index_for_a2 <= 851;
        o_index_for_a3 <= 891;
        o_index_for_a4 <= 1492;
        o_index_for_a5 <= 1588; 
        o_index_for_a6 <= 2304; 
    end
    341: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 88;
        o_index_for_a1 <= 198;
        o_index_for_a2 <= 852;
        o_index_for_a3 <= 892;
        o_index_for_a4 <= 1493;
        o_index_for_a5 <= 1589; 
        o_index_for_a6 <= 2304; 
    end
    342: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 89;
        o_index_for_a1 <= 199;
        o_index_for_a2 <= 853;
        o_index_for_a3 <= 893;
        o_index_for_a4 <= 1494;
        o_index_for_a5 <= 1590; 
        o_index_for_a6 <= 2304; 
    end
    343: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 90;
        o_index_for_a1 <= 200;
        o_index_for_a2 <= 854;
        o_index_for_a3 <= 894;
        o_index_for_a4 <= 1495;
        o_index_for_a5 <= 1591; 
        o_index_for_a6 <= 2304; 
    end
    344: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 91;
        o_index_for_a1 <= 201;
        o_index_for_a2 <= 855;
        o_index_for_a3 <= 895;
        o_index_for_a4 <= 1496;
        o_index_for_a5 <= 1592; 
        o_index_for_a6 <= 2304; 
    end
    345: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 92;
        o_index_for_a1 <= 202;
        o_index_for_a2 <= 856;
        o_index_for_a3 <= 896;
        o_index_for_a4 <= 1497;
        o_index_for_a5 <= 1593; 
        o_index_for_a6 <= 2304; 
    end
    346: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 93;
        o_index_for_a1 <= 203;
        o_index_for_a2 <= 857;
        o_index_for_a3 <= 897;
        o_index_for_a4 <= 1498;
        o_index_for_a5 <= 1594; 
        o_index_for_a6 <= 2304; 
    end
    347: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 94;
        o_index_for_a1 <= 204;
        o_index_for_a2 <= 858;
        o_index_for_a3 <= 898;
        o_index_for_a4 <= 1499;
        o_index_for_a5 <= 1595; 
        o_index_for_a6 <= 2304; 
    end
    348: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 95;
        o_index_for_a1 <= 205;
        o_index_for_a2 <= 859;
        o_index_for_a3 <= 899;
        o_index_for_a4 <= 1500;
        o_index_for_a5 <= 1596; 
        o_index_for_a6 <= 2304; 
    end
    349: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 0;
        o_index_for_a1 <= 206;
        o_index_for_a2 <= 860;
        o_index_for_a3 <= 900;
        o_index_for_a4 <= 1501;
        o_index_for_a5 <= 1597; 
        o_index_for_a6 <= 2304; 
    end
    350: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 1;
        o_index_for_a1 <= 207;
        o_index_for_a2 <= 861;
        o_index_for_a3 <= 901;
        o_index_for_a4 <= 1502;
        o_index_for_a5 <= 1598; 
        o_index_for_a6 <= 2304; 
    end
    351: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 2;
        o_index_for_a1 <= 208;
        o_index_for_a2 <= 862;
        o_index_for_a3 <= 902;
        o_index_for_a4 <= 1503;
        o_index_for_a5 <= 1599; 
        o_index_for_a6 <= 2304; 
    end
    352: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 3;
        o_index_for_a1 <= 209;
        o_index_for_a2 <= 863;
        o_index_for_a3 <= 903;
        o_index_for_a4 <= 1504;
        o_index_for_a5 <= 1600; 
        o_index_for_a6 <= 2304; 
    end
    353: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 4;
        o_index_for_a1 <= 210;
        o_index_for_a2 <= 768;
        o_index_for_a3 <= 904;
        o_index_for_a4 <= 1505;
        o_index_for_a5 <= 1601; 
        o_index_for_a6 <= 2304; 
    end
    354: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 5;
        o_index_for_a1 <= 211;
        o_index_for_a2 <= 769;
        o_index_for_a3 <= 905;
        o_index_for_a4 <= 1506;
        o_index_for_a5 <= 1602; 
        o_index_for_a6 <= 2304; 
    end
    355: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 6;
        o_index_for_a1 <= 212;
        o_index_for_a2 <= 770;
        o_index_for_a3 <= 906;
        o_index_for_a4 <= 1507;
        o_index_for_a5 <= 1603; 
        o_index_for_a6 <= 2304; 
    end
    356: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 7;
        o_index_for_a1 <= 213;
        o_index_for_a2 <= 771;
        o_index_for_a3 <= 907;
        o_index_for_a4 <= 1508;
        o_index_for_a5 <= 1604; 
        o_index_for_a6 <= 2304; 
    end
    357: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 8;
        o_index_for_a1 <= 214;
        o_index_for_a2 <= 772;
        o_index_for_a3 <= 908;
        o_index_for_a4 <= 1509;
        o_index_for_a5 <= 1605; 
        o_index_for_a6 <= 2304; 
    end
    358: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 9;
        o_index_for_a1 <= 215;
        o_index_for_a2 <= 773;
        o_index_for_a3 <= 909;
        o_index_for_a4 <= 1510;
        o_index_for_a5 <= 1606; 
        o_index_for_a6 <= 2304; 
    end
    359: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 10;
        o_index_for_a1 <= 216;
        o_index_for_a2 <= 774;
        o_index_for_a3 <= 910;
        o_index_for_a4 <= 1511;
        o_index_for_a5 <= 1607; 
        o_index_for_a6 <= 2304; 
    end
    360: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 11;
        o_index_for_a1 <= 217;
        o_index_for_a2 <= 775;
        o_index_for_a3 <= 911;
        o_index_for_a4 <= 1512;
        o_index_for_a5 <= 1608; 
        o_index_for_a6 <= 2304; 
    end
    361: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 12;
        o_index_for_a1 <= 218;
        o_index_for_a2 <= 776;
        o_index_for_a3 <= 912;
        o_index_for_a4 <= 1513;
        o_index_for_a5 <= 1609; 
        o_index_for_a6 <= 2304; 
    end
    362: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 13;
        o_index_for_a1 <= 219;
        o_index_for_a2 <= 777;
        o_index_for_a3 <= 913;
        o_index_for_a4 <= 1514;
        o_index_for_a5 <= 1610; 
        o_index_for_a6 <= 2304; 
    end
    363: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 14;
        o_index_for_a1 <= 220;
        o_index_for_a2 <= 778;
        o_index_for_a3 <= 914;
        o_index_for_a4 <= 1515;
        o_index_for_a5 <= 1611; 
        o_index_for_a6 <= 2304; 
    end
    364: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 15;
        o_index_for_a1 <= 221;
        o_index_for_a2 <= 779;
        o_index_for_a3 <= 915;
        o_index_for_a4 <= 1516;
        o_index_for_a5 <= 1612; 
        o_index_for_a6 <= 2304; 
    end
    365: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 16;
        o_index_for_a1 <= 222;
        o_index_for_a2 <= 780;
        o_index_for_a3 <= 916;
        o_index_for_a4 <= 1517;
        o_index_for_a5 <= 1613; 
        o_index_for_a6 <= 2304; 
    end
    366: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 17;
        o_index_for_a1 <= 223;
        o_index_for_a2 <= 781;
        o_index_for_a3 <= 917;
        o_index_for_a4 <= 1518;
        o_index_for_a5 <= 1614; 
        o_index_for_a6 <= 2304; 
    end
    367: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 18;
        o_index_for_a1 <= 224;
        o_index_for_a2 <= 782;
        o_index_for_a3 <= 918;
        o_index_for_a4 <= 1519;
        o_index_for_a5 <= 1615; 
        o_index_for_a6 <= 2304; 
    end
    368: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 19;
        o_index_for_a1 <= 225;
        o_index_for_a2 <= 783;
        o_index_for_a3 <= 919;
        o_index_for_a4 <= 1520;
        o_index_for_a5 <= 1616; 
        o_index_for_a6 <= 2304; 
    end
    369: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 20;
        o_index_for_a1 <= 226;
        o_index_for_a2 <= 784;
        o_index_for_a3 <= 920;
        o_index_for_a4 <= 1521;
        o_index_for_a5 <= 1617; 
        o_index_for_a6 <= 2304; 
    end
    370: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 21;
        o_index_for_a1 <= 227;
        o_index_for_a2 <= 785;
        o_index_for_a3 <= 921;
        o_index_for_a4 <= 1522;
        o_index_for_a5 <= 1618; 
        o_index_for_a6 <= 2304; 
    end
    371: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 22;
        o_index_for_a1 <= 228;
        o_index_for_a2 <= 786;
        o_index_for_a3 <= 922;
        o_index_for_a4 <= 1523;
        o_index_for_a5 <= 1619; 
        o_index_for_a6 <= 2304; 
    end
    372: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 23;
        o_index_for_a1 <= 229;
        o_index_for_a2 <= 787;
        o_index_for_a3 <= 923;
        o_index_for_a4 <= 1524;
        o_index_for_a5 <= 1620; 
        o_index_for_a6 <= 2304; 
    end
    373: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 24;
        o_index_for_a1 <= 230;
        o_index_for_a2 <= 788;
        o_index_for_a3 <= 924;
        o_index_for_a4 <= 1525;
        o_index_for_a5 <= 1621; 
        o_index_for_a6 <= 2304; 
    end
    374: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 25;
        o_index_for_a1 <= 231;
        o_index_for_a2 <= 789;
        o_index_for_a3 <= 925;
        o_index_for_a4 <= 1526;
        o_index_for_a5 <= 1622; 
        o_index_for_a6 <= 2304; 
    end
    375: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 26;
        o_index_for_a1 <= 232;
        o_index_for_a2 <= 790;
        o_index_for_a3 <= 926;
        o_index_for_a4 <= 1527;
        o_index_for_a5 <= 1623; 
        o_index_for_a6 <= 2304; 
    end
    376: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 27;
        o_index_for_a1 <= 233;
        o_index_for_a2 <= 791;
        o_index_for_a3 <= 927;
        o_index_for_a4 <= 1528;
        o_index_for_a5 <= 1624; 
        o_index_for_a6 <= 2304; 
    end
    377: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 28;
        o_index_for_a1 <= 234;
        o_index_for_a2 <= 792;
        o_index_for_a3 <= 928;
        o_index_for_a4 <= 1529;
        o_index_for_a5 <= 1625; 
        o_index_for_a6 <= 2304; 
    end
    378: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 29;
        o_index_for_a1 <= 235;
        o_index_for_a2 <= 793;
        o_index_for_a3 <= 929;
        o_index_for_a4 <= 1530;
        o_index_for_a5 <= 1626; 
        o_index_for_a6 <= 2304; 
    end
    379: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 30;
        o_index_for_a1 <= 236;
        o_index_for_a2 <= 794;
        o_index_for_a3 <= 930;
        o_index_for_a4 <= 1531;
        o_index_for_a5 <= 1627; 
        o_index_for_a6 <= 2304; 
    end
    380: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 31;
        o_index_for_a1 <= 237;
        o_index_for_a2 <= 795;
        o_index_for_a3 <= 931;
        o_index_for_a4 <= 1532;
        o_index_for_a5 <= 1628; 
        o_index_for_a6 <= 2304; 
    end
    381: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 32;
        o_index_for_a1 <= 238;
        o_index_for_a2 <= 796;
        o_index_for_a3 <= 932;
        o_index_for_a4 <= 1533;
        o_index_for_a5 <= 1629; 
        o_index_for_a6 <= 2304; 
    end
    382: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 33;
        o_index_for_a1 <= 239;
        o_index_for_a2 <= 797;
        o_index_for_a3 <= 933;
        o_index_for_a4 <= 1534;
        o_index_for_a5 <= 1630; 
        o_index_for_a6 <= 2304; 
    end
    383: begin
        o_branch_for_a0 <= 0;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 1;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 34;
        o_index_for_a1 <= 240;
        o_index_for_a2 <= 798;
        o_index_for_a3 <= 934;
        o_index_for_a4 <= 1535;
        o_index_for_a5 <= 1631; 
        o_index_for_a6 <= 2304; 
    end
    384: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 249;
        o_index_for_a1 <= 588;
        o_index_for_a2 <= 919;
        o_index_for_a3 <= 984;
        o_index_for_a4 <= 1536;
        o_index_for_a5 <= 1632; 
        o_index_for_a6 <= 2304; 
    end
    385: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 250;
        o_index_for_a1 <= 589;
        o_index_for_a2 <= 920;
        o_index_for_a3 <= 985;
        o_index_for_a4 <= 1537;
        o_index_for_a5 <= 1633; 
        o_index_for_a6 <= 2304; 
    end
    386: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 251;
        o_index_for_a1 <= 590;
        o_index_for_a2 <= 921;
        o_index_for_a3 <= 986;
        o_index_for_a4 <= 1538;
        o_index_for_a5 <= 1634; 
        o_index_for_a6 <= 2304; 
    end
    387: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 252;
        o_index_for_a1 <= 591;
        o_index_for_a2 <= 922;
        o_index_for_a3 <= 987;
        o_index_for_a4 <= 1539;
        o_index_for_a5 <= 1635; 
        o_index_for_a6 <= 2304; 
    end
    388: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 253;
        o_index_for_a1 <= 592;
        o_index_for_a2 <= 923;
        o_index_for_a3 <= 988;
        o_index_for_a4 <= 1540;
        o_index_for_a5 <= 1636; 
        o_index_for_a6 <= 2304; 
    end
    389: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 254;
        o_index_for_a1 <= 593;
        o_index_for_a2 <= 924;
        o_index_for_a3 <= 989;
        o_index_for_a4 <= 1541;
        o_index_for_a5 <= 1637; 
        o_index_for_a6 <= 2304; 
    end
    390: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 255;
        o_index_for_a1 <= 594;
        o_index_for_a2 <= 925;
        o_index_for_a3 <= 990;
        o_index_for_a4 <= 1542;
        o_index_for_a5 <= 1638; 
        o_index_for_a6 <= 2304; 
    end
    391: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 256;
        o_index_for_a1 <= 595;
        o_index_for_a2 <= 926;
        o_index_for_a3 <= 991;
        o_index_for_a4 <= 1543;
        o_index_for_a5 <= 1639; 
        o_index_for_a6 <= 2304; 
    end
    392: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 257;
        o_index_for_a1 <= 596;
        o_index_for_a2 <= 927;
        o_index_for_a3 <= 992;
        o_index_for_a4 <= 1544;
        o_index_for_a5 <= 1640; 
        o_index_for_a6 <= 2304; 
    end
    393: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 258;
        o_index_for_a1 <= 597;
        o_index_for_a2 <= 928;
        o_index_for_a3 <= 993;
        o_index_for_a4 <= 1545;
        o_index_for_a5 <= 1641; 
        o_index_for_a6 <= 2304; 
    end
    394: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 259;
        o_index_for_a1 <= 598;
        o_index_for_a2 <= 929;
        o_index_for_a3 <= 994;
        o_index_for_a4 <= 1546;
        o_index_for_a5 <= 1642; 
        o_index_for_a6 <= 2304; 
    end
    395: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 260;
        o_index_for_a1 <= 599;
        o_index_for_a2 <= 930;
        o_index_for_a3 <= 995;
        o_index_for_a4 <= 1547;
        o_index_for_a5 <= 1643; 
        o_index_for_a6 <= 2304; 
    end
    396: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 261;
        o_index_for_a1 <= 600;
        o_index_for_a2 <= 931;
        o_index_for_a3 <= 996;
        o_index_for_a4 <= 1548;
        o_index_for_a5 <= 1644; 
        o_index_for_a6 <= 2304; 
    end
    397: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 262;
        o_index_for_a1 <= 601;
        o_index_for_a2 <= 932;
        o_index_for_a3 <= 997;
        o_index_for_a4 <= 1549;
        o_index_for_a5 <= 1645; 
        o_index_for_a6 <= 2304; 
    end
    398: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 263;
        o_index_for_a1 <= 602;
        o_index_for_a2 <= 933;
        o_index_for_a3 <= 998;
        o_index_for_a4 <= 1550;
        o_index_for_a5 <= 1646; 
        o_index_for_a6 <= 2304; 
    end
    399: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 264;
        o_index_for_a1 <= 603;
        o_index_for_a2 <= 934;
        o_index_for_a3 <= 999;
        o_index_for_a4 <= 1551;
        o_index_for_a5 <= 1647; 
        o_index_for_a6 <= 2304; 
    end
    400: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 265;
        o_index_for_a1 <= 604;
        o_index_for_a2 <= 935;
        o_index_for_a3 <= 1000;
        o_index_for_a4 <= 1552;
        o_index_for_a5 <= 1648; 
        o_index_for_a6 <= 2304; 
    end
    401: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 266;
        o_index_for_a1 <= 605;
        o_index_for_a2 <= 936;
        o_index_for_a3 <= 1001;
        o_index_for_a4 <= 1553;
        o_index_for_a5 <= 1649; 
        o_index_for_a6 <= 2304; 
    end
    402: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 267;
        o_index_for_a1 <= 606;
        o_index_for_a2 <= 937;
        o_index_for_a3 <= 1002;
        o_index_for_a4 <= 1554;
        o_index_for_a5 <= 1650; 
        o_index_for_a6 <= 2304; 
    end
    403: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 268;
        o_index_for_a1 <= 607;
        o_index_for_a2 <= 938;
        o_index_for_a3 <= 1003;
        o_index_for_a4 <= 1555;
        o_index_for_a5 <= 1651; 
        o_index_for_a6 <= 2304; 
    end
    404: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 269;
        o_index_for_a1 <= 608;
        o_index_for_a2 <= 939;
        o_index_for_a3 <= 1004;
        o_index_for_a4 <= 1556;
        o_index_for_a5 <= 1652; 
        o_index_for_a6 <= 2304; 
    end
    405: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 270;
        o_index_for_a1 <= 609;
        o_index_for_a2 <= 940;
        o_index_for_a3 <= 1005;
        o_index_for_a4 <= 1557;
        o_index_for_a5 <= 1653; 
        o_index_for_a6 <= 2304; 
    end
    406: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 271;
        o_index_for_a1 <= 610;
        o_index_for_a2 <= 941;
        o_index_for_a3 <= 1006;
        o_index_for_a4 <= 1558;
        o_index_for_a5 <= 1654; 
        o_index_for_a6 <= 2304; 
    end
    407: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 272;
        o_index_for_a1 <= 611;
        o_index_for_a2 <= 942;
        o_index_for_a3 <= 1007;
        o_index_for_a4 <= 1559;
        o_index_for_a5 <= 1655; 
        o_index_for_a6 <= 2304; 
    end
    408: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 273;
        o_index_for_a1 <= 612;
        o_index_for_a2 <= 943;
        o_index_for_a3 <= 1008;
        o_index_for_a4 <= 1560;
        o_index_for_a5 <= 1656; 
        o_index_for_a6 <= 2304; 
    end
    409: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 274;
        o_index_for_a1 <= 613;
        o_index_for_a2 <= 944;
        o_index_for_a3 <= 1009;
        o_index_for_a4 <= 1561;
        o_index_for_a5 <= 1657; 
        o_index_for_a6 <= 2304; 
    end
    410: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 275;
        o_index_for_a1 <= 614;
        o_index_for_a2 <= 945;
        o_index_for_a3 <= 1010;
        o_index_for_a4 <= 1562;
        o_index_for_a5 <= 1658; 
        o_index_for_a6 <= 2304; 
    end
    411: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 276;
        o_index_for_a1 <= 615;
        o_index_for_a2 <= 946;
        o_index_for_a3 <= 1011;
        o_index_for_a4 <= 1563;
        o_index_for_a5 <= 1659; 
        o_index_for_a6 <= 2304; 
    end
    412: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 277;
        o_index_for_a1 <= 616;
        o_index_for_a2 <= 947;
        o_index_for_a3 <= 1012;
        o_index_for_a4 <= 1564;
        o_index_for_a5 <= 1660; 
        o_index_for_a6 <= 2304; 
    end
    413: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 278;
        o_index_for_a1 <= 617;
        o_index_for_a2 <= 948;
        o_index_for_a3 <= 1013;
        o_index_for_a4 <= 1565;
        o_index_for_a5 <= 1661; 
        o_index_for_a6 <= 2304; 
    end
    414: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 279;
        o_index_for_a1 <= 618;
        o_index_for_a2 <= 949;
        o_index_for_a3 <= 1014;
        o_index_for_a4 <= 1566;
        o_index_for_a5 <= 1662; 
        o_index_for_a6 <= 2304; 
    end
    415: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 280;
        o_index_for_a1 <= 619;
        o_index_for_a2 <= 950;
        o_index_for_a3 <= 1015;
        o_index_for_a4 <= 1567;
        o_index_for_a5 <= 1663; 
        o_index_for_a6 <= 2304; 
    end
    416: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 281;
        o_index_for_a1 <= 620;
        o_index_for_a2 <= 951;
        o_index_for_a3 <= 1016;
        o_index_for_a4 <= 1568;
        o_index_for_a5 <= 1664; 
        o_index_for_a6 <= 2304; 
    end
    417: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 282;
        o_index_for_a1 <= 621;
        o_index_for_a2 <= 952;
        o_index_for_a3 <= 1017;
        o_index_for_a4 <= 1569;
        o_index_for_a5 <= 1665; 
        o_index_for_a6 <= 2304; 
    end
    418: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 283;
        o_index_for_a1 <= 622;
        o_index_for_a2 <= 953;
        o_index_for_a3 <= 1018;
        o_index_for_a4 <= 1570;
        o_index_for_a5 <= 1666; 
        o_index_for_a6 <= 2304; 
    end
    419: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 284;
        o_index_for_a1 <= 623;
        o_index_for_a2 <= 954;
        o_index_for_a3 <= 1019;
        o_index_for_a4 <= 1571;
        o_index_for_a5 <= 1667; 
        o_index_for_a6 <= 2304; 
    end
    420: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 285;
        o_index_for_a1 <= 624;
        o_index_for_a2 <= 955;
        o_index_for_a3 <= 1020;
        o_index_for_a4 <= 1572;
        o_index_for_a5 <= 1668; 
        o_index_for_a6 <= 2304; 
    end
    421: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 286;
        o_index_for_a1 <= 625;
        o_index_for_a2 <= 956;
        o_index_for_a3 <= 1021;
        o_index_for_a4 <= 1573;
        o_index_for_a5 <= 1669; 
        o_index_for_a6 <= 2304; 
    end
    422: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 287;
        o_index_for_a1 <= 626;
        o_index_for_a2 <= 957;
        o_index_for_a3 <= 1022;
        o_index_for_a4 <= 1574;
        o_index_for_a5 <= 1670; 
        o_index_for_a6 <= 2304; 
    end
    423: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 192;
        o_index_for_a1 <= 627;
        o_index_for_a2 <= 958;
        o_index_for_a3 <= 1023;
        o_index_for_a4 <= 1575;
        o_index_for_a5 <= 1671; 
        o_index_for_a6 <= 2304; 
    end
    424: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 193;
        o_index_for_a1 <= 628;
        o_index_for_a2 <= 959;
        o_index_for_a3 <= 1024;
        o_index_for_a4 <= 1576;
        o_index_for_a5 <= 1672; 
        o_index_for_a6 <= 2304; 
    end
    425: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 194;
        o_index_for_a1 <= 629;
        o_index_for_a2 <= 864;
        o_index_for_a3 <= 1025;
        o_index_for_a4 <= 1577;
        o_index_for_a5 <= 1673; 
        o_index_for_a6 <= 2304; 
    end
    426: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 195;
        o_index_for_a1 <= 630;
        o_index_for_a2 <= 865;
        o_index_for_a3 <= 1026;
        o_index_for_a4 <= 1578;
        o_index_for_a5 <= 1674; 
        o_index_for_a6 <= 2304; 
    end
    427: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 196;
        o_index_for_a1 <= 631;
        o_index_for_a2 <= 866;
        o_index_for_a3 <= 1027;
        o_index_for_a4 <= 1579;
        o_index_for_a5 <= 1675; 
        o_index_for_a6 <= 2304; 
    end
    428: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 197;
        o_index_for_a1 <= 632;
        o_index_for_a2 <= 867;
        o_index_for_a3 <= 1028;
        o_index_for_a4 <= 1580;
        o_index_for_a5 <= 1676; 
        o_index_for_a6 <= 2304; 
    end
    429: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 198;
        o_index_for_a1 <= 633;
        o_index_for_a2 <= 868;
        o_index_for_a3 <= 1029;
        o_index_for_a4 <= 1581;
        o_index_for_a5 <= 1677; 
        o_index_for_a6 <= 2304; 
    end
    430: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 199;
        o_index_for_a1 <= 634;
        o_index_for_a2 <= 869;
        o_index_for_a3 <= 1030;
        o_index_for_a4 <= 1582;
        o_index_for_a5 <= 1678; 
        o_index_for_a6 <= 2304; 
    end
    431: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 200;
        o_index_for_a1 <= 635;
        o_index_for_a2 <= 870;
        o_index_for_a3 <= 1031;
        o_index_for_a4 <= 1583;
        o_index_for_a5 <= 1679; 
        o_index_for_a6 <= 2304; 
    end
    432: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 201;
        o_index_for_a1 <= 636;
        o_index_for_a2 <= 871;
        o_index_for_a3 <= 1032;
        o_index_for_a4 <= 1584;
        o_index_for_a5 <= 1680; 
        o_index_for_a6 <= 2304; 
    end
    433: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 202;
        o_index_for_a1 <= 637;
        o_index_for_a2 <= 872;
        o_index_for_a3 <= 1033;
        o_index_for_a4 <= 1585;
        o_index_for_a5 <= 1681; 
        o_index_for_a6 <= 2304; 
    end
    434: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 203;
        o_index_for_a1 <= 638;
        o_index_for_a2 <= 873;
        o_index_for_a3 <= 1034;
        o_index_for_a4 <= 1586;
        o_index_for_a5 <= 1682; 
        o_index_for_a6 <= 2304; 
    end
    435: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 204;
        o_index_for_a1 <= 639;
        o_index_for_a2 <= 874;
        o_index_for_a3 <= 1035;
        o_index_for_a4 <= 1587;
        o_index_for_a5 <= 1683; 
        o_index_for_a6 <= 2304; 
    end
    436: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 205;
        o_index_for_a1 <= 640;
        o_index_for_a2 <= 875;
        o_index_for_a3 <= 1036;
        o_index_for_a4 <= 1588;
        o_index_for_a5 <= 1684; 
        o_index_for_a6 <= 2304; 
    end
    437: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 206;
        o_index_for_a1 <= 641;
        o_index_for_a2 <= 876;
        o_index_for_a3 <= 1037;
        o_index_for_a4 <= 1589;
        o_index_for_a5 <= 1685; 
        o_index_for_a6 <= 2304; 
    end
    438: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 207;
        o_index_for_a1 <= 642;
        o_index_for_a2 <= 877;
        o_index_for_a3 <= 1038;
        o_index_for_a4 <= 1590;
        o_index_for_a5 <= 1686; 
        o_index_for_a6 <= 2304; 
    end
    439: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 208;
        o_index_for_a1 <= 643;
        o_index_for_a2 <= 878;
        o_index_for_a3 <= 1039;
        o_index_for_a4 <= 1591;
        o_index_for_a5 <= 1687; 
        o_index_for_a6 <= 2304; 
    end
    440: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 209;
        o_index_for_a1 <= 644;
        o_index_for_a2 <= 879;
        o_index_for_a3 <= 1040;
        o_index_for_a4 <= 1592;
        o_index_for_a5 <= 1688; 
        o_index_for_a6 <= 2304; 
    end
    441: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 210;
        o_index_for_a1 <= 645;
        o_index_for_a2 <= 880;
        o_index_for_a3 <= 1041;
        o_index_for_a4 <= 1593;
        o_index_for_a5 <= 1689; 
        o_index_for_a6 <= 2304; 
    end
    442: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 211;
        o_index_for_a1 <= 646;
        o_index_for_a2 <= 881;
        o_index_for_a3 <= 1042;
        o_index_for_a4 <= 1594;
        o_index_for_a5 <= 1690; 
        o_index_for_a6 <= 2304; 
    end
    443: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 212;
        o_index_for_a1 <= 647;
        o_index_for_a2 <= 882;
        o_index_for_a3 <= 1043;
        o_index_for_a4 <= 1595;
        o_index_for_a5 <= 1691; 
        o_index_for_a6 <= 2304; 
    end
    444: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 213;
        o_index_for_a1 <= 648;
        o_index_for_a2 <= 883;
        o_index_for_a3 <= 1044;
        o_index_for_a4 <= 1596;
        o_index_for_a5 <= 1692; 
        o_index_for_a6 <= 2304; 
    end
    445: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 214;
        o_index_for_a1 <= 649;
        o_index_for_a2 <= 884;
        o_index_for_a3 <= 1045;
        o_index_for_a4 <= 1597;
        o_index_for_a5 <= 1693; 
        o_index_for_a6 <= 2304; 
    end
    446: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 215;
        o_index_for_a1 <= 650;
        o_index_for_a2 <= 885;
        o_index_for_a3 <= 1046;
        o_index_for_a4 <= 1598;
        o_index_for_a5 <= 1694; 
        o_index_for_a6 <= 2304; 
    end
    447: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 216;
        o_index_for_a1 <= 651;
        o_index_for_a2 <= 886;
        o_index_for_a3 <= 1047;
        o_index_for_a4 <= 1599;
        o_index_for_a5 <= 1695; 
        o_index_for_a6 <= 2304; 
    end
    448: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 217;
        o_index_for_a1 <= 652;
        o_index_for_a2 <= 887;
        o_index_for_a3 <= 1048;
        o_index_for_a4 <= 1600;
        o_index_for_a5 <= 1696; 
        o_index_for_a6 <= 2304; 
    end
    449: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 218;
        o_index_for_a1 <= 653;
        o_index_for_a2 <= 888;
        o_index_for_a3 <= 1049;
        o_index_for_a4 <= 1601;
        o_index_for_a5 <= 1697; 
        o_index_for_a6 <= 2304; 
    end
    450: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 219;
        o_index_for_a1 <= 654;
        o_index_for_a2 <= 889;
        o_index_for_a3 <= 1050;
        o_index_for_a4 <= 1602;
        o_index_for_a5 <= 1698; 
        o_index_for_a6 <= 2304; 
    end
    451: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 220;
        o_index_for_a1 <= 655;
        o_index_for_a2 <= 890;
        o_index_for_a3 <= 1051;
        o_index_for_a4 <= 1603;
        o_index_for_a5 <= 1699; 
        o_index_for_a6 <= 2304; 
    end
    452: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 221;
        o_index_for_a1 <= 656;
        o_index_for_a2 <= 891;
        o_index_for_a3 <= 1052;
        o_index_for_a4 <= 1604;
        o_index_for_a5 <= 1700; 
        o_index_for_a6 <= 2304; 
    end
    453: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 222;
        o_index_for_a1 <= 657;
        o_index_for_a2 <= 892;
        o_index_for_a3 <= 1053;
        o_index_for_a4 <= 1605;
        o_index_for_a5 <= 1701; 
        o_index_for_a6 <= 2304; 
    end
    454: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 223;
        o_index_for_a1 <= 658;
        o_index_for_a2 <= 893;
        o_index_for_a3 <= 1054;
        o_index_for_a4 <= 1606;
        o_index_for_a5 <= 1702; 
        o_index_for_a6 <= 2304; 
    end
    455: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 224;
        o_index_for_a1 <= 659;
        o_index_for_a2 <= 894;
        o_index_for_a3 <= 1055;
        o_index_for_a4 <= 1607;
        o_index_for_a5 <= 1703; 
        o_index_for_a6 <= 2304; 
    end
    456: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 225;
        o_index_for_a1 <= 660;
        o_index_for_a2 <= 895;
        o_index_for_a3 <= 960;
        o_index_for_a4 <= 1608;
        o_index_for_a5 <= 1704; 
        o_index_for_a6 <= 2304; 
    end
    457: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 226;
        o_index_for_a1 <= 661;
        o_index_for_a2 <= 896;
        o_index_for_a3 <= 961;
        o_index_for_a4 <= 1609;
        o_index_for_a5 <= 1705; 
        o_index_for_a6 <= 2304; 
    end
    458: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 227;
        o_index_for_a1 <= 662;
        o_index_for_a2 <= 897;
        o_index_for_a3 <= 962;
        o_index_for_a4 <= 1610;
        o_index_for_a5 <= 1706; 
        o_index_for_a6 <= 2304; 
    end
    459: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 228;
        o_index_for_a1 <= 663;
        o_index_for_a2 <= 898;
        o_index_for_a3 <= 963;
        o_index_for_a4 <= 1611;
        o_index_for_a5 <= 1707; 
        o_index_for_a6 <= 2304; 
    end
    460: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 229;
        o_index_for_a1 <= 664;
        o_index_for_a2 <= 899;
        o_index_for_a3 <= 964;
        o_index_for_a4 <= 1612;
        o_index_for_a5 <= 1708; 
        o_index_for_a6 <= 2304; 
    end
    461: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 230;
        o_index_for_a1 <= 665;
        o_index_for_a2 <= 900;
        o_index_for_a3 <= 965;
        o_index_for_a4 <= 1613;
        o_index_for_a5 <= 1709; 
        o_index_for_a6 <= 2304; 
    end
    462: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 231;
        o_index_for_a1 <= 666;
        o_index_for_a2 <= 901;
        o_index_for_a3 <= 966;
        o_index_for_a4 <= 1614;
        o_index_for_a5 <= 1710; 
        o_index_for_a6 <= 2304; 
    end
    463: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 232;
        o_index_for_a1 <= 667;
        o_index_for_a2 <= 902;
        o_index_for_a3 <= 967;
        o_index_for_a4 <= 1615;
        o_index_for_a5 <= 1711; 
        o_index_for_a6 <= 2304; 
    end
    464: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 233;
        o_index_for_a1 <= 668;
        o_index_for_a2 <= 903;
        o_index_for_a3 <= 968;
        o_index_for_a4 <= 1616;
        o_index_for_a5 <= 1712; 
        o_index_for_a6 <= 2304; 
    end
    465: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 234;
        o_index_for_a1 <= 669;
        o_index_for_a2 <= 904;
        o_index_for_a3 <= 969;
        o_index_for_a4 <= 1617;
        o_index_for_a5 <= 1713; 
        o_index_for_a6 <= 2304; 
    end
    466: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 235;
        o_index_for_a1 <= 670;
        o_index_for_a2 <= 905;
        o_index_for_a3 <= 970;
        o_index_for_a4 <= 1618;
        o_index_for_a5 <= 1714; 
        o_index_for_a6 <= 2304; 
    end
    467: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 236;
        o_index_for_a1 <= 671;
        o_index_for_a2 <= 906;
        o_index_for_a3 <= 971;
        o_index_for_a4 <= 1619;
        o_index_for_a5 <= 1715; 
        o_index_for_a6 <= 2304; 
    end
    468: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 237;
        o_index_for_a1 <= 576;
        o_index_for_a2 <= 907;
        o_index_for_a3 <= 972;
        o_index_for_a4 <= 1620;
        o_index_for_a5 <= 1716; 
        o_index_for_a6 <= 2304; 
    end
    469: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 238;
        o_index_for_a1 <= 577;
        o_index_for_a2 <= 908;
        o_index_for_a3 <= 973;
        o_index_for_a4 <= 1621;
        o_index_for_a5 <= 1717; 
        o_index_for_a6 <= 2304; 
    end
    470: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 239;
        o_index_for_a1 <= 578;
        o_index_for_a2 <= 909;
        o_index_for_a3 <= 974;
        o_index_for_a4 <= 1622;
        o_index_for_a5 <= 1718; 
        o_index_for_a6 <= 2304; 
    end
    471: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 240;
        o_index_for_a1 <= 579;
        o_index_for_a2 <= 910;
        o_index_for_a3 <= 975;
        o_index_for_a4 <= 1623;
        o_index_for_a5 <= 1719; 
        o_index_for_a6 <= 2304; 
    end
    472: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 241;
        o_index_for_a1 <= 580;
        o_index_for_a2 <= 911;
        o_index_for_a3 <= 976;
        o_index_for_a4 <= 1624;
        o_index_for_a5 <= 1720; 
        o_index_for_a6 <= 2304; 
    end
    473: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 242;
        o_index_for_a1 <= 581;
        o_index_for_a2 <= 912;
        o_index_for_a3 <= 977;
        o_index_for_a4 <= 1625;
        o_index_for_a5 <= 1721; 
        o_index_for_a6 <= 2304; 
    end
    474: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 243;
        o_index_for_a1 <= 582;
        o_index_for_a2 <= 913;
        o_index_for_a3 <= 978;
        o_index_for_a4 <= 1626;
        o_index_for_a5 <= 1722; 
        o_index_for_a6 <= 2304; 
    end
    475: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 244;
        o_index_for_a1 <= 583;
        o_index_for_a2 <= 914;
        o_index_for_a3 <= 979;
        o_index_for_a4 <= 1627;
        o_index_for_a5 <= 1723; 
        o_index_for_a6 <= 2304; 
    end
    476: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 245;
        o_index_for_a1 <= 584;
        o_index_for_a2 <= 915;
        o_index_for_a3 <= 980;
        o_index_for_a4 <= 1628;
        o_index_for_a5 <= 1724; 
        o_index_for_a6 <= 2304; 
    end
    477: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 246;
        o_index_for_a1 <= 585;
        o_index_for_a2 <= 916;
        o_index_for_a3 <= 981;
        o_index_for_a4 <= 1629;
        o_index_for_a5 <= 1725; 
        o_index_for_a6 <= 2304; 
    end
    478: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 247;
        o_index_for_a1 <= 586;
        o_index_for_a2 <= 917;
        o_index_for_a3 <= 982;
        o_index_for_a4 <= 1630;
        o_index_for_a5 <= 1726; 
        o_index_for_a6 <= 2304; 
    end
    479: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 0;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 248;
        o_index_for_a1 <= 587;
        o_index_for_a2 <= 918;
        o_index_for_a3 <= 983;
        o_index_for_a4 <= 1631;
        o_index_for_a5 <= 1727; 
        o_index_for_a6 <= 2304; 
    end
    480: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 434;
        o_index_for_a1 <= 536;
        o_index_for_a2 <= 686;
        o_index_for_a3 <= 1073;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 1632; 
        o_index_for_a6 <= 1728; 
    end
    481: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 435;
        o_index_for_a1 <= 537;
        o_index_for_a2 <= 687;
        o_index_for_a3 <= 1074;
        o_index_for_a4 <= 1153;
        o_index_for_a5 <= 1633; 
        o_index_for_a6 <= 1729; 
    end
    482: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 436;
        o_index_for_a1 <= 538;
        o_index_for_a2 <= 688;
        o_index_for_a3 <= 1075;
        o_index_for_a4 <= 1154;
        o_index_for_a5 <= 1634; 
        o_index_for_a6 <= 1730; 
    end
    483: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 437;
        o_index_for_a1 <= 539;
        o_index_for_a2 <= 689;
        o_index_for_a3 <= 1076;
        o_index_for_a4 <= 1155;
        o_index_for_a5 <= 1635; 
        o_index_for_a6 <= 1731; 
    end
    484: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 438;
        o_index_for_a1 <= 540;
        o_index_for_a2 <= 690;
        o_index_for_a3 <= 1077;
        o_index_for_a4 <= 1156;
        o_index_for_a5 <= 1636; 
        o_index_for_a6 <= 1732; 
    end
    485: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 439;
        o_index_for_a1 <= 541;
        o_index_for_a2 <= 691;
        o_index_for_a3 <= 1078;
        o_index_for_a4 <= 1157;
        o_index_for_a5 <= 1637; 
        o_index_for_a6 <= 1733; 
    end
    486: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 440;
        o_index_for_a1 <= 542;
        o_index_for_a2 <= 692;
        o_index_for_a3 <= 1079;
        o_index_for_a4 <= 1158;
        o_index_for_a5 <= 1638; 
        o_index_for_a6 <= 1734; 
    end
    487: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 441;
        o_index_for_a1 <= 543;
        o_index_for_a2 <= 693;
        o_index_for_a3 <= 1080;
        o_index_for_a4 <= 1159;
        o_index_for_a5 <= 1639; 
        o_index_for_a6 <= 1735; 
    end
    488: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 442;
        o_index_for_a1 <= 544;
        o_index_for_a2 <= 694;
        o_index_for_a3 <= 1081;
        o_index_for_a4 <= 1160;
        o_index_for_a5 <= 1640; 
        o_index_for_a6 <= 1736; 
    end
    489: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 443;
        o_index_for_a1 <= 545;
        o_index_for_a2 <= 695;
        o_index_for_a3 <= 1082;
        o_index_for_a4 <= 1161;
        o_index_for_a5 <= 1641; 
        o_index_for_a6 <= 1737; 
    end
    490: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 444;
        o_index_for_a1 <= 546;
        o_index_for_a2 <= 696;
        o_index_for_a3 <= 1083;
        o_index_for_a4 <= 1162;
        o_index_for_a5 <= 1642; 
        o_index_for_a6 <= 1738; 
    end
    491: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 445;
        o_index_for_a1 <= 547;
        o_index_for_a2 <= 697;
        o_index_for_a3 <= 1084;
        o_index_for_a4 <= 1163;
        o_index_for_a5 <= 1643; 
        o_index_for_a6 <= 1739; 
    end
    492: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 446;
        o_index_for_a1 <= 548;
        o_index_for_a2 <= 698;
        o_index_for_a3 <= 1085;
        o_index_for_a4 <= 1164;
        o_index_for_a5 <= 1644; 
        o_index_for_a6 <= 1740; 
    end
    493: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 447;
        o_index_for_a1 <= 549;
        o_index_for_a2 <= 699;
        o_index_for_a3 <= 1086;
        o_index_for_a4 <= 1165;
        o_index_for_a5 <= 1645; 
        o_index_for_a6 <= 1741; 
    end
    494: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 448;
        o_index_for_a1 <= 550;
        o_index_for_a2 <= 700;
        o_index_for_a3 <= 1087;
        o_index_for_a4 <= 1166;
        o_index_for_a5 <= 1646; 
        o_index_for_a6 <= 1742; 
    end
    495: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 449;
        o_index_for_a1 <= 551;
        o_index_for_a2 <= 701;
        o_index_for_a3 <= 1088;
        o_index_for_a4 <= 1167;
        o_index_for_a5 <= 1647; 
        o_index_for_a6 <= 1743; 
    end
    496: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 450;
        o_index_for_a1 <= 552;
        o_index_for_a2 <= 702;
        o_index_for_a3 <= 1089;
        o_index_for_a4 <= 1168;
        o_index_for_a5 <= 1648; 
        o_index_for_a6 <= 1744; 
    end
    497: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 451;
        o_index_for_a1 <= 553;
        o_index_for_a2 <= 703;
        o_index_for_a3 <= 1090;
        o_index_for_a4 <= 1169;
        o_index_for_a5 <= 1649; 
        o_index_for_a6 <= 1745; 
    end
    498: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 452;
        o_index_for_a1 <= 554;
        o_index_for_a2 <= 704;
        o_index_for_a3 <= 1091;
        o_index_for_a4 <= 1170;
        o_index_for_a5 <= 1650; 
        o_index_for_a6 <= 1746; 
    end
    499: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 453;
        o_index_for_a1 <= 555;
        o_index_for_a2 <= 705;
        o_index_for_a3 <= 1092;
        o_index_for_a4 <= 1171;
        o_index_for_a5 <= 1651; 
        o_index_for_a6 <= 1747; 
    end
    500: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 454;
        o_index_for_a1 <= 556;
        o_index_for_a2 <= 706;
        o_index_for_a3 <= 1093;
        o_index_for_a4 <= 1172;
        o_index_for_a5 <= 1652; 
        o_index_for_a6 <= 1748; 
    end
    501: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 455;
        o_index_for_a1 <= 557;
        o_index_for_a2 <= 707;
        o_index_for_a3 <= 1094;
        o_index_for_a4 <= 1173;
        o_index_for_a5 <= 1653; 
        o_index_for_a6 <= 1749; 
    end
    502: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 456;
        o_index_for_a1 <= 558;
        o_index_for_a2 <= 708;
        o_index_for_a3 <= 1095;
        o_index_for_a4 <= 1174;
        o_index_for_a5 <= 1654; 
        o_index_for_a6 <= 1750; 
    end
    503: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 457;
        o_index_for_a1 <= 559;
        o_index_for_a2 <= 709;
        o_index_for_a3 <= 1096;
        o_index_for_a4 <= 1175;
        o_index_for_a5 <= 1655; 
        o_index_for_a6 <= 1751; 
    end
    504: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 458;
        o_index_for_a1 <= 560;
        o_index_for_a2 <= 710;
        o_index_for_a3 <= 1097;
        o_index_for_a4 <= 1176;
        o_index_for_a5 <= 1656; 
        o_index_for_a6 <= 1752; 
    end
    505: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 459;
        o_index_for_a1 <= 561;
        o_index_for_a2 <= 711;
        o_index_for_a3 <= 1098;
        o_index_for_a4 <= 1177;
        o_index_for_a5 <= 1657; 
        o_index_for_a6 <= 1753; 
    end
    506: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 460;
        o_index_for_a1 <= 562;
        o_index_for_a2 <= 712;
        o_index_for_a3 <= 1099;
        o_index_for_a4 <= 1178;
        o_index_for_a5 <= 1658; 
        o_index_for_a6 <= 1754; 
    end
    507: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 461;
        o_index_for_a1 <= 563;
        o_index_for_a2 <= 713;
        o_index_for_a3 <= 1100;
        o_index_for_a4 <= 1179;
        o_index_for_a5 <= 1659; 
        o_index_for_a6 <= 1755; 
    end
    508: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 462;
        o_index_for_a1 <= 564;
        o_index_for_a2 <= 714;
        o_index_for_a3 <= 1101;
        o_index_for_a4 <= 1180;
        o_index_for_a5 <= 1660; 
        o_index_for_a6 <= 1756; 
    end
    509: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 463;
        o_index_for_a1 <= 565;
        o_index_for_a2 <= 715;
        o_index_for_a3 <= 1102;
        o_index_for_a4 <= 1181;
        o_index_for_a5 <= 1661; 
        o_index_for_a6 <= 1757; 
    end
    510: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 464;
        o_index_for_a1 <= 566;
        o_index_for_a2 <= 716;
        o_index_for_a3 <= 1103;
        o_index_for_a4 <= 1182;
        o_index_for_a5 <= 1662; 
        o_index_for_a6 <= 1758; 
    end
    511: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 465;
        o_index_for_a1 <= 567;
        o_index_for_a2 <= 717;
        o_index_for_a3 <= 1104;
        o_index_for_a4 <= 1183;
        o_index_for_a5 <= 1663; 
        o_index_for_a6 <= 1759; 
    end
    512: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 466;
        o_index_for_a1 <= 568;
        o_index_for_a2 <= 718;
        o_index_for_a3 <= 1105;
        o_index_for_a4 <= 1184;
        o_index_for_a5 <= 1664; 
        o_index_for_a6 <= 1760; 
    end
    513: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 467;
        o_index_for_a1 <= 569;
        o_index_for_a2 <= 719;
        o_index_for_a3 <= 1106;
        o_index_for_a4 <= 1185;
        o_index_for_a5 <= 1665; 
        o_index_for_a6 <= 1761; 
    end
    514: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 468;
        o_index_for_a1 <= 570;
        o_index_for_a2 <= 720;
        o_index_for_a3 <= 1107;
        o_index_for_a4 <= 1186;
        o_index_for_a5 <= 1666; 
        o_index_for_a6 <= 1762; 
    end
    515: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 469;
        o_index_for_a1 <= 571;
        o_index_for_a2 <= 721;
        o_index_for_a3 <= 1108;
        o_index_for_a4 <= 1187;
        o_index_for_a5 <= 1667; 
        o_index_for_a6 <= 1763; 
    end
    516: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 470;
        o_index_for_a1 <= 572;
        o_index_for_a2 <= 722;
        o_index_for_a3 <= 1109;
        o_index_for_a4 <= 1188;
        o_index_for_a5 <= 1668; 
        o_index_for_a6 <= 1764; 
    end
    517: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 471;
        o_index_for_a1 <= 573;
        o_index_for_a2 <= 723;
        o_index_for_a3 <= 1110;
        o_index_for_a4 <= 1189;
        o_index_for_a5 <= 1669; 
        o_index_for_a6 <= 1765; 
    end
    518: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 472;
        o_index_for_a1 <= 574;
        o_index_for_a2 <= 724;
        o_index_for_a3 <= 1111;
        o_index_for_a4 <= 1190;
        o_index_for_a5 <= 1670; 
        o_index_for_a6 <= 1766; 
    end
    519: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 473;
        o_index_for_a1 <= 575;
        o_index_for_a2 <= 725;
        o_index_for_a3 <= 1112;
        o_index_for_a4 <= 1191;
        o_index_for_a5 <= 1671; 
        o_index_for_a6 <= 1767; 
    end
    520: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 474;
        o_index_for_a1 <= 480;
        o_index_for_a2 <= 726;
        o_index_for_a3 <= 1113;
        o_index_for_a4 <= 1192;
        o_index_for_a5 <= 1672; 
        o_index_for_a6 <= 1768; 
    end
    521: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 475;
        o_index_for_a1 <= 481;
        o_index_for_a2 <= 727;
        o_index_for_a3 <= 1114;
        o_index_for_a4 <= 1193;
        o_index_for_a5 <= 1673; 
        o_index_for_a6 <= 1769; 
    end
    522: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 476;
        o_index_for_a1 <= 482;
        o_index_for_a2 <= 728;
        o_index_for_a3 <= 1115;
        o_index_for_a4 <= 1194;
        o_index_for_a5 <= 1674; 
        o_index_for_a6 <= 1770; 
    end
    523: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 477;
        o_index_for_a1 <= 483;
        o_index_for_a2 <= 729;
        o_index_for_a3 <= 1116;
        o_index_for_a4 <= 1195;
        o_index_for_a5 <= 1675; 
        o_index_for_a6 <= 1771; 
    end
    524: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 478;
        o_index_for_a1 <= 484;
        o_index_for_a2 <= 730;
        o_index_for_a3 <= 1117;
        o_index_for_a4 <= 1196;
        o_index_for_a5 <= 1676; 
        o_index_for_a6 <= 1772; 
    end
    525: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 479;
        o_index_for_a1 <= 485;
        o_index_for_a2 <= 731;
        o_index_for_a3 <= 1118;
        o_index_for_a4 <= 1197;
        o_index_for_a5 <= 1677; 
        o_index_for_a6 <= 1773; 
    end
    526: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 384;
        o_index_for_a1 <= 486;
        o_index_for_a2 <= 732;
        o_index_for_a3 <= 1119;
        o_index_for_a4 <= 1198;
        o_index_for_a5 <= 1678; 
        o_index_for_a6 <= 1774; 
    end
    527: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 385;
        o_index_for_a1 <= 487;
        o_index_for_a2 <= 733;
        o_index_for_a3 <= 1120;
        o_index_for_a4 <= 1199;
        o_index_for_a5 <= 1679; 
        o_index_for_a6 <= 1775; 
    end
    528: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 386;
        o_index_for_a1 <= 488;
        o_index_for_a2 <= 734;
        o_index_for_a3 <= 1121;
        o_index_for_a4 <= 1200;
        o_index_for_a5 <= 1680; 
        o_index_for_a6 <= 1776; 
    end
    529: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 387;
        o_index_for_a1 <= 489;
        o_index_for_a2 <= 735;
        o_index_for_a3 <= 1122;
        o_index_for_a4 <= 1201;
        o_index_for_a5 <= 1681; 
        o_index_for_a6 <= 1777; 
    end
    530: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 388;
        o_index_for_a1 <= 490;
        o_index_for_a2 <= 736;
        o_index_for_a3 <= 1123;
        o_index_for_a4 <= 1202;
        o_index_for_a5 <= 1682; 
        o_index_for_a6 <= 1778; 
    end
    531: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 389;
        o_index_for_a1 <= 491;
        o_index_for_a2 <= 737;
        o_index_for_a3 <= 1124;
        o_index_for_a4 <= 1203;
        o_index_for_a5 <= 1683; 
        o_index_for_a6 <= 1779; 
    end
    532: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 390;
        o_index_for_a1 <= 492;
        o_index_for_a2 <= 738;
        o_index_for_a3 <= 1125;
        o_index_for_a4 <= 1204;
        o_index_for_a5 <= 1684; 
        o_index_for_a6 <= 1780; 
    end
    533: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 391;
        o_index_for_a1 <= 493;
        o_index_for_a2 <= 739;
        o_index_for_a3 <= 1126;
        o_index_for_a4 <= 1205;
        o_index_for_a5 <= 1685; 
        o_index_for_a6 <= 1781; 
    end
    534: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 392;
        o_index_for_a1 <= 494;
        o_index_for_a2 <= 740;
        o_index_for_a3 <= 1127;
        o_index_for_a4 <= 1206;
        o_index_for_a5 <= 1686; 
        o_index_for_a6 <= 1782; 
    end
    535: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 393;
        o_index_for_a1 <= 495;
        o_index_for_a2 <= 741;
        o_index_for_a3 <= 1128;
        o_index_for_a4 <= 1207;
        o_index_for_a5 <= 1687; 
        o_index_for_a6 <= 1783; 
    end
    536: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 394;
        o_index_for_a1 <= 496;
        o_index_for_a2 <= 742;
        o_index_for_a3 <= 1129;
        o_index_for_a4 <= 1208;
        o_index_for_a5 <= 1688; 
        o_index_for_a6 <= 1784; 
    end
    537: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 395;
        o_index_for_a1 <= 497;
        o_index_for_a2 <= 743;
        o_index_for_a3 <= 1130;
        o_index_for_a4 <= 1209;
        o_index_for_a5 <= 1689; 
        o_index_for_a6 <= 1785; 
    end
    538: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 396;
        o_index_for_a1 <= 498;
        o_index_for_a2 <= 744;
        o_index_for_a3 <= 1131;
        o_index_for_a4 <= 1210;
        o_index_for_a5 <= 1690; 
        o_index_for_a6 <= 1786; 
    end
    539: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 397;
        o_index_for_a1 <= 499;
        o_index_for_a2 <= 745;
        o_index_for_a3 <= 1132;
        o_index_for_a4 <= 1211;
        o_index_for_a5 <= 1691; 
        o_index_for_a6 <= 1787; 
    end
    540: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 398;
        o_index_for_a1 <= 500;
        o_index_for_a2 <= 746;
        o_index_for_a3 <= 1133;
        o_index_for_a4 <= 1212;
        o_index_for_a5 <= 1692; 
        o_index_for_a6 <= 1788; 
    end
    541: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 399;
        o_index_for_a1 <= 501;
        o_index_for_a2 <= 747;
        o_index_for_a3 <= 1134;
        o_index_for_a4 <= 1213;
        o_index_for_a5 <= 1693; 
        o_index_for_a6 <= 1789; 
    end
    542: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 400;
        o_index_for_a1 <= 502;
        o_index_for_a2 <= 748;
        o_index_for_a3 <= 1135;
        o_index_for_a4 <= 1214;
        o_index_for_a5 <= 1694; 
        o_index_for_a6 <= 1790; 
    end
    543: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 401;
        o_index_for_a1 <= 503;
        o_index_for_a2 <= 749;
        o_index_for_a3 <= 1136;
        o_index_for_a4 <= 1215;
        o_index_for_a5 <= 1695; 
        o_index_for_a6 <= 1791; 
    end
    544: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 402;
        o_index_for_a1 <= 504;
        o_index_for_a2 <= 750;
        o_index_for_a3 <= 1137;
        o_index_for_a4 <= 1216;
        o_index_for_a5 <= 1696; 
        o_index_for_a6 <= 1792; 
    end
    545: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 403;
        o_index_for_a1 <= 505;
        o_index_for_a2 <= 751;
        o_index_for_a3 <= 1138;
        o_index_for_a4 <= 1217;
        o_index_for_a5 <= 1697; 
        o_index_for_a6 <= 1793; 
    end
    546: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 404;
        o_index_for_a1 <= 506;
        o_index_for_a2 <= 752;
        o_index_for_a3 <= 1139;
        o_index_for_a4 <= 1218;
        o_index_for_a5 <= 1698; 
        o_index_for_a6 <= 1794; 
    end
    547: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 405;
        o_index_for_a1 <= 507;
        o_index_for_a2 <= 753;
        o_index_for_a3 <= 1140;
        o_index_for_a4 <= 1219;
        o_index_for_a5 <= 1699; 
        o_index_for_a6 <= 1795; 
    end
    548: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 406;
        o_index_for_a1 <= 508;
        o_index_for_a2 <= 754;
        o_index_for_a3 <= 1141;
        o_index_for_a4 <= 1220;
        o_index_for_a5 <= 1700; 
        o_index_for_a6 <= 1796; 
    end
    549: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 407;
        o_index_for_a1 <= 509;
        o_index_for_a2 <= 755;
        o_index_for_a3 <= 1142;
        o_index_for_a4 <= 1221;
        o_index_for_a5 <= 1701; 
        o_index_for_a6 <= 1797; 
    end
    550: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 408;
        o_index_for_a1 <= 510;
        o_index_for_a2 <= 756;
        o_index_for_a3 <= 1143;
        o_index_for_a4 <= 1222;
        o_index_for_a5 <= 1702; 
        o_index_for_a6 <= 1798; 
    end
    551: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 409;
        o_index_for_a1 <= 511;
        o_index_for_a2 <= 757;
        o_index_for_a3 <= 1144;
        o_index_for_a4 <= 1223;
        o_index_for_a5 <= 1703; 
        o_index_for_a6 <= 1799; 
    end
    552: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 410;
        o_index_for_a1 <= 512;
        o_index_for_a2 <= 758;
        o_index_for_a3 <= 1145;
        o_index_for_a4 <= 1224;
        o_index_for_a5 <= 1704; 
        o_index_for_a6 <= 1800; 
    end
    553: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 411;
        o_index_for_a1 <= 513;
        o_index_for_a2 <= 759;
        o_index_for_a3 <= 1146;
        o_index_for_a4 <= 1225;
        o_index_for_a5 <= 1705; 
        o_index_for_a6 <= 1801; 
    end
    554: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 412;
        o_index_for_a1 <= 514;
        o_index_for_a2 <= 760;
        o_index_for_a3 <= 1147;
        o_index_for_a4 <= 1226;
        o_index_for_a5 <= 1706; 
        o_index_for_a6 <= 1802; 
    end
    555: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 413;
        o_index_for_a1 <= 515;
        o_index_for_a2 <= 761;
        o_index_for_a3 <= 1148;
        o_index_for_a4 <= 1227;
        o_index_for_a5 <= 1707; 
        o_index_for_a6 <= 1803; 
    end
    556: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 414;
        o_index_for_a1 <= 516;
        o_index_for_a2 <= 762;
        o_index_for_a3 <= 1149;
        o_index_for_a4 <= 1228;
        o_index_for_a5 <= 1708; 
        o_index_for_a6 <= 1804; 
    end
    557: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 415;
        o_index_for_a1 <= 517;
        o_index_for_a2 <= 763;
        o_index_for_a3 <= 1150;
        o_index_for_a4 <= 1229;
        o_index_for_a5 <= 1709; 
        o_index_for_a6 <= 1805; 
    end
    558: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 416;
        o_index_for_a1 <= 518;
        o_index_for_a2 <= 764;
        o_index_for_a3 <= 1151;
        o_index_for_a4 <= 1230;
        o_index_for_a5 <= 1710; 
        o_index_for_a6 <= 1806; 
    end
    559: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 417;
        o_index_for_a1 <= 519;
        o_index_for_a2 <= 765;
        o_index_for_a3 <= 1056;
        o_index_for_a4 <= 1231;
        o_index_for_a5 <= 1711; 
        o_index_for_a6 <= 1807; 
    end
    560: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 418;
        o_index_for_a1 <= 520;
        o_index_for_a2 <= 766;
        o_index_for_a3 <= 1057;
        o_index_for_a4 <= 1232;
        o_index_for_a5 <= 1712; 
        o_index_for_a6 <= 1808; 
    end
    561: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 419;
        o_index_for_a1 <= 521;
        o_index_for_a2 <= 767;
        o_index_for_a3 <= 1058;
        o_index_for_a4 <= 1233;
        o_index_for_a5 <= 1713; 
        o_index_for_a6 <= 1809; 
    end
    562: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 420;
        o_index_for_a1 <= 522;
        o_index_for_a2 <= 672;
        o_index_for_a3 <= 1059;
        o_index_for_a4 <= 1234;
        o_index_for_a5 <= 1714; 
        o_index_for_a6 <= 1810; 
    end
    563: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 421;
        o_index_for_a1 <= 523;
        o_index_for_a2 <= 673;
        o_index_for_a3 <= 1060;
        o_index_for_a4 <= 1235;
        o_index_for_a5 <= 1715; 
        o_index_for_a6 <= 1811; 
    end
    564: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 422;
        o_index_for_a1 <= 524;
        o_index_for_a2 <= 674;
        o_index_for_a3 <= 1061;
        o_index_for_a4 <= 1236;
        o_index_for_a5 <= 1716; 
        o_index_for_a6 <= 1812; 
    end
    565: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 423;
        o_index_for_a1 <= 525;
        o_index_for_a2 <= 675;
        o_index_for_a3 <= 1062;
        o_index_for_a4 <= 1237;
        o_index_for_a5 <= 1717; 
        o_index_for_a6 <= 1813; 
    end
    566: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 424;
        o_index_for_a1 <= 526;
        o_index_for_a2 <= 676;
        o_index_for_a3 <= 1063;
        o_index_for_a4 <= 1238;
        o_index_for_a5 <= 1718; 
        o_index_for_a6 <= 1814; 
    end
    567: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 425;
        o_index_for_a1 <= 527;
        o_index_for_a2 <= 677;
        o_index_for_a3 <= 1064;
        o_index_for_a4 <= 1239;
        o_index_for_a5 <= 1719; 
        o_index_for_a6 <= 1815; 
    end
    568: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 426;
        o_index_for_a1 <= 528;
        o_index_for_a2 <= 678;
        o_index_for_a3 <= 1065;
        o_index_for_a4 <= 1240;
        o_index_for_a5 <= 1720; 
        o_index_for_a6 <= 1816; 
    end
    569: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 427;
        o_index_for_a1 <= 529;
        o_index_for_a2 <= 679;
        o_index_for_a3 <= 1066;
        o_index_for_a4 <= 1241;
        o_index_for_a5 <= 1721; 
        o_index_for_a6 <= 1817; 
    end
    570: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 428;
        o_index_for_a1 <= 530;
        o_index_for_a2 <= 680;
        o_index_for_a3 <= 1067;
        o_index_for_a4 <= 1242;
        o_index_for_a5 <= 1722; 
        o_index_for_a6 <= 1818; 
    end
    571: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 429;
        o_index_for_a1 <= 531;
        o_index_for_a2 <= 681;
        o_index_for_a3 <= 1068;
        o_index_for_a4 <= 1243;
        o_index_for_a5 <= 1723; 
        o_index_for_a6 <= 1819; 
    end
    572: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 430;
        o_index_for_a1 <= 532;
        o_index_for_a2 <= 682;
        o_index_for_a3 <= 1069;
        o_index_for_a4 <= 1244;
        o_index_for_a5 <= 1724; 
        o_index_for_a6 <= 1820; 
    end
    573: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 431;
        o_index_for_a1 <= 533;
        o_index_for_a2 <= 683;
        o_index_for_a3 <= 1070;
        o_index_for_a4 <= 1245;
        o_index_for_a5 <= 1725; 
        o_index_for_a6 <= 1821; 
    end
    574: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 432;
        o_index_for_a1 <= 534;
        o_index_for_a2 <= 684;
        o_index_for_a3 <= 1071;
        o_index_for_a4 <= 1246;
        o_index_for_a5 <= 1726; 
        o_index_for_a6 <= 1822; 
    end
    575: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 2;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 433;
        o_index_for_a1 <= 535;
        o_index_for_a2 <= 685;
        o_index_for_a3 <= 1072;
        o_index_for_a4 <= 1247;
        o_index_for_a5 <= 1727; 
        o_index_for_a6 <= 1823; 
    end
    576: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 193;
        o_index_for_a1 <= 331;
        o_index_for_a2 <= 946;
        o_index_for_a3 <= 1038;
        o_index_for_a4 <= 1728;
        o_index_for_a5 <= 1824; 
        o_index_for_a6 <= 2304; 
    end
    577: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 194;
        o_index_for_a1 <= 332;
        o_index_for_a2 <= 947;
        o_index_for_a3 <= 1039;
        o_index_for_a4 <= 1729;
        o_index_for_a5 <= 1825; 
        o_index_for_a6 <= 2304; 
    end
    578: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 195;
        o_index_for_a1 <= 333;
        o_index_for_a2 <= 948;
        o_index_for_a3 <= 1040;
        o_index_for_a4 <= 1730;
        o_index_for_a5 <= 1826; 
        o_index_for_a6 <= 2304; 
    end
    579: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 196;
        o_index_for_a1 <= 334;
        o_index_for_a2 <= 949;
        o_index_for_a3 <= 1041;
        o_index_for_a4 <= 1731;
        o_index_for_a5 <= 1827; 
        o_index_for_a6 <= 2304; 
    end
    580: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 197;
        o_index_for_a1 <= 335;
        o_index_for_a2 <= 950;
        o_index_for_a3 <= 1042;
        o_index_for_a4 <= 1732;
        o_index_for_a5 <= 1828; 
        o_index_for_a6 <= 2304; 
    end
    581: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 198;
        o_index_for_a1 <= 336;
        o_index_for_a2 <= 951;
        o_index_for_a3 <= 1043;
        o_index_for_a4 <= 1733;
        o_index_for_a5 <= 1829; 
        o_index_for_a6 <= 2304; 
    end
    582: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 199;
        o_index_for_a1 <= 337;
        o_index_for_a2 <= 952;
        o_index_for_a3 <= 1044;
        o_index_for_a4 <= 1734;
        o_index_for_a5 <= 1830; 
        o_index_for_a6 <= 2304; 
    end
    583: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 200;
        o_index_for_a1 <= 338;
        o_index_for_a2 <= 953;
        o_index_for_a3 <= 1045;
        o_index_for_a4 <= 1735;
        o_index_for_a5 <= 1831; 
        o_index_for_a6 <= 2304; 
    end
    584: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 201;
        o_index_for_a1 <= 339;
        o_index_for_a2 <= 954;
        o_index_for_a3 <= 1046;
        o_index_for_a4 <= 1736;
        o_index_for_a5 <= 1832; 
        o_index_for_a6 <= 2304; 
    end
    585: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 202;
        o_index_for_a1 <= 340;
        o_index_for_a2 <= 955;
        o_index_for_a3 <= 1047;
        o_index_for_a4 <= 1737;
        o_index_for_a5 <= 1833; 
        o_index_for_a6 <= 2304; 
    end
    586: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 203;
        o_index_for_a1 <= 341;
        o_index_for_a2 <= 956;
        o_index_for_a3 <= 1048;
        o_index_for_a4 <= 1738;
        o_index_for_a5 <= 1834; 
        o_index_for_a6 <= 2304; 
    end
    587: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 204;
        o_index_for_a1 <= 342;
        o_index_for_a2 <= 957;
        o_index_for_a3 <= 1049;
        o_index_for_a4 <= 1739;
        o_index_for_a5 <= 1835; 
        o_index_for_a6 <= 2304; 
    end
    588: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 205;
        o_index_for_a1 <= 343;
        o_index_for_a2 <= 958;
        o_index_for_a3 <= 1050;
        o_index_for_a4 <= 1740;
        o_index_for_a5 <= 1836; 
        o_index_for_a6 <= 2304; 
    end
    589: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 206;
        o_index_for_a1 <= 344;
        o_index_for_a2 <= 959;
        o_index_for_a3 <= 1051;
        o_index_for_a4 <= 1741;
        o_index_for_a5 <= 1837; 
        o_index_for_a6 <= 2304; 
    end
    590: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 207;
        o_index_for_a1 <= 345;
        o_index_for_a2 <= 864;
        o_index_for_a3 <= 1052;
        o_index_for_a4 <= 1742;
        o_index_for_a5 <= 1838; 
        o_index_for_a6 <= 2304; 
    end
    591: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 208;
        o_index_for_a1 <= 346;
        o_index_for_a2 <= 865;
        o_index_for_a3 <= 1053;
        o_index_for_a4 <= 1743;
        o_index_for_a5 <= 1839; 
        o_index_for_a6 <= 2304; 
    end
    592: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 209;
        o_index_for_a1 <= 347;
        o_index_for_a2 <= 866;
        o_index_for_a3 <= 1054;
        o_index_for_a4 <= 1744;
        o_index_for_a5 <= 1840; 
        o_index_for_a6 <= 2304; 
    end
    593: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 210;
        o_index_for_a1 <= 348;
        o_index_for_a2 <= 867;
        o_index_for_a3 <= 1055;
        o_index_for_a4 <= 1745;
        o_index_for_a5 <= 1841; 
        o_index_for_a6 <= 2304; 
    end
    594: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 211;
        o_index_for_a1 <= 349;
        o_index_for_a2 <= 868;
        o_index_for_a3 <= 960;
        o_index_for_a4 <= 1746;
        o_index_for_a5 <= 1842; 
        o_index_for_a6 <= 2304; 
    end
    595: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 212;
        o_index_for_a1 <= 350;
        o_index_for_a2 <= 869;
        o_index_for_a3 <= 961;
        o_index_for_a4 <= 1747;
        o_index_for_a5 <= 1843; 
        o_index_for_a6 <= 2304; 
    end
    596: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 213;
        o_index_for_a1 <= 351;
        o_index_for_a2 <= 870;
        o_index_for_a3 <= 962;
        o_index_for_a4 <= 1748;
        o_index_for_a5 <= 1844; 
        o_index_for_a6 <= 2304; 
    end
    597: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 214;
        o_index_for_a1 <= 352;
        o_index_for_a2 <= 871;
        o_index_for_a3 <= 963;
        o_index_for_a4 <= 1749;
        o_index_for_a5 <= 1845; 
        o_index_for_a6 <= 2304; 
    end
    598: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 215;
        o_index_for_a1 <= 353;
        o_index_for_a2 <= 872;
        o_index_for_a3 <= 964;
        o_index_for_a4 <= 1750;
        o_index_for_a5 <= 1846; 
        o_index_for_a6 <= 2304; 
    end
    599: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 216;
        o_index_for_a1 <= 354;
        o_index_for_a2 <= 873;
        o_index_for_a3 <= 965;
        o_index_for_a4 <= 1751;
        o_index_for_a5 <= 1847; 
        o_index_for_a6 <= 2304; 
    end
    600: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 217;
        o_index_for_a1 <= 355;
        o_index_for_a2 <= 874;
        o_index_for_a3 <= 966;
        o_index_for_a4 <= 1752;
        o_index_for_a5 <= 1848; 
        o_index_for_a6 <= 2304; 
    end
    601: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 218;
        o_index_for_a1 <= 356;
        o_index_for_a2 <= 875;
        o_index_for_a3 <= 967;
        o_index_for_a4 <= 1753;
        o_index_for_a5 <= 1849; 
        o_index_for_a6 <= 2304; 
    end
    602: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 219;
        o_index_for_a1 <= 357;
        o_index_for_a2 <= 876;
        o_index_for_a3 <= 968;
        o_index_for_a4 <= 1754;
        o_index_for_a5 <= 1850; 
        o_index_for_a6 <= 2304; 
    end
    603: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 220;
        o_index_for_a1 <= 358;
        o_index_for_a2 <= 877;
        o_index_for_a3 <= 969;
        o_index_for_a4 <= 1755;
        o_index_for_a5 <= 1851; 
        o_index_for_a6 <= 2304; 
    end
    604: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 221;
        o_index_for_a1 <= 359;
        o_index_for_a2 <= 878;
        o_index_for_a3 <= 970;
        o_index_for_a4 <= 1756;
        o_index_for_a5 <= 1852; 
        o_index_for_a6 <= 2304; 
    end
    605: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 222;
        o_index_for_a1 <= 360;
        o_index_for_a2 <= 879;
        o_index_for_a3 <= 971;
        o_index_for_a4 <= 1757;
        o_index_for_a5 <= 1853; 
        o_index_for_a6 <= 2304; 
    end
    606: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 223;
        o_index_for_a1 <= 361;
        o_index_for_a2 <= 880;
        o_index_for_a3 <= 972;
        o_index_for_a4 <= 1758;
        o_index_for_a5 <= 1854; 
        o_index_for_a6 <= 2304; 
    end
    607: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 224;
        o_index_for_a1 <= 362;
        o_index_for_a2 <= 881;
        o_index_for_a3 <= 973;
        o_index_for_a4 <= 1759;
        o_index_for_a5 <= 1855; 
        o_index_for_a6 <= 2304; 
    end
    608: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 225;
        o_index_for_a1 <= 363;
        o_index_for_a2 <= 882;
        o_index_for_a3 <= 974;
        o_index_for_a4 <= 1760;
        o_index_for_a5 <= 1856; 
        o_index_for_a6 <= 2304; 
    end
    609: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 226;
        o_index_for_a1 <= 364;
        o_index_for_a2 <= 883;
        o_index_for_a3 <= 975;
        o_index_for_a4 <= 1761;
        o_index_for_a5 <= 1857; 
        o_index_for_a6 <= 2304; 
    end
    610: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 227;
        o_index_for_a1 <= 365;
        o_index_for_a2 <= 884;
        o_index_for_a3 <= 976;
        o_index_for_a4 <= 1762;
        o_index_for_a5 <= 1858; 
        o_index_for_a6 <= 2304; 
    end
    611: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 228;
        o_index_for_a1 <= 366;
        o_index_for_a2 <= 885;
        o_index_for_a3 <= 977;
        o_index_for_a4 <= 1763;
        o_index_for_a5 <= 1859; 
        o_index_for_a6 <= 2304; 
    end
    612: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 229;
        o_index_for_a1 <= 367;
        o_index_for_a2 <= 886;
        o_index_for_a3 <= 978;
        o_index_for_a4 <= 1764;
        o_index_for_a5 <= 1860; 
        o_index_for_a6 <= 2304; 
    end
    613: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 230;
        o_index_for_a1 <= 368;
        o_index_for_a2 <= 887;
        o_index_for_a3 <= 979;
        o_index_for_a4 <= 1765;
        o_index_for_a5 <= 1861; 
        o_index_for_a6 <= 2304; 
    end
    614: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 231;
        o_index_for_a1 <= 369;
        o_index_for_a2 <= 888;
        o_index_for_a3 <= 980;
        o_index_for_a4 <= 1766;
        o_index_for_a5 <= 1862; 
        o_index_for_a6 <= 2304; 
    end
    615: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 232;
        o_index_for_a1 <= 370;
        o_index_for_a2 <= 889;
        o_index_for_a3 <= 981;
        o_index_for_a4 <= 1767;
        o_index_for_a5 <= 1863; 
        o_index_for_a6 <= 2304; 
    end
    616: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 233;
        o_index_for_a1 <= 371;
        o_index_for_a2 <= 890;
        o_index_for_a3 <= 982;
        o_index_for_a4 <= 1768;
        o_index_for_a5 <= 1864; 
        o_index_for_a6 <= 2304; 
    end
    617: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 234;
        o_index_for_a1 <= 372;
        o_index_for_a2 <= 891;
        o_index_for_a3 <= 983;
        o_index_for_a4 <= 1769;
        o_index_for_a5 <= 1865; 
        o_index_for_a6 <= 2304; 
    end
    618: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 235;
        o_index_for_a1 <= 373;
        o_index_for_a2 <= 892;
        o_index_for_a3 <= 984;
        o_index_for_a4 <= 1770;
        o_index_for_a5 <= 1866; 
        o_index_for_a6 <= 2304; 
    end
    619: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 236;
        o_index_for_a1 <= 374;
        o_index_for_a2 <= 893;
        o_index_for_a3 <= 985;
        o_index_for_a4 <= 1771;
        o_index_for_a5 <= 1867; 
        o_index_for_a6 <= 2304; 
    end
    620: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 237;
        o_index_for_a1 <= 375;
        o_index_for_a2 <= 894;
        o_index_for_a3 <= 986;
        o_index_for_a4 <= 1772;
        o_index_for_a5 <= 1868; 
        o_index_for_a6 <= 2304; 
    end
    621: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 238;
        o_index_for_a1 <= 376;
        o_index_for_a2 <= 895;
        o_index_for_a3 <= 987;
        o_index_for_a4 <= 1773;
        o_index_for_a5 <= 1869; 
        o_index_for_a6 <= 2304; 
    end
    622: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 239;
        o_index_for_a1 <= 377;
        o_index_for_a2 <= 896;
        o_index_for_a3 <= 988;
        o_index_for_a4 <= 1774;
        o_index_for_a5 <= 1870; 
        o_index_for_a6 <= 2304; 
    end
    623: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 240;
        o_index_for_a1 <= 378;
        o_index_for_a2 <= 897;
        o_index_for_a3 <= 989;
        o_index_for_a4 <= 1775;
        o_index_for_a5 <= 1871; 
        o_index_for_a6 <= 2304; 
    end
    624: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 241;
        o_index_for_a1 <= 379;
        o_index_for_a2 <= 898;
        o_index_for_a3 <= 990;
        o_index_for_a4 <= 1776;
        o_index_for_a5 <= 1872; 
        o_index_for_a6 <= 2304; 
    end
    625: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 242;
        o_index_for_a1 <= 380;
        o_index_for_a2 <= 899;
        o_index_for_a3 <= 991;
        o_index_for_a4 <= 1777;
        o_index_for_a5 <= 1873; 
        o_index_for_a6 <= 2304; 
    end
    626: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 243;
        o_index_for_a1 <= 381;
        o_index_for_a2 <= 900;
        o_index_for_a3 <= 992;
        o_index_for_a4 <= 1778;
        o_index_for_a5 <= 1874; 
        o_index_for_a6 <= 2304; 
    end
    627: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 244;
        o_index_for_a1 <= 382;
        o_index_for_a2 <= 901;
        o_index_for_a3 <= 993;
        o_index_for_a4 <= 1779;
        o_index_for_a5 <= 1875; 
        o_index_for_a6 <= 2304; 
    end
    628: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 245;
        o_index_for_a1 <= 383;
        o_index_for_a2 <= 902;
        o_index_for_a3 <= 994;
        o_index_for_a4 <= 1780;
        o_index_for_a5 <= 1876; 
        o_index_for_a6 <= 2304; 
    end
    629: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 246;
        o_index_for_a1 <= 288;
        o_index_for_a2 <= 903;
        o_index_for_a3 <= 995;
        o_index_for_a4 <= 1781;
        o_index_for_a5 <= 1877; 
        o_index_for_a6 <= 2304; 
    end
    630: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 247;
        o_index_for_a1 <= 289;
        o_index_for_a2 <= 904;
        o_index_for_a3 <= 996;
        o_index_for_a4 <= 1782;
        o_index_for_a5 <= 1878; 
        o_index_for_a6 <= 2304; 
    end
    631: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 248;
        o_index_for_a1 <= 290;
        o_index_for_a2 <= 905;
        o_index_for_a3 <= 997;
        o_index_for_a4 <= 1783;
        o_index_for_a5 <= 1879; 
        o_index_for_a6 <= 2304; 
    end
    632: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 249;
        o_index_for_a1 <= 291;
        o_index_for_a2 <= 906;
        o_index_for_a3 <= 998;
        o_index_for_a4 <= 1784;
        o_index_for_a5 <= 1880; 
        o_index_for_a6 <= 2304; 
    end
    633: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 250;
        o_index_for_a1 <= 292;
        o_index_for_a2 <= 907;
        o_index_for_a3 <= 999;
        o_index_for_a4 <= 1785;
        o_index_for_a5 <= 1881; 
        o_index_for_a6 <= 2304; 
    end
    634: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 251;
        o_index_for_a1 <= 293;
        o_index_for_a2 <= 908;
        o_index_for_a3 <= 1000;
        o_index_for_a4 <= 1786;
        o_index_for_a5 <= 1882; 
        o_index_for_a6 <= 2304; 
    end
    635: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 252;
        o_index_for_a1 <= 294;
        o_index_for_a2 <= 909;
        o_index_for_a3 <= 1001;
        o_index_for_a4 <= 1787;
        o_index_for_a5 <= 1883; 
        o_index_for_a6 <= 2304; 
    end
    636: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 253;
        o_index_for_a1 <= 295;
        o_index_for_a2 <= 910;
        o_index_for_a3 <= 1002;
        o_index_for_a4 <= 1788;
        o_index_for_a5 <= 1884; 
        o_index_for_a6 <= 2304; 
    end
    637: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 254;
        o_index_for_a1 <= 296;
        o_index_for_a2 <= 911;
        o_index_for_a3 <= 1003;
        o_index_for_a4 <= 1789;
        o_index_for_a5 <= 1885; 
        o_index_for_a6 <= 2304; 
    end
    638: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 255;
        o_index_for_a1 <= 297;
        o_index_for_a2 <= 912;
        o_index_for_a3 <= 1004;
        o_index_for_a4 <= 1790;
        o_index_for_a5 <= 1886; 
        o_index_for_a6 <= 2304; 
    end
    639: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 256;
        o_index_for_a1 <= 298;
        o_index_for_a2 <= 913;
        o_index_for_a3 <= 1005;
        o_index_for_a4 <= 1791;
        o_index_for_a5 <= 1887; 
        o_index_for_a6 <= 2304; 
    end
    640: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 257;
        o_index_for_a1 <= 299;
        o_index_for_a2 <= 914;
        o_index_for_a3 <= 1006;
        o_index_for_a4 <= 1792;
        o_index_for_a5 <= 1888; 
        o_index_for_a6 <= 2304; 
    end
    641: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 258;
        o_index_for_a1 <= 300;
        o_index_for_a2 <= 915;
        o_index_for_a3 <= 1007;
        o_index_for_a4 <= 1793;
        o_index_for_a5 <= 1889; 
        o_index_for_a6 <= 2304; 
    end
    642: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 259;
        o_index_for_a1 <= 301;
        o_index_for_a2 <= 916;
        o_index_for_a3 <= 1008;
        o_index_for_a4 <= 1794;
        o_index_for_a5 <= 1890; 
        o_index_for_a6 <= 2304; 
    end
    643: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 260;
        o_index_for_a1 <= 302;
        o_index_for_a2 <= 917;
        o_index_for_a3 <= 1009;
        o_index_for_a4 <= 1795;
        o_index_for_a5 <= 1891; 
        o_index_for_a6 <= 2304; 
    end
    644: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 261;
        o_index_for_a1 <= 303;
        o_index_for_a2 <= 918;
        o_index_for_a3 <= 1010;
        o_index_for_a4 <= 1796;
        o_index_for_a5 <= 1892; 
        o_index_for_a6 <= 2304; 
    end
    645: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 262;
        o_index_for_a1 <= 304;
        o_index_for_a2 <= 919;
        o_index_for_a3 <= 1011;
        o_index_for_a4 <= 1797;
        o_index_for_a5 <= 1893; 
        o_index_for_a6 <= 2304; 
    end
    646: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 263;
        o_index_for_a1 <= 305;
        o_index_for_a2 <= 920;
        o_index_for_a3 <= 1012;
        o_index_for_a4 <= 1798;
        o_index_for_a5 <= 1894; 
        o_index_for_a6 <= 2304; 
    end
    647: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 264;
        o_index_for_a1 <= 306;
        o_index_for_a2 <= 921;
        o_index_for_a3 <= 1013;
        o_index_for_a4 <= 1799;
        o_index_for_a5 <= 1895; 
        o_index_for_a6 <= 2304; 
    end
    648: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 265;
        o_index_for_a1 <= 307;
        o_index_for_a2 <= 922;
        o_index_for_a3 <= 1014;
        o_index_for_a4 <= 1800;
        o_index_for_a5 <= 1896; 
        o_index_for_a6 <= 2304; 
    end
    649: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 266;
        o_index_for_a1 <= 308;
        o_index_for_a2 <= 923;
        o_index_for_a3 <= 1015;
        o_index_for_a4 <= 1801;
        o_index_for_a5 <= 1897; 
        o_index_for_a6 <= 2304; 
    end
    650: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 267;
        o_index_for_a1 <= 309;
        o_index_for_a2 <= 924;
        o_index_for_a3 <= 1016;
        o_index_for_a4 <= 1802;
        o_index_for_a5 <= 1898; 
        o_index_for_a6 <= 2304; 
    end
    651: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 268;
        o_index_for_a1 <= 310;
        o_index_for_a2 <= 925;
        o_index_for_a3 <= 1017;
        o_index_for_a4 <= 1803;
        o_index_for_a5 <= 1899; 
        o_index_for_a6 <= 2304; 
    end
    652: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 269;
        o_index_for_a1 <= 311;
        o_index_for_a2 <= 926;
        o_index_for_a3 <= 1018;
        o_index_for_a4 <= 1804;
        o_index_for_a5 <= 1900; 
        o_index_for_a6 <= 2304; 
    end
    653: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 270;
        o_index_for_a1 <= 312;
        o_index_for_a2 <= 927;
        o_index_for_a3 <= 1019;
        o_index_for_a4 <= 1805;
        o_index_for_a5 <= 1901; 
        o_index_for_a6 <= 2304; 
    end
    654: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 271;
        o_index_for_a1 <= 313;
        o_index_for_a2 <= 928;
        o_index_for_a3 <= 1020;
        o_index_for_a4 <= 1806;
        o_index_for_a5 <= 1902; 
        o_index_for_a6 <= 2304; 
    end
    655: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 272;
        o_index_for_a1 <= 314;
        o_index_for_a2 <= 929;
        o_index_for_a3 <= 1021;
        o_index_for_a4 <= 1807;
        o_index_for_a5 <= 1903; 
        o_index_for_a6 <= 2304; 
    end
    656: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 273;
        o_index_for_a1 <= 315;
        o_index_for_a2 <= 930;
        o_index_for_a3 <= 1022;
        o_index_for_a4 <= 1808;
        o_index_for_a5 <= 1904; 
        o_index_for_a6 <= 2304; 
    end
    657: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 274;
        o_index_for_a1 <= 316;
        o_index_for_a2 <= 931;
        o_index_for_a3 <= 1023;
        o_index_for_a4 <= 1809;
        o_index_for_a5 <= 1905; 
        o_index_for_a6 <= 2304; 
    end
    658: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 275;
        o_index_for_a1 <= 317;
        o_index_for_a2 <= 932;
        o_index_for_a3 <= 1024;
        o_index_for_a4 <= 1810;
        o_index_for_a5 <= 1906; 
        o_index_for_a6 <= 2304; 
    end
    659: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 276;
        o_index_for_a1 <= 318;
        o_index_for_a2 <= 933;
        o_index_for_a3 <= 1025;
        o_index_for_a4 <= 1811;
        o_index_for_a5 <= 1907; 
        o_index_for_a6 <= 2304; 
    end
    660: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 277;
        o_index_for_a1 <= 319;
        o_index_for_a2 <= 934;
        o_index_for_a3 <= 1026;
        o_index_for_a4 <= 1812;
        o_index_for_a5 <= 1908; 
        o_index_for_a6 <= 2304; 
    end
    661: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 278;
        o_index_for_a1 <= 320;
        o_index_for_a2 <= 935;
        o_index_for_a3 <= 1027;
        o_index_for_a4 <= 1813;
        o_index_for_a5 <= 1909; 
        o_index_for_a6 <= 2304; 
    end
    662: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 279;
        o_index_for_a1 <= 321;
        o_index_for_a2 <= 936;
        o_index_for_a3 <= 1028;
        o_index_for_a4 <= 1814;
        o_index_for_a5 <= 1910; 
        o_index_for_a6 <= 2304; 
    end
    663: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 280;
        o_index_for_a1 <= 322;
        o_index_for_a2 <= 937;
        o_index_for_a3 <= 1029;
        o_index_for_a4 <= 1815;
        o_index_for_a5 <= 1911; 
        o_index_for_a6 <= 2304; 
    end
    664: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 281;
        o_index_for_a1 <= 323;
        o_index_for_a2 <= 938;
        o_index_for_a3 <= 1030;
        o_index_for_a4 <= 1816;
        o_index_for_a5 <= 1912; 
        o_index_for_a6 <= 2304; 
    end
    665: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 282;
        o_index_for_a1 <= 324;
        o_index_for_a2 <= 939;
        o_index_for_a3 <= 1031;
        o_index_for_a4 <= 1817;
        o_index_for_a5 <= 1913; 
        o_index_for_a6 <= 2304; 
    end
    666: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 283;
        o_index_for_a1 <= 325;
        o_index_for_a2 <= 940;
        o_index_for_a3 <= 1032;
        o_index_for_a4 <= 1818;
        o_index_for_a5 <= 1914; 
        o_index_for_a6 <= 2304; 
    end
    667: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 284;
        o_index_for_a1 <= 326;
        o_index_for_a2 <= 941;
        o_index_for_a3 <= 1033;
        o_index_for_a4 <= 1819;
        o_index_for_a5 <= 1915; 
        o_index_for_a6 <= 2304; 
    end
    668: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 285;
        o_index_for_a1 <= 327;
        o_index_for_a2 <= 942;
        o_index_for_a3 <= 1034;
        o_index_for_a4 <= 1820;
        o_index_for_a5 <= 1916; 
        o_index_for_a6 <= 2304; 
    end
    669: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 286;
        o_index_for_a1 <= 328;
        o_index_for_a2 <= 943;
        o_index_for_a3 <= 1035;
        o_index_for_a4 <= 1821;
        o_index_for_a5 <= 1917; 
        o_index_for_a6 <= 2304; 
    end
    670: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 287;
        o_index_for_a1 <= 329;
        o_index_for_a2 <= 944;
        o_index_for_a3 <= 1036;
        o_index_for_a4 <= 1822;
        o_index_for_a5 <= 1918; 
        o_index_for_a6 <= 2304; 
    end
    671: begin
        o_branch_for_a0 <= 3;
        o_branch_for_a1 <= 1;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 1;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 192;
        o_index_for_a1 <= 330;
        o_index_for_a2 <= 945;
        o_index_for_a3 <= 1037;
        o_index_for_a4 <= 1823;
        o_index_for_a5 <= 1919; 
        o_index_for_a6 <= 2304; 
    end
    672: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 181;
        o_index_for_a1 <= 215;
        o_index_for_a2 <= 670;
        o_index_for_a3 <= 913;
        o_index_for_a4 <= 1824;
        o_index_for_a5 <= 1920; 
        o_index_for_a6 <= 2304; 
    end
    673: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 182;
        o_index_for_a1 <= 216;
        o_index_for_a2 <= 671;
        o_index_for_a3 <= 914;
        o_index_for_a4 <= 1825;
        o_index_for_a5 <= 1921; 
        o_index_for_a6 <= 2304; 
    end
    674: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 183;
        o_index_for_a1 <= 217;
        o_index_for_a2 <= 576;
        o_index_for_a3 <= 915;
        o_index_for_a4 <= 1826;
        o_index_for_a5 <= 1922; 
        o_index_for_a6 <= 2304; 
    end
    675: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 184;
        o_index_for_a1 <= 218;
        o_index_for_a2 <= 577;
        o_index_for_a3 <= 916;
        o_index_for_a4 <= 1827;
        o_index_for_a5 <= 1923; 
        o_index_for_a6 <= 2304; 
    end
    676: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 185;
        o_index_for_a1 <= 219;
        o_index_for_a2 <= 578;
        o_index_for_a3 <= 917;
        o_index_for_a4 <= 1828;
        o_index_for_a5 <= 1924; 
        o_index_for_a6 <= 2304; 
    end
    677: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 186;
        o_index_for_a1 <= 220;
        o_index_for_a2 <= 579;
        o_index_for_a3 <= 918;
        o_index_for_a4 <= 1829;
        o_index_for_a5 <= 1925; 
        o_index_for_a6 <= 2304; 
    end
    678: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 187;
        o_index_for_a1 <= 221;
        o_index_for_a2 <= 580;
        o_index_for_a3 <= 919;
        o_index_for_a4 <= 1830;
        o_index_for_a5 <= 1926; 
        o_index_for_a6 <= 2304; 
    end
    679: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 188;
        o_index_for_a1 <= 222;
        o_index_for_a2 <= 581;
        o_index_for_a3 <= 920;
        o_index_for_a4 <= 1831;
        o_index_for_a5 <= 1927; 
        o_index_for_a6 <= 2304; 
    end
    680: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 189;
        o_index_for_a1 <= 223;
        o_index_for_a2 <= 582;
        o_index_for_a3 <= 921;
        o_index_for_a4 <= 1832;
        o_index_for_a5 <= 1928; 
        o_index_for_a6 <= 2304; 
    end
    681: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 190;
        o_index_for_a1 <= 224;
        o_index_for_a2 <= 583;
        o_index_for_a3 <= 922;
        o_index_for_a4 <= 1833;
        o_index_for_a5 <= 1929; 
        o_index_for_a6 <= 2304; 
    end
    682: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 191;
        o_index_for_a1 <= 225;
        o_index_for_a2 <= 584;
        o_index_for_a3 <= 923;
        o_index_for_a4 <= 1834;
        o_index_for_a5 <= 1930; 
        o_index_for_a6 <= 2304; 
    end
    683: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 96;
        o_index_for_a1 <= 226;
        o_index_for_a2 <= 585;
        o_index_for_a3 <= 924;
        o_index_for_a4 <= 1835;
        o_index_for_a5 <= 1931; 
        o_index_for_a6 <= 2304; 
    end
    684: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 97;
        o_index_for_a1 <= 227;
        o_index_for_a2 <= 586;
        o_index_for_a3 <= 925;
        o_index_for_a4 <= 1836;
        o_index_for_a5 <= 1932; 
        o_index_for_a6 <= 2304; 
    end
    685: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 98;
        o_index_for_a1 <= 228;
        o_index_for_a2 <= 587;
        o_index_for_a3 <= 926;
        o_index_for_a4 <= 1837;
        o_index_for_a5 <= 1933; 
        o_index_for_a6 <= 2304; 
    end
    686: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 99;
        o_index_for_a1 <= 229;
        o_index_for_a2 <= 588;
        o_index_for_a3 <= 927;
        o_index_for_a4 <= 1838;
        o_index_for_a5 <= 1934; 
        o_index_for_a6 <= 2304; 
    end
    687: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 100;
        o_index_for_a1 <= 230;
        o_index_for_a2 <= 589;
        o_index_for_a3 <= 928;
        o_index_for_a4 <= 1839;
        o_index_for_a5 <= 1935; 
        o_index_for_a6 <= 2304; 
    end
    688: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 101;
        o_index_for_a1 <= 231;
        o_index_for_a2 <= 590;
        o_index_for_a3 <= 929;
        o_index_for_a4 <= 1840;
        o_index_for_a5 <= 1936; 
        o_index_for_a6 <= 2304; 
    end
    689: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 102;
        o_index_for_a1 <= 232;
        o_index_for_a2 <= 591;
        o_index_for_a3 <= 930;
        o_index_for_a4 <= 1841;
        o_index_for_a5 <= 1937; 
        o_index_for_a6 <= 2304; 
    end
    690: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 103;
        o_index_for_a1 <= 233;
        o_index_for_a2 <= 592;
        o_index_for_a3 <= 931;
        o_index_for_a4 <= 1842;
        o_index_for_a5 <= 1938; 
        o_index_for_a6 <= 2304; 
    end
    691: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 104;
        o_index_for_a1 <= 234;
        o_index_for_a2 <= 593;
        o_index_for_a3 <= 932;
        o_index_for_a4 <= 1843;
        o_index_for_a5 <= 1939; 
        o_index_for_a6 <= 2304; 
    end
    692: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 105;
        o_index_for_a1 <= 235;
        o_index_for_a2 <= 594;
        o_index_for_a3 <= 933;
        o_index_for_a4 <= 1844;
        o_index_for_a5 <= 1940; 
        o_index_for_a6 <= 2304; 
    end
    693: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 106;
        o_index_for_a1 <= 236;
        o_index_for_a2 <= 595;
        o_index_for_a3 <= 934;
        o_index_for_a4 <= 1845;
        o_index_for_a5 <= 1941; 
        o_index_for_a6 <= 2304; 
    end
    694: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 107;
        o_index_for_a1 <= 237;
        o_index_for_a2 <= 596;
        o_index_for_a3 <= 935;
        o_index_for_a4 <= 1846;
        o_index_for_a5 <= 1942; 
        o_index_for_a6 <= 2304; 
    end
    695: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 108;
        o_index_for_a1 <= 238;
        o_index_for_a2 <= 597;
        o_index_for_a3 <= 936;
        o_index_for_a4 <= 1847;
        o_index_for_a5 <= 1943; 
        o_index_for_a6 <= 2304; 
    end
    696: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 109;
        o_index_for_a1 <= 239;
        o_index_for_a2 <= 598;
        o_index_for_a3 <= 937;
        o_index_for_a4 <= 1848;
        o_index_for_a5 <= 1944; 
        o_index_for_a6 <= 2304; 
    end
    697: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 110;
        o_index_for_a1 <= 240;
        o_index_for_a2 <= 599;
        o_index_for_a3 <= 938;
        o_index_for_a4 <= 1849;
        o_index_for_a5 <= 1945; 
        o_index_for_a6 <= 2304; 
    end
    698: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 111;
        o_index_for_a1 <= 241;
        o_index_for_a2 <= 600;
        o_index_for_a3 <= 939;
        o_index_for_a4 <= 1850;
        o_index_for_a5 <= 1946; 
        o_index_for_a6 <= 2304; 
    end
    699: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 112;
        o_index_for_a1 <= 242;
        o_index_for_a2 <= 601;
        o_index_for_a3 <= 940;
        o_index_for_a4 <= 1851;
        o_index_for_a5 <= 1947; 
        o_index_for_a6 <= 2304; 
    end
    700: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 113;
        o_index_for_a1 <= 243;
        o_index_for_a2 <= 602;
        o_index_for_a3 <= 941;
        o_index_for_a4 <= 1852;
        o_index_for_a5 <= 1948; 
        o_index_for_a6 <= 2304; 
    end
    701: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 114;
        o_index_for_a1 <= 244;
        o_index_for_a2 <= 603;
        o_index_for_a3 <= 942;
        o_index_for_a4 <= 1853;
        o_index_for_a5 <= 1949; 
        o_index_for_a6 <= 2304; 
    end
    702: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 115;
        o_index_for_a1 <= 245;
        o_index_for_a2 <= 604;
        o_index_for_a3 <= 943;
        o_index_for_a4 <= 1854;
        o_index_for_a5 <= 1950; 
        o_index_for_a6 <= 2304; 
    end
    703: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 116;
        o_index_for_a1 <= 246;
        o_index_for_a2 <= 605;
        o_index_for_a3 <= 944;
        o_index_for_a4 <= 1855;
        o_index_for_a5 <= 1951; 
        o_index_for_a6 <= 2304; 
    end
    704: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 117;
        o_index_for_a1 <= 247;
        o_index_for_a2 <= 606;
        o_index_for_a3 <= 945;
        o_index_for_a4 <= 1856;
        o_index_for_a5 <= 1952; 
        o_index_for_a6 <= 2304; 
    end
    705: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 118;
        o_index_for_a1 <= 248;
        o_index_for_a2 <= 607;
        o_index_for_a3 <= 946;
        o_index_for_a4 <= 1857;
        o_index_for_a5 <= 1953; 
        o_index_for_a6 <= 2304; 
    end
    706: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 119;
        o_index_for_a1 <= 249;
        o_index_for_a2 <= 608;
        o_index_for_a3 <= 947;
        o_index_for_a4 <= 1858;
        o_index_for_a5 <= 1954; 
        o_index_for_a6 <= 2304; 
    end
    707: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 120;
        o_index_for_a1 <= 250;
        o_index_for_a2 <= 609;
        o_index_for_a3 <= 948;
        o_index_for_a4 <= 1859;
        o_index_for_a5 <= 1955; 
        o_index_for_a6 <= 2304; 
    end
    708: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 121;
        o_index_for_a1 <= 251;
        o_index_for_a2 <= 610;
        o_index_for_a3 <= 949;
        o_index_for_a4 <= 1860;
        o_index_for_a5 <= 1956; 
        o_index_for_a6 <= 2304; 
    end
    709: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 122;
        o_index_for_a1 <= 252;
        o_index_for_a2 <= 611;
        o_index_for_a3 <= 950;
        o_index_for_a4 <= 1861;
        o_index_for_a5 <= 1957; 
        o_index_for_a6 <= 2304; 
    end
    710: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 123;
        o_index_for_a1 <= 253;
        o_index_for_a2 <= 612;
        o_index_for_a3 <= 951;
        o_index_for_a4 <= 1862;
        o_index_for_a5 <= 1958; 
        o_index_for_a6 <= 2304; 
    end
    711: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 124;
        o_index_for_a1 <= 254;
        o_index_for_a2 <= 613;
        o_index_for_a3 <= 952;
        o_index_for_a4 <= 1863;
        o_index_for_a5 <= 1959; 
        o_index_for_a6 <= 2304; 
    end
    712: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 125;
        o_index_for_a1 <= 255;
        o_index_for_a2 <= 614;
        o_index_for_a3 <= 953;
        o_index_for_a4 <= 1864;
        o_index_for_a5 <= 1960; 
        o_index_for_a6 <= 2304; 
    end
    713: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 126;
        o_index_for_a1 <= 256;
        o_index_for_a2 <= 615;
        o_index_for_a3 <= 954;
        o_index_for_a4 <= 1865;
        o_index_for_a5 <= 1961; 
        o_index_for_a6 <= 2304; 
    end
    714: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 127;
        o_index_for_a1 <= 257;
        o_index_for_a2 <= 616;
        o_index_for_a3 <= 955;
        o_index_for_a4 <= 1866;
        o_index_for_a5 <= 1962; 
        o_index_for_a6 <= 2304; 
    end
    715: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 128;
        o_index_for_a1 <= 258;
        o_index_for_a2 <= 617;
        o_index_for_a3 <= 956;
        o_index_for_a4 <= 1867;
        o_index_for_a5 <= 1963; 
        o_index_for_a6 <= 2304; 
    end
    716: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 129;
        o_index_for_a1 <= 259;
        o_index_for_a2 <= 618;
        o_index_for_a3 <= 957;
        o_index_for_a4 <= 1868;
        o_index_for_a5 <= 1964; 
        o_index_for_a6 <= 2304; 
    end
    717: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 130;
        o_index_for_a1 <= 260;
        o_index_for_a2 <= 619;
        o_index_for_a3 <= 958;
        o_index_for_a4 <= 1869;
        o_index_for_a5 <= 1965; 
        o_index_for_a6 <= 2304; 
    end
    718: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 131;
        o_index_for_a1 <= 261;
        o_index_for_a2 <= 620;
        o_index_for_a3 <= 959;
        o_index_for_a4 <= 1870;
        o_index_for_a5 <= 1966; 
        o_index_for_a6 <= 2304; 
    end
    719: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 132;
        o_index_for_a1 <= 262;
        o_index_for_a2 <= 621;
        o_index_for_a3 <= 864;
        o_index_for_a4 <= 1871;
        o_index_for_a5 <= 1967; 
        o_index_for_a6 <= 2304; 
    end
    720: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 133;
        o_index_for_a1 <= 263;
        o_index_for_a2 <= 622;
        o_index_for_a3 <= 865;
        o_index_for_a4 <= 1872;
        o_index_for_a5 <= 1968; 
        o_index_for_a6 <= 2304; 
    end
    721: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 134;
        o_index_for_a1 <= 264;
        o_index_for_a2 <= 623;
        o_index_for_a3 <= 866;
        o_index_for_a4 <= 1873;
        o_index_for_a5 <= 1969; 
        o_index_for_a6 <= 2304; 
    end
    722: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 135;
        o_index_for_a1 <= 265;
        o_index_for_a2 <= 624;
        o_index_for_a3 <= 867;
        o_index_for_a4 <= 1874;
        o_index_for_a5 <= 1970; 
        o_index_for_a6 <= 2304; 
    end
    723: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 136;
        o_index_for_a1 <= 266;
        o_index_for_a2 <= 625;
        o_index_for_a3 <= 868;
        o_index_for_a4 <= 1875;
        o_index_for_a5 <= 1971; 
        o_index_for_a6 <= 2304; 
    end
    724: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 137;
        o_index_for_a1 <= 267;
        o_index_for_a2 <= 626;
        o_index_for_a3 <= 869;
        o_index_for_a4 <= 1876;
        o_index_for_a5 <= 1972; 
        o_index_for_a6 <= 2304; 
    end
    725: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 138;
        o_index_for_a1 <= 268;
        o_index_for_a2 <= 627;
        o_index_for_a3 <= 870;
        o_index_for_a4 <= 1877;
        o_index_for_a5 <= 1973; 
        o_index_for_a6 <= 2304; 
    end
    726: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 139;
        o_index_for_a1 <= 269;
        o_index_for_a2 <= 628;
        o_index_for_a3 <= 871;
        o_index_for_a4 <= 1878;
        o_index_for_a5 <= 1974; 
        o_index_for_a6 <= 2304; 
    end
    727: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 140;
        o_index_for_a1 <= 270;
        o_index_for_a2 <= 629;
        o_index_for_a3 <= 872;
        o_index_for_a4 <= 1879;
        o_index_for_a5 <= 1975; 
        o_index_for_a6 <= 2304; 
    end
    728: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 141;
        o_index_for_a1 <= 271;
        o_index_for_a2 <= 630;
        o_index_for_a3 <= 873;
        o_index_for_a4 <= 1880;
        o_index_for_a5 <= 1976; 
        o_index_for_a6 <= 2304; 
    end
    729: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 142;
        o_index_for_a1 <= 272;
        o_index_for_a2 <= 631;
        o_index_for_a3 <= 874;
        o_index_for_a4 <= 1881;
        o_index_for_a5 <= 1977; 
        o_index_for_a6 <= 2304; 
    end
    730: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 143;
        o_index_for_a1 <= 273;
        o_index_for_a2 <= 632;
        o_index_for_a3 <= 875;
        o_index_for_a4 <= 1882;
        o_index_for_a5 <= 1978; 
        o_index_for_a6 <= 2304; 
    end
    731: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 144;
        o_index_for_a1 <= 274;
        o_index_for_a2 <= 633;
        o_index_for_a3 <= 876;
        o_index_for_a4 <= 1883;
        o_index_for_a5 <= 1979; 
        o_index_for_a6 <= 2304; 
    end
    732: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 145;
        o_index_for_a1 <= 275;
        o_index_for_a2 <= 634;
        o_index_for_a3 <= 877;
        o_index_for_a4 <= 1884;
        o_index_for_a5 <= 1980; 
        o_index_for_a6 <= 2304; 
    end
    733: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 146;
        o_index_for_a1 <= 276;
        o_index_for_a2 <= 635;
        o_index_for_a3 <= 878;
        o_index_for_a4 <= 1885;
        o_index_for_a5 <= 1981; 
        o_index_for_a6 <= 2304; 
    end
    734: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 147;
        o_index_for_a1 <= 277;
        o_index_for_a2 <= 636;
        o_index_for_a3 <= 879;
        o_index_for_a4 <= 1886;
        o_index_for_a5 <= 1982; 
        o_index_for_a6 <= 2304; 
    end
    735: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 148;
        o_index_for_a1 <= 278;
        o_index_for_a2 <= 637;
        o_index_for_a3 <= 880;
        o_index_for_a4 <= 1887;
        o_index_for_a5 <= 1983; 
        o_index_for_a6 <= 2304; 
    end
    736: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 149;
        o_index_for_a1 <= 279;
        o_index_for_a2 <= 638;
        o_index_for_a3 <= 881;
        o_index_for_a4 <= 1888;
        o_index_for_a5 <= 1984; 
        o_index_for_a6 <= 2304; 
    end
    737: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 150;
        o_index_for_a1 <= 280;
        o_index_for_a2 <= 639;
        o_index_for_a3 <= 882;
        o_index_for_a4 <= 1889;
        o_index_for_a5 <= 1985; 
        o_index_for_a6 <= 2304; 
    end
    738: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 151;
        o_index_for_a1 <= 281;
        o_index_for_a2 <= 640;
        o_index_for_a3 <= 883;
        o_index_for_a4 <= 1890;
        o_index_for_a5 <= 1986; 
        o_index_for_a6 <= 2304; 
    end
    739: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 152;
        o_index_for_a1 <= 282;
        o_index_for_a2 <= 641;
        o_index_for_a3 <= 884;
        o_index_for_a4 <= 1891;
        o_index_for_a5 <= 1987; 
        o_index_for_a6 <= 2304; 
    end
    740: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 153;
        o_index_for_a1 <= 283;
        o_index_for_a2 <= 642;
        o_index_for_a3 <= 885;
        o_index_for_a4 <= 1892;
        o_index_for_a5 <= 1988; 
        o_index_for_a6 <= 2304; 
    end
    741: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 154;
        o_index_for_a1 <= 284;
        o_index_for_a2 <= 643;
        o_index_for_a3 <= 886;
        o_index_for_a4 <= 1893;
        o_index_for_a5 <= 1989; 
        o_index_for_a6 <= 2304; 
    end
    742: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 155;
        o_index_for_a1 <= 285;
        o_index_for_a2 <= 644;
        o_index_for_a3 <= 887;
        o_index_for_a4 <= 1894;
        o_index_for_a5 <= 1990; 
        o_index_for_a6 <= 2304; 
    end
    743: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 156;
        o_index_for_a1 <= 286;
        o_index_for_a2 <= 645;
        o_index_for_a3 <= 888;
        o_index_for_a4 <= 1895;
        o_index_for_a5 <= 1991; 
        o_index_for_a6 <= 2304; 
    end
    744: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 157;
        o_index_for_a1 <= 287;
        o_index_for_a2 <= 646;
        o_index_for_a3 <= 889;
        o_index_for_a4 <= 1896;
        o_index_for_a5 <= 1992; 
        o_index_for_a6 <= 2304; 
    end
    745: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 158;
        o_index_for_a1 <= 192;
        o_index_for_a2 <= 647;
        o_index_for_a3 <= 890;
        o_index_for_a4 <= 1897;
        o_index_for_a5 <= 1993; 
        o_index_for_a6 <= 2304; 
    end
    746: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 159;
        o_index_for_a1 <= 193;
        o_index_for_a2 <= 648;
        o_index_for_a3 <= 891;
        o_index_for_a4 <= 1898;
        o_index_for_a5 <= 1994; 
        o_index_for_a6 <= 2304; 
    end
    747: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 160;
        o_index_for_a1 <= 194;
        o_index_for_a2 <= 649;
        o_index_for_a3 <= 892;
        o_index_for_a4 <= 1899;
        o_index_for_a5 <= 1995; 
        o_index_for_a6 <= 2304; 
    end
    748: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 161;
        o_index_for_a1 <= 195;
        o_index_for_a2 <= 650;
        o_index_for_a3 <= 893;
        o_index_for_a4 <= 1900;
        o_index_for_a5 <= 1996; 
        o_index_for_a6 <= 2304; 
    end
    749: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 162;
        o_index_for_a1 <= 196;
        o_index_for_a2 <= 651;
        o_index_for_a3 <= 894;
        o_index_for_a4 <= 1901;
        o_index_for_a5 <= 1997; 
        o_index_for_a6 <= 2304; 
    end
    750: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 163;
        o_index_for_a1 <= 197;
        o_index_for_a2 <= 652;
        o_index_for_a3 <= 895;
        o_index_for_a4 <= 1902;
        o_index_for_a5 <= 1998; 
        o_index_for_a6 <= 2304; 
    end
    751: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 164;
        o_index_for_a1 <= 198;
        o_index_for_a2 <= 653;
        o_index_for_a3 <= 896;
        o_index_for_a4 <= 1903;
        o_index_for_a5 <= 1999; 
        o_index_for_a6 <= 2304; 
    end
    752: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 165;
        o_index_for_a1 <= 199;
        o_index_for_a2 <= 654;
        o_index_for_a3 <= 897;
        o_index_for_a4 <= 1904;
        o_index_for_a5 <= 2000; 
        o_index_for_a6 <= 2304; 
    end
    753: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 166;
        o_index_for_a1 <= 200;
        o_index_for_a2 <= 655;
        o_index_for_a3 <= 898;
        o_index_for_a4 <= 1905;
        o_index_for_a5 <= 2001; 
        o_index_for_a6 <= 2304; 
    end
    754: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 167;
        o_index_for_a1 <= 201;
        o_index_for_a2 <= 656;
        o_index_for_a3 <= 899;
        o_index_for_a4 <= 1906;
        o_index_for_a5 <= 2002; 
        o_index_for_a6 <= 2304; 
    end
    755: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 168;
        o_index_for_a1 <= 202;
        o_index_for_a2 <= 657;
        o_index_for_a3 <= 900;
        o_index_for_a4 <= 1907;
        o_index_for_a5 <= 2003; 
        o_index_for_a6 <= 2304; 
    end
    756: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 169;
        o_index_for_a1 <= 203;
        o_index_for_a2 <= 658;
        o_index_for_a3 <= 901;
        o_index_for_a4 <= 1908;
        o_index_for_a5 <= 2004; 
        o_index_for_a6 <= 2304; 
    end
    757: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 170;
        o_index_for_a1 <= 204;
        o_index_for_a2 <= 659;
        o_index_for_a3 <= 902;
        o_index_for_a4 <= 1909;
        o_index_for_a5 <= 2005; 
        o_index_for_a6 <= 2304; 
    end
    758: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 171;
        o_index_for_a1 <= 205;
        o_index_for_a2 <= 660;
        o_index_for_a3 <= 903;
        o_index_for_a4 <= 1910;
        o_index_for_a5 <= 2006; 
        o_index_for_a6 <= 2304; 
    end
    759: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 172;
        o_index_for_a1 <= 206;
        o_index_for_a2 <= 661;
        o_index_for_a3 <= 904;
        o_index_for_a4 <= 1911;
        o_index_for_a5 <= 2007; 
        o_index_for_a6 <= 2304; 
    end
    760: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 173;
        o_index_for_a1 <= 207;
        o_index_for_a2 <= 662;
        o_index_for_a3 <= 905;
        o_index_for_a4 <= 1912;
        o_index_for_a5 <= 2008; 
        o_index_for_a6 <= 2304; 
    end
    761: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 174;
        o_index_for_a1 <= 208;
        o_index_for_a2 <= 663;
        o_index_for_a3 <= 906;
        o_index_for_a4 <= 1913;
        o_index_for_a5 <= 2009; 
        o_index_for_a6 <= 2304; 
    end
    762: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 175;
        o_index_for_a1 <= 209;
        o_index_for_a2 <= 664;
        o_index_for_a3 <= 907;
        o_index_for_a4 <= 1914;
        o_index_for_a5 <= 2010; 
        o_index_for_a6 <= 2304; 
    end
    763: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 176;
        o_index_for_a1 <= 210;
        o_index_for_a2 <= 665;
        o_index_for_a3 <= 908;
        o_index_for_a4 <= 1915;
        o_index_for_a5 <= 2011; 
        o_index_for_a6 <= 2304; 
    end
    764: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 177;
        o_index_for_a1 <= 211;
        o_index_for_a2 <= 666;
        o_index_for_a3 <= 909;
        o_index_for_a4 <= 1916;
        o_index_for_a5 <= 2012; 
        o_index_for_a6 <= 2304; 
    end
    765: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 178;
        o_index_for_a1 <= 212;
        o_index_for_a2 <= 667;
        o_index_for_a3 <= 910;
        o_index_for_a4 <= 1917;
        o_index_for_a5 <= 2013; 
        o_index_for_a6 <= 2304; 
    end
    766: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 179;
        o_index_for_a1 <= 213;
        o_index_for_a2 <= 668;
        o_index_for_a3 <= 911;
        o_index_for_a4 <= 1918;
        o_index_for_a5 <= 2014; 
        o_index_for_a6 <= 2304; 
    end
    767: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 180;
        o_index_for_a1 <= 214;
        o_index_for_a2 <= 669;
        o_index_for_a3 <= 912;
        o_index_for_a4 <= 1919;
        o_index_for_a5 <= 2015; 
        o_index_for_a6 <= 2304; 
    end
    768: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 84;
        o_index_for_a1 <= 397;
        o_index_for_a2 <= 552;
        o_index_for_a3 <= 725;
        o_index_for_a4 <= 1101;
        o_index_for_a5 <= 1920; 
        o_index_for_a6 <= 2016; 
    end
    769: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 85;
        o_index_for_a1 <= 398;
        o_index_for_a2 <= 553;
        o_index_for_a3 <= 726;
        o_index_for_a4 <= 1102;
        o_index_for_a5 <= 1921; 
        o_index_for_a6 <= 2017; 
    end
    770: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 86;
        o_index_for_a1 <= 399;
        o_index_for_a2 <= 554;
        o_index_for_a3 <= 727;
        o_index_for_a4 <= 1103;
        o_index_for_a5 <= 1922; 
        o_index_for_a6 <= 2018; 
    end
    771: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 87;
        o_index_for_a1 <= 400;
        o_index_for_a2 <= 555;
        o_index_for_a3 <= 728;
        o_index_for_a4 <= 1104;
        o_index_for_a5 <= 1923; 
        o_index_for_a6 <= 2019; 
    end
    772: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 88;
        o_index_for_a1 <= 401;
        o_index_for_a2 <= 556;
        o_index_for_a3 <= 729;
        o_index_for_a4 <= 1105;
        o_index_for_a5 <= 1924; 
        o_index_for_a6 <= 2020; 
    end
    773: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 89;
        o_index_for_a1 <= 402;
        o_index_for_a2 <= 557;
        o_index_for_a3 <= 730;
        o_index_for_a4 <= 1106;
        o_index_for_a5 <= 1925; 
        o_index_for_a6 <= 2021; 
    end
    774: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 90;
        o_index_for_a1 <= 403;
        o_index_for_a2 <= 558;
        o_index_for_a3 <= 731;
        o_index_for_a4 <= 1107;
        o_index_for_a5 <= 1926; 
        o_index_for_a6 <= 2022; 
    end
    775: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 91;
        o_index_for_a1 <= 404;
        o_index_for_a2 <= 559;
        o_index_for_a3 <= 732;
        o_index_for_a4 <= 1108;
        o_index_for_a5 <= 1927; 
        o_index_for_a6 <= 2023; 
    end
    776: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 92;
        o_index_for_a1 <= 405;
        o_index_for_a2 <= 560;
        o_index_for_a3 <= 733;
        o_index_for_a4 <= 1109;
        o_index_for_a5 <= 1928; 
        o_index_for_a6 <= 2024; 
    end
    777: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 93;
        o_index_for_a1 <= 406;
        o_index_for_a2 <= 561;
        o_index_for_a3 <= 734;
        o_index_for_a4 <= 1110;
        o_index_for_a5 <= 1929; 
        o_index_for_a6 <= 2025; 
    end
    778: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 94;
        o_index_for_a1 <= 407;
        o_index_for_a2 <= 562;
        o_index_for_a3 <= 735;
        o_index_for_a4 <= 1111;
        o_index_for_a5 <= 1930; 
        o_index_for_a6 <= 2026; 
    end
    779: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 95;
        o_index_for_a1 <= 408;
        o_index_for_a2 <= 563;
        o_index_for_a3 <= 736;
        o_index_for_a4 <= 1112;
        o_index_for_a5 <= 1931; 
        o_index_for_a6 <= 2027; 
    end
    780: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 0;
        o_index_for_a1 <= 409;
        o_index_for_a2 <= 564;
        o_index_for_a3 <= 737;
        o_index_for_a4 <= 1113;
        o_index_for_a5 <= 1932; 
        o_index_for_a6 <= 2028; 
    end
    781: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 1;
        o_index_for_a1 <= 410;
        o_index_for_a2 <= 565;
        o_index_for_a3 <= 738;
        o_index_for_a4 <= 1114;
        o_index_for_a5 <= 1933; 
        o_index_for_a6 <= 2029; 
    end
    782: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 2;
        o_index_for_a1 <= 411;
        o_index_for_a2 <= 566;
        o_index_for_a3 <= 739;
        o_index_for_a4 <= 1115;
        o_index_for_a5 <= 1934; 
        o_index_for_a6 <= 2030; 
    end
    783: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 3;
        o_index_for_a1 <= 412;
        o_index_for_a2 <= 567;
        o_index_for_a3 <= 740;
        o_index_for_a4 <= 1116;
        o_index_for_a5 <= 1935; 
        o_index_for_a6 <= 2031; 
    end
    784: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 4;
        o_index_for_a1 <= 413;
        o_index_for_a2 <= 568;
        o_index_for_a3 <= 741;
        o_index_for_a4 <= 1117;
        o_index_for_a5 <= 1936; 
        o_index_for_a6 <= 2032; 
    end
    785: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 5;
        o_index_for_a1 <= 414;
        o_index_for_a2 <= 569;
        o_index_for_a3 <= 742;
        o_index_for_a4 <= 1118;
        o_index_for_a5 <= 1937; 
        o_index_for_a6 <= 2033; 
    end
    786: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 6;
        o_index_for_a1 <= 415;
        o_index_for_a2 <= 570;
        o_index_for_a3 <= 743;
        o_index_for_a4 <= 1119;
        o_index_for_a5 <= 1938; 
        o_index_for_a6 <= 2034; 
    end
    787: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 7;
        o_index_for_a1 <= 416;
        o_index_for_a2 <= 571;
        o_index_for_a3 <= 744;
        o_index_for_a4 <= 1120;
        o_index_for_a5 <= 1939; 
        o_index_for_a6 <= 2035; 
    end
    788: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 8;
        o_index_for_a1 <= 417;
        o_index_for_a2 <= 572;
        o_index_for_a3 <= 745;
        o_index_for_a4 <= 1121;
        o_index_for_a5 <= 1940; 
        o_index_for_a6 <= 2036; 
    end
    789: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 9;
        o_index_for_a1 <= 418;
        o_index_for_a2 <= 573;
        o_index_for_a3 <= 746;
        o_index_for_a4 <= 1122;
        o_index_for_a5 <= 1941; 
        o_index_for_a6 <= 2037; 
    end
    790: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 10;
        o_index_for_a1 <= 419;
        o_index_for_a2 <= 574;
        o_index_for_a3 <= 747;
        o_index_for_a4 <= 1123;
        o_index_for_a5 <= 1942; 
        o_index_for_a6 <= 2038; 
    end
    791: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 11;
        o_index_for_a1 <= 420;
        o_index_for_a2 <= 575;
        o_index_for_a3 <= 748;
        o_index_for_a4 <= 1124;
        o_index_for_a5 <= 1943; 
        o_index_for_a6 <= 2039; 
    end
    792: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 12;
        o_index_for_a1 <= 421;
        o_index_for_a2 <= 480;
        o_index_for_a3 <= 749;
        o_index_for_a4 <= 1125;
        o_index_for_a5 <= 1944; 
        o_index_for_a6 <= 2040; 
    end
    793: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 13;
        o_index_for_a1 <= 422;
        o_index_for_a2 <= 481;
        o_index_for_a3 <= 750;
        o_index_for_a4 <= 1126;
        o_index_for_a5 <= 1945; 
        o_index_for_a6 <= 2041; 
    end
    794: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 14;
        o_index_for_a1 <= 423;
        o_index_for_a2 <= 482;
        o_index_for_a3 <= 751;
        o_index_for_a4 <= 1127;
        o_index_for_a5 <= 1946; 
        o_index_for_a6 <= 2042; 
    end
    795: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 15;
        o_index_for_a1 <= 424;
        o_index_for_a2 <= 483;
        o_index_for_a3 <= 752;
        o_index_for_a4 <= 1128;
        o_index_for_a5 <= 1947; 
        o_index_for_a6 <= 2043; 
    end
    796: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 16;
        o_index_for_a1 <= 425;
        o_index_for_a2 <= 484;
        o_index_for_a3 <= 753;
        o_index_for_a4 <= 1129;
        o_index_for_a5 <= 1948; 
        o_index_for_a6 <= 2044; 
    end
    797: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 17;
        o_index_for_a1 <= 426;
        o_index_for_a2 <= 485;
        o_index_for_a3 <= 754;
        o_index_for_a4 <= 1130;
        o_index_for_a5 <= 1949; 
        o_index_for_a6 <= 2045; 
    end
    798: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 18;
        o_index_for_a1 <= 427;
        o_index_for_a2 <= 486;
        o_index_for_a3 <= 755;
        o_index_for_a4 <= 1131;
        o_index_for_a5 <= 1950; 
        o_index_for_a6 <= 2046; 
    end
    799: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 19;
        o_index_for_a1 <= 428;
        o_index_for_a2 <= 487;
        o_index_for_a3 <= 756;
        o_index_for_a4 <= 1132;
        o_index_for_a5 <= 1951; 
        o_index_for_a6 <= 2047; 
    end
    800: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 20;
        o_index_for_a1 <= 429;
        o_index_for_a2 <= 488;
        o_index_for_a3 <= 757;
        o_index_for_a4 <= 1133;
        o_index_for_a5 <= 1952; 
        o_index_for_a6 <= 2048; 
    end
    801: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 21;
        o_index_for_a1 <= 430;
        o_index_for_a2 <= 489;
        o_index_for_a3 <= 758;
        o_index_for_a4 <= 1134;
        o_index_for_a5 <= 1953; 
        o_index_for_a6 <= 2049; 
    end
    802: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 22;
        o_index_for_a1 <= 431;
        o_index_for_a2 <= 490;
        o_index_for_a3 <= 759;
        o_index_for_a4 <= 1135;
        o_index_for_a5 <= 1954; 
        o_index_for_a6 <= 2050; 
    end
    803: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 23;
        o_index_for_a1 <= 432;
        o_index_for_a2 <= 491;
        o_index_for_a3 <= 760;
        o_index_for_a4 <= 1136;
        o_index_for_a5 <= 1955; 
        o_index_for_a6 <= 2051; 
    end
    804: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 24;
        o_index_for_a1 <= 433;
        o_index_for_a2 <= 492;
        o_index_for_a3 <= 761;
        o_index_for_a4 <= 1137;
        o_index_for_a5 <= 1956; 
        o_index_for_a6 <= 2052; 
    end
    805: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 25;
        o_index_for_a1 <= 434;
        o_index_for_a2 <= 493;
        o_index_for_a3 <= 762;
        o_index_for_a4 <= 1138;
        o_index_for_a5 <= 1957; 
        o_index_for_a6 <= 2053; 
    end
    806: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 26;
        o_index_for_a1 <= 435;
        o_index_for_a2 <= 494;
        o_index_for_a3 <= 763;
        o_index_for_a4 <= 1139;
        o_index_for_a5 <= 1958; 
        o_index_for_a6 <= 2054; 
    end
    807: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 27;
        o_index_for_a1 <= 436;
        o_index_for_a2 <= 495;
        o_index_for_a3 <= 764;
        o_index_for_a4 <= 1140;
        o_index_for_a5 <= 1959; 
        o_index_for_a6 <= 2055; 
    end
    808: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 28;
        o_index_for_a1 <= 437;
        o_index_for_a2 <= 496;
        o_index_for_a3 <= 765;
        o_index_for_a4 <= 1141;
        o_index_for_a5 <= 1960; 
        o_index_for_a6 <= 2056; 
    end
    809: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 29;
        o_index_for_a1 <= 438;
        o_index_for_a2 <= 497;
        o_index_for_a3 <= 766;
        o_index_for_a4 <= 1142;
        o_index_for_a5 <= 1961; 
        o_index_for_a6 <= 2057; 
    end
    810: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 30;
        o_index_for_a1 <= 439;
        o_index_for_a2 <= 498;
        o_index_for_a3 <= 767;
        o_index_for_a4 <= 1143;
        o_index_for_a5 <= 1962; 
        o_index_for_a6 <= 2058; 
    end
    811: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 31;
        o_index_for_a1 <= 440;
        o_index_for_a2 <= 499;
        o_index_for_a3 <= 672;
        o_index_for_a4 <= 1144;
        o_index_for_a5 <= 1963; 
        o_index_for_a6 <= 2059; 
    end
    812: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 32;
        o_index_for_a1 <= 441;
        o_index_for_a2 <= 500;
        o_index_for_a3 <= 673;
        o_index_for_a4 <= 1145;
        o_index_for_a5 <= 1964; 
        o_index_for_a6 <= 2060; 
    end
    813: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 33;
        o_index_for_a1 <= 442;
        o_index_for_a2 <= 501;
        o_index_for_a3 <= 674;
        o_index_for_a4 <= 1146;
        o_index_for_a5 <= 1965; 
        o_index_for_a6 <= 2061; 
    end
    814: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 34;
        o_index_for_a1 <= 443;
        o_index_for_a2 <= 502;
        o_index_for_a3 <= 675;
        o_index_for_a4 <= 1147;
        o_index_for_a5 <= 1966; 
        o_index_for_a6 <= 2062; 
    end
    815: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 35;
        o_index_for_a1 <= 444;
        o_index_for_a2 <= 503;
        o_index_for_a3 <= 676;
        o_index_for_a4 <= 1148;
        o_index_for_a5 <= 1967; 
        o_index_for_a6 <= 2063; 
    end
    816: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 36;
        o_index_for_a1 <= 445;
        o_index_for_a2 <= 504;
        o_index_for_a3 <= 677;
        o_index_for_a4 <= 1149;
        o_index_for_a5 <= 1968; 
        o_index_for_a6 <= 2064; 
    end
    817: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 37;
        o_index_for_a1 <= 446;
        o_index_for_a2 <= 505;
        o_index_for_a3 <= 678;
        o_index_for_a4 <= 1150;
        o_index_for_a5 <= 1969; 
        o_index_for_a6 <= 2065; 
    end
    818: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 38;
        o_index_for_a1 <= 447;
        o_index_for_a2 <= 506;
        o_index_for_a3 <= 679;
        o_index_for_a4 <= 1151;
        o_index_for_a5 <= 1970; 
        o_index_for_a6 <= 2066; 
    end
    819: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 39;
        o_index_for_a1 <= 448;
        o_index_for_a2 <= 507;
        o_index_for_a3 <= 680;
        o_index_for_a4 <= 1056;
        o_index_for_a5 <= 1971; 
        o_index_for_a6 <= 2067; 
    end
    820: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 40;
        o_index_for_a1 <= 449;
        o_index_for_a2 <= 508;
        o_index_for_a3 <= 681;
        o_index_for_a4 <= 1057;
        o_index_for_a5 <= 1972; 
        o_index_for_a6 <= 2068; 
    end
    821: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 41;
        o_index_for_a1 <= 450;
        o_index_for_a2 <= 509;
        o_index_for_a3 <= 682;
        o_index_for_a4 <= 1058;
        o_index_for_a5 <= 1973; 
        o_index_for_a6 <= 2069; 
    end
    822: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 42;
        o_index_for_a1 <= 451;
        o_index_for_a2 <= 510;
        o_index_for_a3 <= 683;
        o_index_for_a4 <= 1059;
        o_index_for_a5 <= 1974; 
        o_index_for_a6 <= 2070; 
    end
    823: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 43;
        o_index_for_a1 <= 452;
        o_index_for_a2 <= 511;
        o_index_for_a3 <= 684;
        o_index_for_a4 <= 1060;
        o_index_for_a5 <= 1975; 
        o_index_for_a6 <= 2071; 
    end
    824: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 44;
        o_index_for_a1 <= 453;
        o_index_for_a2 <= 512;
        o_index_for_a3 <= 685;
        o_index_for_a4 <= 1061;
        o_index_for_a5 <= 1976; 
        o_index_for_a6 <= 2072; 
    end
    825: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 45;
        o_index_for_a1 <= 454;
        o_index_for_a2 <= 513;
        o_index_for_a3 <= 686;
        o_index_for_a4 <= 1062;
        o_index_for_a5 <= 1977; 
        o_index_for_a6 <= 2073; 
    end
    826: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 46;
        o_index_for_a1 <= 455;
        o_index_for_a2 <= 514;
        o_index_for_a3 <= 687;
        o_index_for_a4 <= 1063;
        o_index_for_a5 <= 1978; 
        o_index_for_a6 <= 2074; 
    end
    827: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 47;
        o_index_for_a1 <= 456;
        o_index_for_a2 <= 515;
        o_index_for_a3 <= 688;
        o_index_for_a4 <= 1064;
        o_index_for_a5 <= 1979; 
        o_index_for_a6 <= 2075; 
    end
    828: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 48;
        o_index_for_a1 <= 457;
        o_index_for_a2 <= 516;
        o_index_for_a3 <= 689;
        o_index_for_a4 <= 1065;
        o_index_for_a5 <= 1980; 
        o_index_for_a6 <= 2076; 
    end
    829: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 49;
        o_index_for_a1 <= 458;
        o_index_for_a2 <= 517;
        o_index_for_a3 <= 690;
        o_index_for_a4 <= 1066;
        o_index_for_a5 <= 1981; 
        o_index_for_a6 <= 2077; 
    end
    830: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 50;
        o_index_for_a1 <= 459;
        o_index_for_a2 <= 518;
        o_index_for_a3 <= 691;
        o_index_for_a4 <= 1067;
        o_index_for_a5 <= 1982; 
        o_index_for_a6 <= 2078; 
    end
    831: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 51;
        o_index_for_a1 <= 460;
        o_index_for_a2 <= 519;
        o_index_for_a3 <= 692;
        o_index_for_a4 <= 1068;
        o_index_for_a5 <= 1983; 
        o_index_for_a6 <= 2079; 
    end
    832: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 52;
        o_index_for_a1 <= 461;
        o_index_for_a2 <= 520;
        o_index_for_a3 <= 693;
        o_index_for_a4 <= 1069;
        o_index_for_a5 <= 1984; 
        o_index_for_a6 <= 2080; 
    end
    833: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 53;
        o_index_for_a1 <= 462;
        o_index_for_a2 <= 521;
        o_index_for_a3 <= 694;
        o_index_for_a4 <= 1070;
        o_index_for_a5 <= 1985; 
        o_index_for_a6 <= 2081; 
    end
    834: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 54;
        o_index_for_a1 <= 463;
        o_index_for_a2 <= 522;
        o_index_for_a3 <= 695;
        o_index_for_a4 <= 1071;
        o_index_for_a5 <= 1986; 
        o_index_for_a6 <= 2082; 
    end
    835: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 55;
        o_index_for_a1 <= 464;
        o_index_for_a2 <= 523;
        o_index_for_a3 <= 696;
        o_index_for_a4 <= 1072;
        o_index_for_a5 <= 1987; 
        o_index_for_a6 <= 2083; 
    end
    836: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 56;
        o_index_for_a1 <= 465;
        o_index_for_a2 <= 524;
        o_index_for_a3 <= 697;
        o_index_for_a4 <= 1073;
        o_index_for_a5 <= 1988; 
        o_index_for_a6 <= 2084; 
    end
    837: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 57;
        o_index_for_a1 <= 466;
        o_index_for_a2 <= 525;
        o_index_for_a3 <= 698;
        o_index_for_a4 <= 1074;
        o_index_for_a5 <= 1989; 
        o_index_for_a6 <= 2085; 
    end
    838: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 58;
        o_index_for_a1 <= 467;
        o_index_for_a2 <= 526;
        o_index_for_a3 <= 699;
        o_index_for_a4 <= 1075;
        o_index_for_a5 <= 1990; 
        o_index_for_a6 <= 2086; 
    end
    839: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 59;
        o_index_for_a1 <= 468;
        o_index_for_a2 <= 527;
        o_index_for_a3 <= 700;
        o_index_for_a4 <= 1076;
        o_index_for_a5 <= 1991; 
        o_index_for_a6 <= 2087; 
    end
    840: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 60;
        o_index_for_a1 <= 469;
        o_index_for_a2 <= 528;
        o_index_for_a3 <= 701;
        o_index_for_a4 <= 1077;
        o_index_for_a5 <= 1992; 
        o_index_for_a6 <= 2088; 
    end
    841: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 61;
        o_index_for_a1 <= 470;
        o_index_for_a2 <= 529;
        o_index_for_a3 <= 702;
        o_index_for_a4 <= 1078;
        o_index_for_a5 <= 1993; 
        o_index_for_a6 <= 2089; 
    end
    842: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 62;
        o_index_for_a1 <= 471;
        o_index_for_a2 <= 530;
        o_index_for_a3 <= 703;
        o_index_for_a4 <= 1079;
        o_index_for_a5 <= 1994; 
        o_index_for_a6 <= 2090; 
    end
    843: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 63;
        o_index_for_a1 <= 472;
        o_index_for_a2 <= 531;
        o_index_for_a3 <= 704;
        o_index_for_a4 <= 1080;
        o_index_for_a5 <= 1995; 
        o_index_for_a6 <= 2091; 
    end
    844: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 64;
        o_index_for_a1 <= 473;
        o_index_for_a2 <= 532;
        o_index_for_a3 <= 705;
        o_index_for_a4 <= 1081;
        o_index_for_a5 <= 1996; 
        o_index_for_a6 <= 2092; 
    end
    845: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 65;
        o_index_for_a1 <= 474;
        o_index_for_a2 <= 533;
        o_index_for_a3 <= 706;
        o_index_for_a4 <= 1082;
        o_index_for_a5 <= 1997; 
        o_index_for_a6 <= 2093; 
    end
    846: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 66;
        o_index_for_a1 <= 475;
        o_index_for_a2 <= 534;
        o_index_for_a3 <= 707;
        o_index_for_a4 <= 1083;
        o_index_for_a5 <= 1998; 
        o_index_for_a6 <= 2094; 
    end
    847: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 67;
        o_index_for_a1 <= 476;
        o_index_for_a2 <= 535;
        o_index_for_a3 <= 708;
        o_index_for_a4 <= 1084;
        o_index_for_a5 <= 1999; 
        o_index_for_a6 <= 2095; 
    end
    848: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 68;
        o_index_for_a1 <= 477;
        o_index_for_a2 <= 536;
        o_index_for_a3 <= 709;
        o_index_for_a4 <= 1085;
        o_index_for_a5 <= 2000; 
        o_index_for_a6 <= 2096; 
    end
    849: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 69;
        o_index_for_a1 <= 478;
        o_index_for_a2 <= 537;
        o_index_for_a3 <= 710;
        o_index_for_a4 <= 1086;
        o_index_for_a5 <= 2001; 
        o_index_for_a6 <= 2097; 
    end
    850: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 70;
        o_index_for_a1 <= 479;
        o_index_for_a2 <= 538;
        o_index_for_a3 <= 711;
        o_index_for_a4 <= 1087;
        o_index_for_a5 <= 2002; 
        o_index_for_a6 <= 2098; 
    end
    851: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 71;
        o_index_for_a1 <= 384;
        o_index_for_a2 <= 539;
        o_index_for_a3 <= 712;
        o_index_for_a4 <= 1088;
        o_index_for_a5 <= 2003; 
        o_index_for_a6 <= 2099; 
    end
    852: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 72;
        o_index_for_a1 <= 385;
        o_index_for_a2 <= 540;
        o_index_for_a3 <= 713;
        o_index_for_a4 <= 1089;
        o_index_for_a5 <= 2004; 
        o_index_for_a6 <= 2100; 
    end
    853: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 73;
        o_index_for_a1 <= 386;
        o_index_for_a2 <= 541;
        o_index_for_a3 <= 714;
        o_index_for_a4 <= 1090;
        o_index_for_a5 <= 2005; 
        o_index_for_a6 <= 2101; 
    end
    854: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 74;
        o_index_for_a1 <= 387;
        o_index_for_a2 <= 542;
        o_index_for_a3 <= 715;
        o_index_for_a4 <= 1091;
        o_index_for_a5 <= 2006; 
        o_index_for_a6 <= 2102; 
    end
    855: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 75;
        o_index_for_a1 <= 388;
        o_index_for_a2 <= 543;
        o_index_for_a3 <= 716;
        o_index_for_a4 <= 1092;
        o_index_for_a5 <= 2007; 
        o_index_for_a6 <= 2103; 
    end
    856: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 76;
        o_index_for_a1 <= 389;
        o_index_for_a2 <= 544;
        o_index_for_a3 <= 717;
        o_index_for_a4 <= 1093;
        o_index_for_a5 <= 2008; 
        o_index_for_a6 <= 2104; 
    end
    857: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 77;
        o_index_for_a1 <= 390;
        o_index_for_a2 <= 545;
        o_index_for_a3 <= 718;
        o_index_for_a4 <= 1094;
        o_index_for_a5 <= 2009; 
        o_index_for_a6 <= 2105; 
    end
    858: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 78;
        o_index_for_a1 <= 391;
        o_index_for_a2 <= 546;
        o_index_for_a3 <= 719;
        o_index_for_a4 <= 1095;
        o_index_for_a5 <= 2010; 
        o_index_for_a6 <= 2106; 
    end
    859: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 79;
        o_index_for_a1 <= 392;
        o_index_for_a2 <= 547;
        o_index_for_a3 <= 720;
        o_index_for_a4 <= 1096;
        o_index_for_a5 <= 2011; 
        o_index_for_a6 <= 2107; 
    end
    860: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 80;
        o_index_for_a1 <= 393;
        o_index_for_a2 <= 548;
        o_index_for_a3 <= 721;
        o_index_for_a4 <= 1097;
        o_index_for_a5 <= 2012; 
        o_index_for_a6 <= 2108; 
    end
    861: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 81;
        o_index_for_a1 <= 394;
        o_index_for_a2 <= 549;
        o_index_for_a3 <= 722;
        o_index_for_a4 <= 1098;
        o_index_for_a5 <= 2013; 
        o_index_for_a6 <= 2109; 
    end
    862: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 82;
        o_index_for_a1 <= 395;
        o_index_for_a2 <= 550;
        o_index_for_a3 <= 723;
        o_index_for_a4 <= 1099;
        o_index_for_a5 <= 2014; 
        o_index_for_a6 <= 2110; 
    end
    863: begin
        o_branch_for_a0 <= 1;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 3;
        o_branch_for_a3 <= 3;
        o_branch_for_a4 <= 3;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 0; 
        o_index_for_a0 <= 83;
        o_index_for_a1 <= 396;
        o_index_for_a2 <= 551;
        o_index_for_a3 <= 724;
        o_index_for_a4 <= 1100;
        o_index_for_a5 <= 2015; 
        o_index_for_a6 <= 2111; 
    end
    864: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 482;
        o_index_for_a1 <= 709;
        o_index_for_a2 <= 986;
        o_index_for_a3 <= 1080;
        o_index_for_a4 <= 2016;
        o_index_for_a5 <= 2112; 
        o_index_for_a6 <= 2304; 
    end
    865: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 483;
        o_index_for_a1 <= 710;
        o_index_for_a2 <= 987;
        o_index_for_a3 <= 1081;
        o_index_for_a4 <= 2017;
        o_index_for_a5 <= 2113; 
        o_index_for_a6 <= 2304; 
    end
    866: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 484;
        o_index_for_a1 <= 711;
        o_index_for_a2 <= 988;
        o_index_for_a3 <= 1082;
        o_index_for_a4 <= 2018;
        o_index_for_a5 <= 2114; 
        o_index_for_a6 <= 2304; 
    end
    867: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 485;
        o_index_for_a1 <= 712;
        o_index_for_a2 <= 989;
        o_index_for_a3 <= 1083;
        o_index_for_a4 <= 2019;
        o_index_for_a5 <= 2115; 
        o_index_for_a6 <= 2304; 
    end
    868: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 486;
        o_index_for_a1 <= 713;
        o_index_for_a2 <= 990;
        o_index_for_a3 <= 1084;
        o_index_for_a4 <= 2020;
        o_index_for_a5 <= 2116; 
        o_index_for_a6 <= 2304; 
    end
    869: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 487;
        o_index_for_a1 <= 714;
        o_index_for_a2 <= 991;
        o_index_for_a3 <= 1085;
        o_index_for_a4 <= 2021;
        o_index_for_a5 <= 2117; 
        o_index_for_a6 <= 2304; 
    end
    870: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 488;
        o_index_for_a1 <= 715;
        o_index_for_a2 <= 992;
        o_index_for_a3 <= 1086;
        o_index_for_a4 <= 2022;
        o_index_for_a5 <= 2118; 
        o_index_for_a6 <= 2304; 
    end
    871: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 489;
        o_index_for_a1 <= 716;
        o_index_for_a2 <= 993;
        o_index_for_a3 <= 1087;
        o_index_for_a4 <= 2023;
        o_index_for_a5 <= 2119; 
        o_index_for_a6 <= 2304; 
    end
    872: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 490;
        o_index_for_a1 <= 717;
        o_index_for_a2 <= 994;
        o_index_for_a3 <= 1088;
        o_index_for_a4 <= 2024;
        o_index_for_a5 <= 2120; 
        o_index_for_a6 <= 2304; 
    end
    873: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 491;
        o_index_for_a1 <= 718;
        o_index_for_a2 <= 995;
        o_index_for_a3 <= 1089;
        o_index_for_a4 <= 2025;
        o_index_for_a5 <= 2121; 
        o_index_for_a6 <= 2304; 
    end
    874: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 492;
        o_index_for_a1 <= 719;
        o_index_for_a2 <= 996;
        o_index_for_a3 <= 1090;
        o_index_for_a4 <= 2026;
        o_index_for_a5 <= 2122; 
        o_index_for_a6 <= 2304; 
    end
    875: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 493;
        o_index_for_a1 <= 720;
        o_index_for_a2 <= 997;
        o_index_for_a3 <= 1091;
        o_index_for_a4 <= 2027;
        o_index_for_a5 <= 2123; 
        o_index_for_a6 <= 2304; 
    end
    876: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 494;
        o_index_for_a1 <= 721;
        o_index_for_a2 <= 998;
        o_index_for_a3 <= 1092;
        o_index_for_a4 <= 2028;
        o_index_for_a5 <= 2124; 
        o_index_for_a6 <= 2304; 
    end
    877: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 495;
        o_index_for_a1 <= 722;
        o_index_for_a2 <= 999;
        o_index_for_a3 <= 1093;
        o_index_for_a4 <= 2029;
        o_index_for_a5 <= 2125; 
        o_index_for_a6 <= 2304; 
    end
    878: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 496;
        o_index_for_a1 <= 723;
        o_index_for_a2 <= 1000;
        o_index_for_a3 <= 1094;
        o_index_for_a4 <= 2030;
        o_index_for_a5 <= 2126; 
        o_index_for_a6 <= 2304; 
    end
    879: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 497;
        o_index_for_a1 <= 724;
        o_index_for_a2 <= 1001;
        o_index_for_a3 <= 1095;
        o_index_for_a4 <= 2031;
        o_index_for_a5 <= 2127; 
        o_index_for_a6 <= 2304; 
    end
    880: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 498;
        o_index_for_a1 <= 725;
        o_index_for_a2 <= 1002;
        o_index_for_a3 <= 1096;
        o_index_for_a4 <= 2032;
        o_index_for_a5 <= 2128; 
        o_index_for_a6 <= 2304; 
    end
    881: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 499;
        o_index_for_a1 <= 726;
        o_index_for_a2 <= 1003;
        o_index_for_a3 <= 1097;
        o_index_for_a4 <= 2033;
        o_index_for_a5 <= 2129; 
        o_index_for_a6 <= 2304; 
    end
    882: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 500;
        o_index_for_a1 <= 727;
        o_index_for_a2 <= 1004;
        o_index_for_a3 <= 1098;
        o_index_for_a4 <= 2034;
        o_index_for_a5 <= 2130; 
        o_index_for_a6 <= 2304; 
    end
    883: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 501;
        o_index_for_a1 <= 728;
        o_index_for_a2 <= 1005;
        o_index_for_a3 <= 1099;
        o_index_for_a4 <= 2035;
        o_index_for_a5 <= 2131; 
        o_index_for_a6 <= 2304; 
    end
    884: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 502;
        o_index_for_a1 <= 729;
        o_index_for_a2 <= 1006;
        o_index_for_a3 <= 1100;
        o_index_for_a4 <= 2036;
        o_index_for_a5 <= 2132; 
        o_index_for_a6 <= 2304; 
    end
    885: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 503;
        o_index_for_a1 <= 730;
        o_index_for_a2 <= 1007;
        o_index_for_a3 <= 1101;
        o_index_for_a4 <= 2037;
        o_index_for_a5 <= 2133; 
        o_index_for_a6 <= 2304; 
    end
    886: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 504;
        o_index_for_a1 <= 731;
        o_index_for_a2 <= 1008;
        o_index_for_a3 <= 1102;
        o_index_for_a4 <= 2038;
        o_index_for_a5 <= 2134; 
        o_index_for_a6 <= 2304; 
    end
    887: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 505;
        o_index_for_a1 <= 732;
        o_index_for_a2 <= 1009;
        o_index_for_a3 <= 1103;
        o_index_for_a4 <= 2039;
        o_index_for_a5 <= 2135; 
        o_index_for_a6 <= 2304; 
    end
    888: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 506;
        o_index_for_a1 <= 733;
        o_index_for_a2 <= 1010;
        o_index_for_a3 <= 1104;
        o_index_for_a4 <= 2040;
        o_index_for_a5 <= 2136; 
        o_index_for_a6 <= 2304; 
    end
    889: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 507;
        o_index_for_a1 <= 734;
        o_index_for_a2 <= 1011;
        o_index_for_a3 <= 1105;
        o_index_for_a4 <= 2041;
        o_index_for_a5 <= 2137; 
        o_index_for_a6 <= 2304; 
    end
    890: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 508;
        o_index_for_a1 <= 735;
        o_index_for_a2 <= 1012;
        o_index_for_a3 <= 1106;
        o_index_for_a4 <= 2042;
        o_index_for_a5 <= 2138; 
        o_index_for_a6 <= 2304; 
    end
    891: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 509;
        o_index_for_a1 <= 736;
        o_index_for_a2 <= 1013;
        o_index_for_a3 <= 1107;
        o_index_for_a4 <= 2043;
        o_index_for_a5 <= 2139; 
        o_index_for_a6 <= 2304; 
    end
    892: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 510;
        o_index_for_a1 <= 737;
        o_index_for_a2 <= 1014;
        o_index_for_a3 <= 1108;
        o_index_for_a4 <= 2044;
        o_index_for_a5 <= 2140; 
        o_index_for_a6 <= 2304; 
    end
    893: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 511;
        o_index_for_a1 <= 738;
        o_index_for_a2 <= 1015;
        o_index_for_a3 <= 1109;
        o_index_for_a4 <= 2045;
        o_index_for_a5 <= 2141; 
        o_index_for_a6 <= 2304; 
    end
    894: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 512;
        o_index_for_a1 <= 739;
        o_index_for_a2 <= 1016;
        o_index_for_a3 <= 1110;
        o_index_for_a4 <= 2046;
        o_index_for_a5 <= 2142; 
        o_index_for_a6 <= 2304; 
    end
    895: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 513;
        o_index_for_a1 <= 740;
        o_index_for_a2 <= 1017;
        o_index_for_a3 <= 1111;
        o_index_for_a4 <= 2047;
        o_index_for_a5 <= 2143; 
        o_index_for_a6 <= 2304; 
    end
    896: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 514;
        o_index_for_a1 <= 741;
        o_index_for_a2 <= 1018;
        o_index_for_a3 <= 1112;
        o_index_for_a4 <= 2048;
        o_index_for_a5 <= 2144; 
        o_index_for_a6 <= 2304; 
    end
    897: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 515;
        o_index_for_a1 <= 742;
        o_index_for_a2 <= 1019;
        o_index_for_a3 <= 1113;
        o_index_for_a4 <= 2049;
        o_index_for_a5 <= 2145; 
        o_index_for_a6 <= 2304; 
    end
    898: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 516;
        o_index_for_a1 <= 743;
        o_index_for_a2 <= 1020;
        o_index_for_a3 <= 1114;
        o_index_for_a4 <= 2050;
        o_index_for_a5 <= 2146; 
        o_index_for_a6 <= 2304; 
    end
    899: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 517;
        o_index_for_a1 <= 744;
        o_index_for_a2 <= 1021;
        o_index_for_a3 <= 1115;
        o_index_for_a4 <= 2051;
        o_index_for_a5 <= 2147; 
        o_index_for_a6 <= 2304; 
    end
    900: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 518;
        o_index_for_a1 <= 745;
        o_index_for_a2 <= 1022;
        o_index_for_a3 <= 1116;
        o_index_for_a4 <= 2052;
        o_index_for_a5 <= 2148; 
        o_index_for_a6 <= 2304; 
    end
    901: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 519;
        o_index_for_a1 <= 746;
        o_index_for_a2 <= 1023;
        o_index_for_a3 <= 1117;
        o_index_for_a4 <= 2053;
        o_index_for_a5 <= 2149; 
        o_index_for_a6 <= 2304; 
    end
    902: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 520;
        o_index_for_a1 <= 747;
        o_index_for_a2 <= 1024;
        o_index_for_a3 <= 1118;
        o_index_for_a4 <= 2054;
        o_index_for_a5 <= 2150; 
        o_index_for_a6 <= 2304; 
    end
    903: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 521;
        o_index_for_a1 <= 748;
        o_index_for_a2 <= 1025;
        o_index_for_a3 <= 1119;
        o_index_for_a4 <= 2055;
        o_index_for_a5 <= 2151; 
        o_index_for_a6 <= 2304; 
    end
    904: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 522;
        o_index_for_a1 <= 749;
        o_index_for_a2 <= 1026;
        o_index_for_a3 <= 1120;
        o_index_for_a4 <= 2056;
        o_index_for_a5 <= 2152; 
        o_index_for_a6 <= 2304; 
    end
    905: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 523;
        o_index_for_a1 <= 750;
        o_index_for_a2 <= 1027;
        o_index_for_a3 <= 1121;
        o_index_for_a4 <= 2057;
        o_index_for_a5 <= 2153; 
        o_index_for_a6 <= 2304; 
    end
    906: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 524;
        o_index_for_a1 <= 751;
        o_index_for_a2 <= 1028;
        o_index_for_a3 <= 1122;
        o_index_for_a4 <= 2058;
        o_index_for_a5 <= 2154; 
        o_index_for_a6 <= 2304; 
    end
    907: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 525;
        o_index_for_a1 <= 752;
        o_index_for_a2 <= 1029;
        o_index_for_a3 <= 1123;
        o_index_for_a4 <= 2059;
        o_index_for_a5 <= 2155; 
        o_index_for_a6 <= 2304; 
    end
    908: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 526;
        o_index_for_a1 <= 753;
        o_index_for_a2 <= 1030;
        o_index_for_a3 <= 1124;
        o_index_for_a4 <= 2060;
        o_index_for_a5 <= 2156; 
        o_index_for_a6 <= 2304; 
    end
    909: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 527;
        o_index_for_a1 <= 754;
        o_index_for_a2 <= 1031;
        o_index_for_a3 <= 1125;
        o_index_for_a4 <= 2061;
        o_index_for_a5 <= 2157; 
        o_index_for_a6 <= 2304; 
    end
    910: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 528;
        o_index_for_a1 <= 755;
        o_index_for_a2 <= 1032;
        o_index_for_a3 <= 1126;
        o_index_for_a4 <= 2062;
        o_index_for_a5 <= 2158; 
        o_index_for_a6 <= 2304; 
    end
    911: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 529;
        o_index_for_a1 <= 756;
        o_index_for_a2 <= 1033;
        o_index_for_a3 <= 1127;
        o_index_for_a4 <= 2063;
        o_index_for_a5 <= 2159; 
        o_index_for_a6 <= 2304; 
    end
    912: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 530;
        o_index_for_a1 <= 757;
        o_index_for_a2 <= 1034;
        o_index_for_a3 <= 1128;
        o_index_for_a4 <= 2064;
        o_index_for_a5 <= 2160; 
        o_index_for_a6 <= 2304; 
    end
    913: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 531;
        o_index_for_a1 <= 758;
        o_index_for_a2 <= 1035;
        o_index_for_a3 <= 1129;
        o_index_for_a4 <= 2065;
        o_index_for_a5 <= 2161; 
        o_index_for_a6 <= 2304; 
    end
    914: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 532;
        o_index_for_a1 <= 759;
        o_index_for_a2 <= 1036;
        o_index_for_a3 <= 1130;
        o_index_for_a4 <= 2066;
        o_index_for_a5 <= 2162; 
        o_index_for_a6 <= 2304; 
    end
    915: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 533;
        o_index_for_a1 <= 760;
        o_index_for_a2 <= 1037;
        o_index_for_a3 <= 1131;
        o_index_for_a4 <= 2067;
        o_index_for_a5 <= 2163; 
        o_index_for_a6 <= 2304; 
    end
    916: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 534;
        o_index_for_a1 <= 761;
        o_index_for_a2 <= 1038;
        o_index_for_a3 <= 1132;
        o_index_for_a4 <= 2068;
        o_index_for_a5 <= 2164; 
        o_index_for_a6 <= 2304; 
    end
    917: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 535;
        o_index_for_a1 <= 762;
        o_index_for_a2 <= 1039;
        o_index_for_a3 <= 1133;
        o_index_for_a4 <= 2069;
        o_index_for_a5 <= 2165; 
        o_index_for_a6 <= 2304; 
    end
    918: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 536;
        o_index_for_a1 <= 763;
        o_index_for_a2 <= 1040;
        o_index_for_a3 <= 1134;
        o_index_for_a4 <= 2070;
        o_index_for_a5 <= 2166; 
        o_index_for_a6 <= 2304; 
    end
    919: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 537;
        o_index_for_a1 <= 764;
        o_index_for_a2 <= 1041;
        o_index_for_a3 <= 1135;
        o_index_for_a4 <= 2071;
        o_index_for_a5 <= 2167; 
        o_index_for_a6 <= 2304; 
    end
    920: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 538;
        o_index_for_a1 <= 765;
        o_index_for_a2 <= 1042;
        o_index_for_a3 <= 1136;
        o_index_for_a4 <= 2072;
        o_index_for_a5 <= 2168; 
        o_index_for_a6 <= 2304; 
    end
    921: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 539;
        o_index_for_a1 <= 766;
        o_index_for_a2 <= 1043;
        o_index_for_a3 <= 1137;
        o_index_for_a4 <= 2073;
        o_index_for_a5 <= 2169; 
        o_index_for_a6 <= 2304; 
    end
    922: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 540;
        o_index_for_a1 <= 767;
        o_index_for_a2 <= 1044;
        o_index_for_a3 <= 1138;
        o_index_for_a4 <= 2074;
        o_index_for_a5 <= 2170; 
        o_index_for_a6 <= 2304; 
    end
    923: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 541;
        o_index_for_a1 <= 672;
        o_index_for_a2 <= 1045;
        o_index_for_a3 <= 1139;
        o_index_for_a4 <= 2075;
        o_index_for_a5 <= 2171; 
        o_index_for_a6 <= 2304; 
    end
    924: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 542;
        o_index_for_a1 <= 673;
        o_index_for_a2 <= 1046;
        o_index_for_a3 <= 1140;
        o_index_for_a4 <= 2076;
        o_index_for_a5 <= 2172; 
        o_index_for_a6 <= 2304; 
    end
    925: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 543;
        o_index_for_a1 <= 674;
        o_index_for_a2 <= 1047;
        o_index_for_a3 <= 1141;
        o_index_for_a4 <= 2077;
        o_index_for_a5 <= 2173; 
        o_index_for_a6 <= 2304; 
    end
    926: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 544;
        o_index_for_a1 <= 675;
        o_index_for_a2 <= 1048;
        o_index_for_a3 <= 1142;
        o_index_for_a4 <= 2078;
        o_index_for_a5 <= 2174; 
        o_index_for_a6 <= 2304; 
    end
    927: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 545;
        o_index_for_a1 <= 676;
        o_index_for_a2 <= 1049;
        o_index_for_a3 <= 1143;
        o_index_for_a4 <= 2079;
        o_index_for_a5 <= 2175; 
        o_index_for_a6 <= 2304; 
    end
    928: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 546;
        o_index_for_a1 <= 677;
        o_index_for_a2 <= 1050;
        o_index_for_a3 <= 1144;
        o_index_for_a4 <= 2080;
        o_index_for_a5 <= 2176; 
        o_index_for_a6 <= 2304; 
    end
    929: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 547;
        o_index_for_a1 <= 678;
        o_index_for_a2 <= 1051;
        o_index_for_a3 <= 1145;
        o_index_for_a4 <= 2081;
        o_index_for_a5 <= 2177; 
        o_index_for_a6 <= 2304; 
    end
    930: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 548;
        o_index_for_a1 <= 679;
        o_index_for_a2 <= 1052;
        o_index_for_a3 <= 1146;
        o_index_for_a4 <= 2082;
        o_index_for_a5 <= 2178; 
        o_index_for_a6 <= 2304; 
    end
    931: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 549;
        o_index_for_a1 <= 680;
        o_index_for_a2 <= 1053;
        o_index_for_a3 <= 1147;
        o_index_for_a4 <= 2083;
        o_index_for_a5 <= 2179; 
        o_index_for_a6 <= 2304; 
    end
    932: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 550;
        o_index_for_a1 <= 681;
        o_index_for_a2 <= 1054;
        o_index_for_a3 <= 1148;
        o_index_for_a4 <= 2084;
        o_index_for_a5 <= 2180; 
        o_index_for_a6 <= 2304; 
    end
    933: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 551;
        o_index_for_a1 <= 682;
        o_index_for_a2 <= 1055;
        o_index_for_a3 <= 1149;
        o_index_for_a4 <= 2085;
        o_index_for_a5 <= 2181; 
        o_index_for_a6 <= 2304; 
    end
    934: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 552;
        o_index_for_a1 <= 683;
        o_index_for_a2 <= 960;
        o_index_for_a3 <= 1150;
        o_index_for_a4 <= 2086;
        o_index_for_a5 <= 2182; 
        o_index_for_a6 <= 2304; 
    end
    935: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 553;
        o_index_for_a1 <= 684;
        o_index_for_a2 <= 961;
        o_index_for_a3 <= 1151;
        o_index_for_a4 <= 2087;
        o_index_for_a5 <= 2183; 
        o_index_for_a6 <= 2304; 
    end
    936: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 554;
        o_index_for_a1 <= 685;
        o_index_for_a2 <= 962;
        o_index_for_a3 <= 1056;
        o_index_for_a4 <= 2088;
        o_index_for_a5 <= 2184; 
        o_index_for_a6 <= 2304; 
    end
    937: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 555;
        o_index_for_a1 <= 686;
        o_index_for_a2 <= 963;
        o_index_for_a3 <= 1057;
        o_index_for_a4 <= 2089;
        o_index_for_a5 <= 2185; 
        o_index_for_a6 <= 2304; 
    end
    938: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 556;
        o_index_for_a1 <= 687;
        o_index_for_a2 <= 964;
        o_index_for_a3 <= 1058;
        o_index_for_a4 <= 2090;
        o_index_for_a5 <= 2186; 
        o_index_for_a6 <= 2304; 
    end
    939: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 557;
        o_index_for_a1 <= 688;
        o_index_for_a2 <= 965;
        o_index_for_a3 <= 1059;
        o_index_for_a4 <= 2091;
        o_index_for_a5 <= 2187; 
        o_index_for_a6 <= 2304; 
    end
    940: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 558;
        o_index_for_a1 <= 689;
        o_index_for_a2 <= 966;
        o_index_for_a3 <= 1060;
        o_index_for_a4 <= 2092;
        o_index_for_a5 <= 2188; 
        o_index_for_a6 <= 2304; 
    end
    941: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 559;
        o_index_for_a1 <= 690;
        o_index_for_a2 <= 967;
        o_index_for_a3 <= 1061;
        o_index_for_a4 <= 2093;
        o_index_for_a5 <= 2189; 
        o_index_for_a6 <= 2304; 
    end
    942: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 560;
        o_index_for_a1 <= 691;
        o_index_for_a2 <= 968;
        o_index_for_a3 <= 1062;
        o_index_for_a4 <= 2094;
        o_index_for_a5 <= 2190; 
        o_index_for_a6 <= 2304; 
    end
    943: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 561;
        o_index_for_a1 <= 692;
        o_index_for_a2 <= 969;
        o_index_for_a3 <= 1063;
        o_index_for_a4 <= 2095;
        o_index_for_a5 <= 2191; 
        o_index_for_a6 <= 2304; 
    end
    944: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 562;
        o_index_for_a1 <= 693;
        o_index_for_a2 <= 970;
        o_index_for_a3 <= 1064;
        o_index_for_a4 <= 2096;
        o_index_for_a5 <= 2192; 
        o_index_for_a6 <= 2304; 
    end
    945: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 563;
        o_index_for_a1 <= 694;
        o_index_for_a2 <= 971;
        o_index_for_a3 <= 1065;
        o_index_for_a4 <= 2097;
        o_index_for_a5 <= 2193; 
        o_index_for_a6 <= 2304; 
    end
    946: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 564;
        o_index_for_a1 <= 695;
        o_index_for_a2 <= 972;
        o_index_for_a3 <= 1066;
        o_index_for_a4 <= 2098;
        o_index_for_a5 <= 2194; 
        o_index_for_a6 <= 2304; 
    end
    947: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 565;
        o_index_for_a1 <= 696;
        o_index_for_a2 <= 973;
        o_index_for_a3 <= 1067;
        o_index_for_a4 <= 2099;
        o_index_for_a5 <= 2195; 
        o_index_for_a6 <= 2304; 
    end
    948: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 566;
        o_index_for_a1 <= 697;
        o_index_for_a2 <= 974;
        o_index_for_a3 <= 1068;
        o_index_for_a4 <= 2100;
        o_index_for_a5 <= 2196; 
        o_index_for_a6 <= 2304; 
    end
    949: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 567;
        o_index_for_a1 <= 698;
        o_index_for_a2 <= 975;
        o_index_for_a3 <= 1069;
        o_index_for_a4 <= 2101;
        o_index_for_a5 <= 2197; 
        o_index_for_a6 <= 2304; 
    end
    950: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 568;
        o_index_for_a1 <= 699;
        o_index_for_a2 <= 976;
        o_index_for_a3 <= 1070;
        o_index_for_a4 <= 2102;
        o_index_for_a5 <= 2198; 
        o_index_for_a6 <= 2304; 
    end
    951: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 569;
        o_index_for_a1 <= 700;
        o_index_for_a2 <= 977;
        o_index_for_a3 <= 1071;
        o_index_for_a4 <= 2103;
        o_index_for_a5 <= 2199; 
        o_index_for_a6 <= 2304; 
    end
    952: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 570;
        o_index_for_a1 <= 701;
        o_index_for_a2 <= 978;
        o_index_for_a3 <= 1072;
        o_index_for_a4 <= 2104;
        o_index_for_a5 <= 2200; 
        o_index_for_a6 <= 2304; 
    end
    953: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 571;
        o_index_for_a1 <= 702;
        o_index_for_a2 <= 979;
        o_index_for_a3 <= 1073;
        o_index_for_a4 <= 2105;
        o_index_for_a5 <= 2201; 
        o_index_for_a6 <= 2304; 
    end
    954: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 572;
        o_index_for_a1 <= 703;
        o_index_for_a2 <= 980;
        o_index_for_a3 <= 1074;
        o_index_for_a4 <= 2106;
        o_index_for_a5 <= 2202; 
        o_index_for_a6 <= 2304; 
    end
    955: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 573;
        o_index_for_a1 <= 704;
        o_index_for_a2 <= 981;
        o_index_for_a3 <= 1075;
        o_index_for_a4 <= 2107;
        o_index_for_a5 <= 2203; 
        o_index_for_a6 <= 2304; 
    end
    956: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 574;
        o_index_for_a1 <= 705;
        o_index_for_a2 <= 982;
        o_index_for_a3 <= 1076;
        o_index_for_a4 <= 2108;
        o_index_for_a5 <= 2204; 
        o_index_for_a6 <= 2304; 
    end
    957: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 575;
        o_index_for_a1 <= 706;
        o_index_for_a2 <= 983;
        o_index_for_a3 <= 1077;
        o_index_for_a4 <= 2109;
        o_index_for_a5 <= 2205; 
        o_index_for_a6 <= 2304; 
    end
    958: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 480;
        o_index_for_a1 <= 707;
        o_index_for_a2 <= 984;
        o_index_for_a3 <= 1078;
        o_index_for_a4 <= 2110;
        o_index_for_a5 <= 2206; 
        o_index_for_a6 <= 2304; 
    end
    959: begin
        o_branch_for_a0 <= 4;
        o_branch_for_a1 <= 4;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 4;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 481;
        o_index_for_a1 <= 708;
        o_index_for_a2 <= 985;
        o_index_for_a3 <= 1079;
        o_index_for_a4 <= 2111;
        o_index_for_a5 <= 2207; 
        o_index_for_a6 <= 2304; 
    end
    960: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 281;
        o_index_for_a1 <= 319;
        o_index_for_a2 <= 825;
        o_index_for_a3 <= 911;
        o_index_for_a4 <= 2112;
        o_index_for_a5 <= 2208; 
        o_index_for_a6 <= 2304; 
    end
    961: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 282;
        o_index_for_a1 <= 320;
        o_index_for_a2 <= 826;
        o_index_for_a3 <= 912;
        o_index_for_a4 <= 2113;
        o_index_for_a5 <= 2209; 
        o_index_for_a6 <= 2304; 
    end
    962: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 283;
        o_index_for_a1 <= 321;
        o_index_for_a2 <= 827;
        o_index_for_a3 <= 913;
        o_index_for_a4 <= 2114;
        o_index_for_a5 <= 2210; 
        o_index_for_a6 <= 2304; 
    end
    963: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 284;
        o_index_for_a1 <= 322;
        o_index_for_a2 <= 828;
        o_index_for_a3 <= 914;
        o_index_for_a4 <= 2115;
        o_index_for_a5 <= 2211; 
        o_index_for_a6 <= 2304; 
    end
    964: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 285;
        o_index_for_a1 <= 323;
        o_index_for_a2 <= 829;
        o_index_for_a3 <= 915;
        o_index_for_a4 <= 2116;
        o_index_for_a5 <= 2212; 
        o_index_for_a6 <= 2304; 
    end
    965: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 286;
        o_index_for_a1 <= 324;
        o_index_for_a2 <= 830;
        o_index_for_a3 <= 916;
        o_index_for_a4 <= 2117;
        o_index_for_a5 <= 2213; 
        o_index_for_a6 <= 2304; 
    end
    966: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 287;
        o_index_for_a1 <= 325;
        o_index_for_a2 <= 831;
        o_index_for_a3 <= 917;
        o_index_for_a4 <= 2118;
        o_index_for_a5 <= 2214; 
        o_index_for_a6 <= 2304; 
    end
    967: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 192;
        o_index_for_a1 <= 326;
        o_index_for_a2 <= 832;
        o_index_for_a3 <= 918;
        o_index_for_a4 <= 2119;
        o_index_for_a5 <= 2215; 
        o_index_for_a6 <= 2304; 
    end
    968: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 193;
        o_index_for_a1 <= 327;
        o_index_for_a2 <= 833;
        o_index_for_a3 <= 919;
        o_index_for_a4 <= 2120;
        o_index_for_a5 <= 2216; 
        o_index_for_a6 <= 2304; 
    end
    969: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 194;
        o_index_for_a1 <= 328;
        o_index_for_a2 <= 834;
        o_index_for_a3 <= 920;
        o_index_for_a4 <= 2121;
        o_index_for_a5 <= 2217; 
        o_index_for_a6 <= 2304; 
    end
    970: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 195;
        o_index_for_a1 <= 329;
        o_index_for_a2 <= 835;
        o_index_for_a3 <= 921;
        o_index_for_a4 <= 2122;
        o_index_for_a5 <= 2218; 
        o_index_for_a6 <= 2304; 
    end
    971: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 196;
        o_index_for_a1 <= 330;
        o_index_for_a2 <= 836;
        o_index_for_a3 <= 922;
        o_index_for_a4 <= 2123;
        o_index_for_a5 <= 2219; 
        o_index_for_a6 <= 2304; 
    end
    972: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 197;
        o_index_for_a1 <= 331;
        o_index_for_a2 <= 837;
        o_index_for_a3 <= 923;
        o_index_for_a4 <= 2124;
        o_index_for_a5 <= 2220; 
        o_index_for_a6 <= 2304; 
    end
    973: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 198;
        o_index_for_a1 <= 332;
        o_index_for_a2 <= 838;
        o_index_for_a3 <= 924;
        o_index_for_a4 <= 2125;
        o_index_for_a5 <= 2221; 
        o_index_for_a6 <= 2304; 
    end
    974: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 199;
        o_index_for_a1 <= 333;
        o_index_for_a2 <= 839;
        o_index_for_a3 <= 925;
        o_index_for_a4 <= 2126;
        o_index_for_a5 <= 2222; 
        o_index_for_a6 <= 2304; 
    end
    975: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 200;
        o_index_for_a1 <= 334;
        o_index_for_a2 <= 840;
        o_index_for_a3 <= 926;
        o_index_for_a4 <= 2127;
        o_index_for_a5 <= 2223; 
        o_index_for_a6 <= 2304; 
    end
    976: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 201;
        o_index_for_a1 <= 335;
        o_index_for_a2 <= 841;
        o_index_for_a3 <= 927;
        o_index_for_a4 <= 2128;
        o_index_for_a5 <= 2224; 
        o_index_for_a6 <= 2304; 
    end
    977: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 202;
        o_index_for_a1 <= 336;
        o_index_for_a2 <= 842;
        o_index_for_a3 <= 928;
        o_index_for_a4 <= 2129;
        o_index_for_a5 <= 2225; 
        o_index_for_a6 <= 2304; 
    end
    978: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 203;
        o_index_for_a1 <= 337;
        o_index_for_a2 <= 843;
        o_index_for_a3 <= 929;
        o_index_for_a4 <= 2130;
        o_index_for_a5 <= 2226; 
        o_index_for_a6 <= 2304; 
    end
    979: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 204;
        o_index_for_a1 <= 338;
        o_index_for_a2 <= 844;
        o_index_for_a3 <= 930;
        o_index_for_a4 <= 2131;
        o_index_for_a5 <= 2227; 
        o_index_for_a6 <= 2304; 
    end
    980: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 205;
        o_index_for_a1 <= 339;
        o_index_for_a2 <= 845;
        o_index_for_a3 <= 931;
        o_index_for_a4 <= 2132;
        o_index_for_a5 <= 2228; 
        o_index_for_a6 <= 2304; 
    end
    981: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 206;
        o_index_for_a1 <= 340;
        o_index_for_a2 <= 846;
        o_index_for_a3 <= 932;
        o_index_for_a4 <= 2133;
        o_index_for_a5 <= 2229; 
        o_index_for_a6 <= 2304; 
    end
    982: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 207;
        o_index_for_a1 <= 341;
        o_index_for_a2 <= 847;
        o_index_for_a3 <= 933;
        o_index_for_a4 <= 2134;
        o_index_for_a5 <= 2230; 
        o_index_for_a6 <= 2304; 
    end
    983: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 208;
        o_index_for_a1 <= 342;
        o_index_for_a2 <= 848;
        o_index_for_a3 <= 934;
        o_index_for_a4 <= 2135;
        o_index_for_a5 <= 2231; 
        o_index_for_a6 <= 2304; 
    end
    984: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 209;
        o_index_for_a1 <= 343;
        o_index_for_a2 <= 849;
        o_index_for_a3 <= 935;
        o_index_for_a4 <= 2136;
        o_index_for_a5 <= 2232; 
        o_index_for_a6 <= 2304; 
    end
    985: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 210;
        o_index_for_a1 <= 344;
        o_index_for_a2 <= 850;
        o_index_for_a3 <= 936;
        o_index_for_a4 <= 2137;
        o_index_for_a5 <= 2233; 
        o_index_for_a6 <= 2304; 
    end
    986: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 211;
        o_index_for_a1 <= 345;
        o_index_for_a2 <= 851;
        o_index_for_a3 <= 937;
        o_index_for_a4 <= 2138;
        o_index_for_a5 <= 2234; 
        o_index_for_a6 <= 2304; 
    end
    987: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 212;
        o_index_for_a1 <= 346;
        o_index_for_a2 <= 852;
        o_index_for_a3 <= 938;
        o_index_for_a4 <= 2139;
        o_index_for_a5 <= 2235; 
        o_index_for_a6 <= 2304; 
    end
    988: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 213;
        o_index_for_a1 <= 347;
        o_index_for_a2 <= 853;
        o_index_for_a3 <= 939;
        o_index_for_a4 <= 2140;
        o_index_for_a5 <= 2236; 
        o_index_for_a6 <= 2304; 
    end
    989: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 214;
        o_index_for_a1 <= 348;
        o_index_for_a2 <= 854;
        o_index_for_a3 <= 940;
        o_index_for_a4 <= 2141;
        o_index_for_a5 <= 2237; 
        o_index_for_a6 <= 2304; 
    end
    990: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 215;
        o_index_for_a1 <= 349;
        o_index_for_a2 <= 855;
        o_index_for_a3 <= 941;
        o_index_for_a4 <= 2142;
        o_index_for_a5 <= 2238; 
        o_index_for_a6 <= 2304; 
    end
    991: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 216;
        o_index_for_a1 <= 350;
        o_index_for_a2 <= 856;
        o_index_for_a3 <= 942;
        o_index_for_a4 <= 2143;
        o_index_for_a5 <= 2239; 
        o_index_for_a6 <= 2304; 
    end
    992: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 217;
        o_index_for_a1 <= 351;
        o_index_for_a2 <= 857;
        o_index_for_a3 <= 943;
        o_index_for_a4 <= 2144;
        o_index_for_a5 <= 2240; 
        o_index_for_a6 <= 2304; 
    end
    993: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 218;
        o_index_for_a1 <= 352;
        o_index_for_a2 <= 858;
        o_index_for_a3 <= 944;
        o_index_for_a4 <= 2145;
        o_index_for_a5 <= 2241; 
        o_index_for_a6 <= 2304; 
    end
    994: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 219;
        o_index_for_a1 <= 353;
        o_index_for_a2 <= 859;
        o_index_for_a3 <= 945;
        o_index_for_a4 <= 2146;
        o_index_for_a5 <= 2242; 
        o_index_for_a6 <= 2304; 
    end
    995: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 220;
        o_index_for_a1 <= 354;
        o_index_for_a2 <= 860;
        o_index_for_a3 <= 946;
        o_index_for_a4 <= 2147;
        o_index_for_a5 <= 2243; 
        o_index_for_a6 <= 2304; 
    end
    996: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 221;
        o_index_for_a1 <= 355;
        o_index_for_a2 <= 861;
        o_index_for_a3 <= 947;
        o_index_for_a4 <= 2148;
        o_index_for_a5 <= 2244; 
        o_index_for_a6 <= 2304; 
    end
    997: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 222;
        o_index_for_a1 <= 356;
        o_index_for_a2 <= 862;
        o_index_for_a3 <= 948;
        o_index_for_a4 <= 2149;
        o_index_for_a5 <= 2245; 
        o_index_for_a6 <= 2304; 
    end
    998: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 223;
        o_index_for_a1 <= 357;
        o_index_for_a2 <= 863;
        o_index_for_a3 <= 949;
        o_index_for_a4 <= 2150;
        o_index_for_a5 <= 2246; 
        o_index_for_a6 <= 2304; 
    end
    999: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 224;
        o_index_for_a1 <= 358;
        o_index_for_a2 <= 768;
        o_index_for_a3 <= 950;
        o_index_for_a4 <= 2151;
        o_index_for_a5 <= 2247; 
        o_index_for_a6 <= 2304; 
    end
    1000: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 225;
        o_index_for_a1 <= 359;
        o_index_for_a2 <= 769;
        o_index_for_a3 <= 951;
        o_index_for_a4 <= 2152;
        o_index_for_a5 <= 2248; 
        o_index_for_a6 <= 2304; 
    end
    1001: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 226;
        o_index_for_a1 <= 360;
        o_index_for_a2 <= 770;
        o_index_for_a3 <= 952;
        o_index_for_a4 <= 2153;
        o_index_for_a5 <= 2249; 
        o_index_for_a6 <= 2304; 
    end
    1002: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 227;
        o_index_for_a1 <= 361;
        o_index_for_a2 <= 771;
        o_index_for_a3 <= 953;
        o_index_for_a4 <= 2154;
        o_index_for_a5 <= 2250; 
        o_index_for_a6 <= 2304; 
    end
    1003: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 228;
        o_index_for_a1 <= 362;
        o_index_for_a2 <= 772;
        o_index_for_a3 <= 954;
        o_index_for_a4 <= 2155;
        o_index_for_a5 <= 2251; 
        o_index_for_a6 <= 2304; 
    end
    1004: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 229;
        o_index_for_a1 <= 363;
        o_index_for_a2 <= 773;
        o_index_for_a3 <= 955;
        o_index_for_a4 <= 2156;
        o_index_for_a5 <= 2252; 
        o_index_for_a6 <= 2304; 
    end
    1005: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 230;
        o_index_for_a1 <= 364;
        o_index_for_a2 <= 774;
        o_index_for_a3 <= 956;
        o_index_for_a4 <= 2157;
        o_index_for_a5 <= 2253; 
        o_index_for_a6 <= 2304; 
    end
    1006: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 231;
        o_index_for_a1 <= 365;
        o_index_for_a2 <= 775;
        o_index_for_a3 <= 957;
        o_index_for_a4 <= 2158;
        o_index_for_a5 <= 2254; 
        o_index_for_a6 <= 2304; 
    end
    1007: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 232;
        o_index_for_a1 <= 366;
        o_index_for_a2 <= 776;
        o_index_for_a3 <= 958;
        o_index_for_a4 <= 2159;
        o_index_for_a5 <= 2255; 
        o_index_for_a6 <= 2304; 
    end
    1008: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 233;
        o_index_for_a1 <= 367;
        o_index_for_a2 <= 777;
        o_index_for_a3 <= 959;
        o_index_for_a4 <= 2160;
        o_index_for_a5 <= 2256; 
        o_index_for_a6 <= 2304; 
    end
    1009: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 234;
        o_index_for_a1 <= 368;
        o_index_for_a2 <= 778;
        o_index_for_a3 <= 864;
        o_index_for_a4 <= 2161;
        o_index_for_a5 <= 2257; 
        o_index_for_a6 <= 2304; 
    end
    1010: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 235;
        o_index_for_a1 <= 369;
        o_index_for_a2 <= 779;
        o_index_for_a3 <= 865;
        o_index_for_a4 <= 2162;
        o_index_for_a5 <= 2258; 
        o_index_for_a6 <= 2304; 
    end
    1011: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 236;
        o_index_for_a1 <= 370;
        o_index_for_a2 <= 780;
        o_index_for_a3 <= 866;
        o_index_for_a4 <= 2163;
        o_index_for_a5 <= 2259; 
        o_index_for_a6 <= 2304; 
    end
    1012: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 237;
        o_index_for_a1 <= 371;
        o_index_for_a2 <= 781;
        o_index_for_a3 <= 867;
        o_index_for_a4 <= 2164;
        o_index_for_a5 <= 2260; 
        o_index_for_a6 <= 2304; 
    end
    1013: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 238;
        o_index_for_a1 <= 372;
        o_index_for_a2 <= 782;
        o_index_for_a3 <= 868;
        o_index_for_a4 <= 2165;
        o_index_for_a5 <= 2261; 
        o_index_for_a6 <= 2304; 
    end
    1014: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 239;
        o_index_for_a1 <= 373;
        o_index_for_a2 <= 783;
        o_index_for_a3 <= 869;
        o_index_for_a4 <= 2166;
        o_index_for_a5 <= 2262; 
        o_index_for_a6 <= 2304; 
    end
    1015: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 240;
        o_index_for_a1 <= 374;
        o_index_for_a2 <= 784;
        o_index_for_a3 <= 870;
        o_index_for_a4 <= 2167;
        o_index_for_a5 <= 2263; 
        o_index_for_a6 <= 2304; 
    end
    1016: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 241;
        o_index_for_a1 <= 375;
        o_index_for_a2 <= 785;
        o_index_for_a3 <= 871;
        o_index_for_a4 <= 2168;
        o_index_for_a5 <= 2264; 
        o_index_for_a6 <= 2304; 
    end
    1017: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 242;
        o_index_for_a1 <= 376;
        o_index_for_a2 <= 786;
        o_index_for_a3 <= 872;
        o_index_for_a4 <= 2169;
        o_index_for_a5 <= 2265; 
        o_index_for_a6 <= 2304; 
    end
    1018: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 243;
        o_index_for_a1 <= 377;
        o_index_for_a2 <= 787;
        o_index_for_a3 <= 873;
        o_index_for_a4 <= 2170;
        o_index_for_a5 <= 2266; 
        o_index_for_a6 <= 2304; 
    end
    1019: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 244;
        o_index_for_a1 <= 378;
        o_index_for_a2 <= 788;
        o_index_for_a3 <= 874;
        o_index_for_a4 <= 2171;
        o_index_for_a5 <= 2267; 
        o_index_for_a6 <= 2304; 
    end
    1020: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 245;
        o_index_for_a1 <= 379;
        o_index_for_a2 <= 789;
        o_index_for_a3 <= 875;
        o_index_for_a4 <= 2172;
        o_index_for_a5 <= 2268; 
        o_index_for_a6 <= 2304; 
    end
    1021: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 246;
        o_index_for_a1 <= 380;
        o_index_for_a2 <= 790;
        o_index_for_a3 <= 876;
        o_index_for_a4 <= 2173;
        o_index_for_a5 <= 2269; 
        o_index_for_a6 <= 2304; 
    end
    1022: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 247;
        o_index_for_a1 <= 381;
        o_index_for_a2 <= 791;
        o_index_for_a3 <= 877;
        o_index_for_a4 <= 2174;
        o_index_for_a5 <= 2270; 
        o_index_for_a6 <= 2304; 
    end
    1023: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 248;
        o_index_for_a1 <= 382;
        o_index_for_a2 <= 792;
        o_index_for_a3 <= 878;
        o_index_for_a4 <= 2175;
        o_index_for_a5 <= 2271; 
        o_index_for_a6 <= 2304; 
    end
    1024: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 249;
        o_index_for_a1 <= 383;
        o_index_for_a2 <= 793;
        o_index_for_a3 <= 879;
        o_index_for_a4 <= 2176;
        o_index_for_a5 <= 2272; 
        o_index_for_a6 <= 2304; 
    end
    1025: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 250;
        o_index_for_a1 <= 288;
        o_index_for_a2 <= 794;
        o_index_for_a3 <= 880;
        o_index_for_a4 <= 2177;
        o_index_for_a5 <= 2273; 
        o_index_for_a6 <= 2304; 
    end
    1026: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 251;
        o_index_for_a1 <= 289;
        o_index_for_a2 <= 795;
        o_index_for_a3 <= 881;
        o_index_for_a4 <= 2178;
        o_index_for_a5 <= 2274; 
        o_index_for_a6 <= 2304; 
    end
    1027: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 252;
        o_index_for_a1 <= 290;
        o_index_for_a2 <= 796;
        o_index_for_a3 <= 882;
        o_index_for_a4 <= 2179;
        o_index_for_a5 <= 2275; 
        o_index_for_a6 <= 2304; 
    end
    1028: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 253;
        o_index_for_a1 <= 291;
        o_index_for_a2 <= 797;
        o_index_for_a3 <= 883;
        o_index_for_a4 <= 2180;
        o_index_for_a5 <= 2276; 
        o_index_for_a6 <= 2304; 
    end
    1029: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 254;
        o_index_for_a1 <= 292;
        o_index_for_a2 <= 798;
        o_index_for_a3 <= 884;
        o_index_for_a4 <= 2181;
        o_index_for_a5 <= 2277; 
        o_index_for_a6 <= 2304; 
    end
    1030: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 255;
        o_index_for_a1 <= 293;
        o_index_for_a2 <= 799;
        o_index_for_a3 <= 885;
        o_index_for_a4 <= 2182;
        o_index_for_a5 <= 2278; 
        o_index_for_a6 <= 2304; 
    end
    1031: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 256;
        o_index_for_a1 <= 294;
        o_index_for_a2 <= 800;
        o_index_for_a3 <= 886;
        o_index_for_a4 <= 2183;
        o_index_for_a5 <= 2279; 
        o_index_for_a6 <= 2304; 
    end
    1032: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 257;
        o_index_for_a1 <= 295;
        o_index_for_a2 <= 801;
        o_index_for_a3 <= 887;
        o_index_for_a4 <= 2184;
        o_index_for_a5 <= 2280; 
        o_index_for_a6 <= 2304; 
    end
    1033: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 258;
        o_index_for_a1 <= 296;
        o_index_for_a2 <= 802;
        o_index_for_a3 <= 888;
        o_index_for_a4 <= 2185;
        o_index_for_a5 <= 2281; 
        o_index_for_a6 <= 2304; 
    end
    1034: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 259;
        o_index_for_a1 <= 297;
        o_index_for_a2 <= 803;
        o_index_for_a3 <= 889;
        o_index_for_a4 <= 2186;
        o_index_for_a5 <= 2282; 
        o_index_for_a6 <= 2304; 
    end
    1035: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 260;
        o_index_for_a1 <= 298;
        o_index_for_a2 <= 804;
        o_index_for_a3 <= 890;
        o_index_for_a4 <= 2187;
        o_index_for_a5 <= 2283; 
        o_index_for_a6 <= 2304; 
    end
    1036: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 261;
        o_index_for_a1 <= 299;
        o_index_for_a2 <= 805;
        o_index_for_a3 <= 891;
        o_index_for_a4 <= 2188;
        o_index_for_a5 <= 2284; 
        o_index_for_a6 <= 2304; 
    end
    1037: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 262;
        o_index_for_a1 <= 300;
        o_index_for_a2 <= 806;
        o_index_for_a3 <= 892;
        o_index_for_a4 <= 2189;
        o_index_for_a5 <= 2285; 
        o_index_for_a6 <= 2304; 
    end
    1038: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 263;
        o_index_for_a1 <= 301;
        o_index_for_a2 <= 807;
        o_index_for_a3 <= 893;
        o_index_for_a4 <= 2190;
        o_index_for_a5 <= 2286; 
        o_index_for_a6 <= 2304; 
    end
    1039: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 264;
        o_index_for_a1 <= 302;
        o_index_for_a2 <= 808;
        o_index_for_a3 <= 894;
        o_index_for_a4 <= 2191;
        o_index_for_a5 <= 2287; 
        o_index_for_a6 <= 2304; 
    end
    1040: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 265;
        o_index_for_a1 <= 303;
        o_index_for_a2 <= 809;
        o_index_for_a3 <= 895;
        o_index_for_a4 <= 2192;
        o_index_for_a5 <= 2288; 
        o_index_for_a6 <= 2304; 
    end
    1041: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 266;
        o_index_for_a1 <= 304;
        o_index_for_a2 <= 810;
        o_index_for_a3 <= 896;
        o_index_for_a4 <= 2193;
        o_index_for_a5 <= 2289; 
        o_index_for_a6 <= 2304; 
    end
    1042: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 267;
        o_index_for_a1 <= 305;
        o_index_for_a2 <= 811;
        o_index_for_a3 <= 897;
        o_index_for_a4 <= 2194;
        o_index_for_a5 <= 2290; 
        o_index_for_a6 <= 2304; 
    end
    1043: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 268;
        o_index_for_a1 <= 306;
        o_index_for_a2 <= 812;
        o_index_for_a3 <= 898;
        o_index_for_a4 <= 2195;
        o_index_for_a5 <= 2291; 
        o_index_for_a6 <= 2304; 
    end
    1044: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 269;
        o_index_for_a1 <= 307;
        o_index_for_a2 <= 813;
        o_index_for_a3 <= 899;
        o_index_for_a4 <= 2196;
        o_index_for_a5 <= 2292; 
        o_index_for_a6 <= 2304; 
    end
    1045: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 270;
        o_index_for_a1 <= 308;
        o_index_for_a2 <= 814;
        o_index_for_a3 <= 900;
        o_index_for_a4 <= 2197;
        o_index_for_a5 <= 2293; 
        o_index_for_a6 <= 2304; 
    end
    1046: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 271;
        o_index_for_a1 <= 309;
        o_index_for_a2 <= 815;
        o_index_for_a3 <= 901;
        o_index_for_a4 <= 2198;
        o_index_for_a5 <= 2294; 
        o_index_for_a6 <= 2304; 
    end
    1047: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 272;
        o_index_for_a1 <= 310;
        o_index_for_a2 <= 816;
        o_index_for_a3 <= 902;
        o_index_for_a4 <= 2199;
        o_index_for_a5 <= 2295; 
        o_index_for_a6 <= 2304; 
    end
    1048: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 273;
        o_index_for_a1 <= 311;
        o_index_for_a2 <= 817;
        o_index_for_a3 <= 903;
        o_index_for_a4 <= 2200;
        o_index_for_a5 <= 2296; 
        o_index_for_a6 <= 2304; 
    end
    1049: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 274;
        o_index_for_a1 <= 312;
        o_index_for_a2 <= 818;
        o_index_for_a3 <= 904;
        o_index_for_a4 <= 2201;
        o_index_for_a5 <= 2297; 
        o_index_for_a6 <= 2304; 
    end
    1050: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 275;
        o_index_for_a1 <= 313;
        o_index_for_a2 <= 819;
        o_index_for_a3 <= 905;
        o_index_for_a4 <= 2202;
        o_index_for_a5 <= 2298; 
        o_index_for_a6 <= 2304; 
    end
    1051: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 276;
        o_index_for_a1 <= 314;
        o_index_for_a2 <= 820;
        o_index_for_a3 <= 906;
        o_index_for_a4 <= 2203;
        o_index_for_a5 <= 2299; 
        o_index_for_a6 <= 2304; 
    end
    1052: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 277;
        o_index_for_a1 <= 315;
        o_index_for_a2 <= 821;
        o_index_for_a3 <= 907;
        o_index_for_a4 <= 2204;
        o_index_for_a5 <= 2300; 
        o_index_for_a6 <= 2304; 
    end
    1053: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 278;
        o_index_for_a1 <= 316;
        o_index_for_a2 <= 822;
        o_index_for_a3 <= 908;
        o_index_for_a4 <= 2205;
        o_index_for_a5 <= 2301; 
        o_index_for_a6 <= 2304; 
    end
    1054: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 279;
        o_index_for_a1 <= 317;
        o_index_for_a2 <= 823;
        o_index_for_a3 <= 909;
        o_index_for_a4 <= 2206;
        o_index_for_a5 <= 2302; 
        o_index_for_a6 <= 2304; 
    end
    1055: begin
        o_branch_for_a0 <= 5;
        o_branch_for_a1 <= 2;
        o_branch_for_a2 <= 2;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 1;
        o_branch_for_a5 <= 0; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 280;
        o_index_for_a1 <= 318;
        o_index_for_a2 <= 824;
        o_index_for_a3 <= 910;
        o_index_for_a4 <= 2207;
        o_index_for_a5 <= 2303; 
        o_index_for_a6 <= 2304; 
    end
    1056: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 53;
        o_index_for_a1 <= 510;
        o_index_for_a2 <= 727;
        o_index_for_a3 <= 1126;
        o_index_for_a4 <= 1241;
        o_index_for_a5 <= 2208; 
        o_index_for_a6 <= 2304; 
    end
    1057: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 54;
        o_index_for_a1 <= 511;
        o_index_for_a2 <= 728;
        o_index_for_a3 <= 1127;
        o_index_for_a4 <= 1242;
        o_index_for_a5 <= 2209; 
        o_index_for_a6 <= 2304; 
    end
    1058: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 55;
        o_index_for_a1 <= 512;
        o_index_for_a2 <= 729;
        o_index_for_a3 <= 1128;
        o_index_for_a4 <= 1243;
        o_index_for_a5 <= 2210; 
        o_index_for_a6 <= 2304; 
    end
    1059: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 56;
        o_index_for_a1 <= 513;
        o_index_for_a2 <= 730;
        o_index_for_a3 <= 1129;
        o_index_for_a4 <= 1244;
        o_index_for_a5 <= 2211; 
        o_index_for_a6 <= 2304; 
    end
    1060: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 57;
        o_index_for_a1 <= 514;
        o_index_for_a2 <= 731;
        o_index_for_a3 <= 1130;
        o_index_for_a4 <= 1245;
        o_index_for_a5 <= 2212; 
        o_index_for_a6 <= 2304; 
    end
    1061: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 58;
        o_index_for_a1 <= 515;
        o_index_for_a2 <= 732;
        o_index_for_a3 <= 1131;
        o_index_for_a4 <= 1246;
        o_index_for_a5 <= 2213; 
        o_index_for_a6 <= 2304; 
    end
    1062: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 59;
        o_index_for_a1 <= 516;
        o_index_for_a2 <= 733;
        o_index_for_a3 <= 1132;
        o_index_for_a4 <= 1247;
        o_index_for_a5 <= 2214; 
        o_index_for_a6 <= 2304; 
    end
    1063: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 60;
        o_index_for_a1 <= 517;
        o_index_for_a2 <= 734;
        o_index_for_a3 <= 1133;
        o_index_for_a4 <= 1152;
        o_index_for_a5 <= 2215; 
        o_index_for_a6 <= 2304; 
    end
    1064: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 61;
        o_index_for_a1 <= 518;
        o_index_for_a2 <= 735;
        o_index_for_a3 <= 1134;
        o_index_for_a4 <= 1153;
        o_index_for_a5 <= 2216; 
        o_index_for_a6 <= 2304; 
    end
    1065: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 62;
        o_index_for_a1 <= 519;
        o_index_for_a2 <= 736;
        o_index_for_a3 <= 1135;
        o_index_for_a4 <= 1154;
        o_index_for_a5 <= 2217; 
        o_index_for_a6 <= 2304; 
    end
    1066: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 63;
        o_index_for_a1 <= 520;
        o_index_for_a2 <= 737;
        o_index_for_a3 <= 1136;
        o_index_for_a4 <= 1155;
        o_index_for_a5 <= 2218; 
        o_index_for_a6 <= 2304; 
    end
    1067: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 64;
        o_index_for_a1 <= 521;
        o_index_for_a2 <= 738;
        o_index_for_a3 <= 1137;
        o_index_for_a4 <= 1156;
        o_index_for_a5 <= 2219; 
        o_index_for_a6 <= 2304; 
    end
    1068: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 65;
        o_index_for_a1 <= 522;
        o_index_for_a2 <= 739;
        o_index_for_a3 <= 1138;
        o_index_for_a4 <= 1157;
        o_index_for_a5 <= 2220; 
        o_index_for_a6 <= 2304; 
    end
    1069: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 66;
        o_index_for_a1 <= 523;
        o_index_for_a2 <= 740;
        o_index_for_a3 <= 1139;
        o_index_for_a4 <= 1158;
        o_index_for_a5 <= 2221; 
        o_index_for_a6 <= 2304; 
    end
    1070: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 67;
        o_index_for_a1 <= 524;
        o_index_for_a2 <= 741;
        o_index_for_a3 <= 1140;
        o_index_for_a4 <= 1159;
        o_index_for_a5 <= 2222; 
        o_index_for_a6 <= 2304; 
    end
    1071: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 68;
        o_index_for_a1 <= 525;
        o_index_for_a2 <= 742;
        o_index_for_a3 <= 1141;
        o_index_for_a4 <= 1160;
        o_index_for_a5 <= 2223; 
        o_index_for_a6 <= 2304; 
    end
    1072: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 69;
        o_index_for_a1 <= 526;
        o_index_for_a2 <= 743;
        o_index_for_a3 <= 1142;
        o_index_for_a4 <= 1161;
        o_index_for_a5 <= 2224; 
        o_index_for_a6 <= 2304; 
    end
    1073: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 70;
        o_index_for_a1 <= 527;
        o_index_for_a2 <= 744;
        o_index_for_a3 <= 1143;
        o_index_for_a4 <= 1162;
        o_index_for_a5 <= 2225; 
        o_index_for_a6 <= 2304; 
    end
    1074: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 71;
        o_index_for_a1 <= 528;
        o_index_for_a2 <= 745;
        o_index_for_a3 <= 1144;
        o_index_for_a4 <= 1163;
        o_index_for_a5 <= 2226; 
        o_index_for_a6 <= 2304; 
    end
    1075: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 72;
        o_index_for_a1 <= 529;
        o_index_for_a2 <= 746;
        o_index_for_a3 <= 1145;
        o_index_for_a4 <= 1164;
        o_index_for_a5 <= 2227; 
        o_index_for_a6 <= 2304; 
    end
    1076: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 73;
        o_index_for_a1 <= 530;
        o_index_for_a2 <= 747;
        o_index_for_a3 <= 1146;
        o_index_for_a4 <= 1165;
        o_index_for_a5 <= 2228; 
        o_index_for_a6 <= 2304; 
    end
    1077: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 74;
        o_index_for_a1 <= 531;
        o_index_for_a2 <= 748;
        o_index_for_a3 <= 1147;
        o_index_for_a4 <= 1166;
        o_index_for_a5 <= 2229; 
        o_index_for_a6 <= 2304; 
    end
    1078: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 75;
        o_index_for_a1 <= 532;
        o_index_for_a2 <= 749;
        o_index_for_a3 <= 1148;
        o_index_for_a4 <= 1167;
        o_index_for_a5 <= 2230; 
        o_index_for_a6 <= 2304; 
    end
    1079: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 76;
        o_index_for_a1 <= 533;
        o_index_for_a2 <= 750;
        o_index_for_a3 <= 1149;
        o_index_for_a4 <= 1168;
        o_index_for_a5 <= 2231; 
        o_index_for_a6 <= 2304; 
    end
    1080: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 77;
        o_index_for_a1 <= 534;
        o_index_for_a2 <= 751;
        o_index_for_a3 <= 1150;
        o_index_for_a4 <= 1169;
        o_index_for_a5 <= 2232; 
        o_index_for_a6 <= 2304; 
    end
    1081: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 78;
        o_index_for_a1 <= 535;
        o_index_for_a2 <= 752;
        o_index_for_a3 <= 1151;
        o_index_for_a4 <= 1170;
        o_index_for_a5 <= 2233; 
        o_index_for_a6 <= 2304; 
    end
    1082: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 79;
        o_index_for_a1 <= 536;
        o_index_for_a2 <= 753;
        o_index_for_a3 <= 1056;
        o_index_for_a4 <= 1171;
        o_index_for_a5 <= 2234; 
        o_index_for_a6 <= 2304; 
    end
    1083: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 80;
        o_index_for_a1 <= 537;
        o_index_for_a2 <= 754;
        o_index_for_a3 <= 1057;
        o_index_for_a4 <= 1172;
        o_index_for_a5 <= 2235; 
        o_index_for_a6 <= 2304; 
    end
    1084: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 81;
        o_index_for_a1 <= 538;
        o_index_for_a2 <= 755;
        o_index_for_a3 <= 1058;
        o_index_for_a4 <= 1173;
        o_index_for_a5 <= 2236; 
        o_index_for_a6 <= 2304; 
    end
    1085: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 82;
        o_index_for_a1 <= 539;
        o_index_for_a2 <= 756;
        o_index_for_a3 <= 1059;
        o_index_for_a4 <= 1174;
        o_index_for_a5 <= 2237; 
        o_index_for_a6 <= 2304; 
    end
    1086: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 83;
        o_index_for_a1 <= 540;
        o_index_for_a2 <= 757;
        o_index_for_a3 <= 1060;
        o_index_for_a4 <= 1175;
        o_index_for_a5 <= 2238; 
        o_index_for_a6 <= 2304; 
    end
    1087: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 84;
        o_index_for_a1 <= 541;
        o_index_for_a2 <= 758;
        o_index_for_a3 <= 1061;
        o_index_for_a4 <= 1176;
        o_index_for_a5 <= 2239; 
        o_index_for_a6 <= 2304; 
    end
    1088: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 85;
        o_index_for_a1 <= 542;
        o_index_for_a2 <= 759;
        o_index_for_a3 <= 1062;
        o_index_for_a4 <= 1177;
        o_index_for_a5 <= 2240; 
        o_index_for_a6 <= 2304; 
    end
    1089: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 86;
        o_index_for_a1 <= 543;
        o_index_for_a2 <= 760;
        o_index_for_a3 <= 1063;
        o_index_for_a4 <= 1178;
        o_index_for_a5 <= 2241; 
        o_index_for_a6 <= 2304; 
    end
    1090: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 87;
        o_index_for_a1 <= 544;
        o_index_for_a2 <= 761;
        o_index_for_a3 <= 1064;
        o_index_for_a4 <= 1179;
        o_index_for_a5 <= 2242; 
        o_index_for_a6 <= 2304; 
    end
    1091: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 88;
        o_index_for_a1 <= 545;
        o_index_for_a2 <= 762;
        o_index_for_a3 <= 1065;
        o_index_for_a4 <= 1180;
        o_index_for_a5 <= 2243; 
        o_index_for_a6 <= 2304; 
    end
    1092: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 89;
        o_index_for_a1 <= 546;
        o_index_for_a2 <= 763;
        o_index_for_a3 <= 1066;
        o_index_for_a4 <= 1181;
        o_index_for_a5 <= 2244; 
        o_index_for_a6 <= 2304; 
    end
    1093: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 90;
        o_index_for_a1 <= 547;
        o_index_for_a2 <= 764;
        o_index_for_a3 <= 1067;
        o_index_for_a4 <= 1182;
        o_index_for_a5 <= 2245; 
        o_index_for_a6 <= 2304; 
    end
    1094: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 91;
        o_index_for_a1 <= 548;
        o_index_for_a2 <= 765;
        o_index_for_a3 <= 1068;
        o_index_for_a4 <= 1183;
        o_index_for_a5 <= 2246; 
        o_index_for_a6 <= 2304; 
    end
    1095: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 92;
        o_index_for_a1 <= 549;
        o_index_for_a2 <= 766;
        o_index_for_a3 <= 1069;
        o_index_for_a4 <= 1184;
        o_index_for_a5 <= 2247; 
        o_index_for_a6 <= 2304; 
    end
    1096: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 93;
        o_index_for_a1 <= 550;
        o_index_for_a2 <= 767;
        o_index_for_a3 <= 1070;
        o_index_for_a4 <= 1185;
        o_index_for_a5 <= 2248; 
        o_index_for_a6 <= 2304; 
    end
    1097: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 94;
        o_index_for_a1 <= 551;
        o_index_for_a2 <= 672;
        o_index_for_a3 <= 1071;
        o_index_for_a4 <= 1186;
        o_index_for_a5 <= 2249; 
        o_index_for_a6 <= 2304; 
    end
    1098: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 95;
        o_index_for_a1 <= 552;
        o_index_for_a2 <= 673;
        o_index_for_a3 <= 1072;
        o_index_for_a4 <= 1187;
        o_index_for_a5 <= 2250; 
        o_index_for_a6 <= 2304; 
    end
    1099: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 0;
        o_index_for_a1 <= 553;
        o_index_for_a2 <= 674;
        o_index_for_a3 <= 1073;
        o_index_for_a4 <= 1188;
        o_index_for_a5 <= 2251; 
        o_index_for_a6 <= 2304; 
    end
    1100: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 1;
        o_index_for_a1 <= 554;
        o_index_for_a2 <= 675;
        o_index_for_a3 <= 1074;
        o_index_for_a4 <= 1189;
        o_index_for_a5 <= 2252; 
        o_index_for_a6 <= 2304; 
    end
    1101: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 2;
        o_index_for_a1 <= 555;
        o_index_for_a2 <= 676;
        o_index_for_a3 <= 1075;
        o_index_for_a4 <= 1190;
        o_index_for_a5 <= 2253; 
        o_index_for_a6 <= 2304; 
    end
    1102: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 3;
        o_index_for_a1 <= 556;
        o_index_for_a2 <= 677;
        o_index_for_a3 <= 1076;
        o_index_for_a4 <= 1191;
        o_index_for_a5 <= 2254; 
        o_index_for_a6 <= 2304; 
    end
    1103: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 4;
        o_index_for_a1 <= 557;
        o_index_for_a2 <= 678;
        o_index_for_a3 <= 1077;
        o_index_for_a4 <= 1192;
        o_index_for_a5 <= 2255; 
        o_index_for_a6 <= 2304; 
    end
    1104: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 5;
        o_index_for_a1 <= 558;
        o_index_for_a2 <= 679;
        o_index_for_a3 <= 1078;
        o_index_for_a4 <= 1193;
        o_index_for_a5 <= 2256; 
        o_index_for_a6 <= 2304; 
    end
    1105: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 6;
        o_index_for_a1 <= 559;
        o_index_for_a2 <= 680;
        o_index_for_a3 <= 1079;
        o_index_for_a4 <= 1194;
        o_index_for_a5 <= 2257; 
        o_index_for_a6 <= 2304; 
    end
    1106: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 7;
        o_index_for_a1 <= 560;
        o_index_for_a2 <= 681;
        o_index_for_a3 <= 1080;
        o_index_for_a4 <= 1195;
        o_index_for_a5 <= 2258; 
        o_index_for_a6 <= 2304; 
    end
    1107: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 8;
        o_index_for_a1 <= 561;
        o_index_for_a2 <= 682;
        o_index_for_a3 <= 1081;
        o_index_for_a4 <= 1196;
        o_index_for_a5 <= 2259; 
        o_index_for_a6 <= 2304; 
    end
    1108: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 9;
        o_index_for_a1 <= 562;
        o_index_for_a2 <= 683;
        o_index_for_a3 <= 1082;
        o_index_for_a4 <= 1197;
        o_index_for_a5 <= 2260; 
        o_index_for_a6 <= 2304; 
    end
    1109: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 10;
        o_index_for_a1 <= 563;
        o_index_for_a2 <= 684;
        o_index_for_a3 <= 1083;
        o_index_for_a4 <= 1198;
        o_index_for_a5 <= 2261; 
        o_index_for_a6 <= 2304; 
    end
    1110: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 11;
        o_index_for_a1 <= 564;
        o_index_for_a2 <= 685;
        o_index_for_a3 <= 1084;
        o_index_for_a4 <= 1199;
        o_index_for_a5 <= 2262; 
        o_index_for_a6 <= 2304; 
    end
    1111: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 12;
        o_index_for_a1 <= 565;
        o_index_for_a2 <= 686;
        o_index_for_a3 <= 1085;
        o_index_for_a4 <= 1200;
        o_index_for_a5 <= 2263; 
        o_index_for_a6 <= 2304; 
    end
    1112: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 13;
        o_index_for_a1 <= 566;
        o_index_for_a2 <= 687;
        o_index_for_a3 <= 1086;
        o_index_for_a4 <= 1201;
        o_index_for_a5 <= 2264; 
        o_index_for_a6 <= 2304; 
    end
    1113: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 14;
        o_index_for_a1 <= 567;
        o_index_for_a2 <= 688;
        o_index_for_a3 <= 1087;
        o_index_for_a4 <= 1202;
        o_index_for_a5 <= 2265; 
        o_index_for_a6 <= 2304; 
    end
    1114: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 15;
        o_index_for_a1 <= 568;
        o_index_for_a2 <= 689;
        o_index_for_a3 <= 1088;
        o_index_for_a4 <= 1203;
        o_index_for_a5 <= 2266; 
        o_index_for_a6 <= 2304; 
    end
    1115: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 16;
        o_index_for_a1 <= 569;
        o_index_for_a2 <= 690;
        o_index_for_a3 <= 1089;
        o_index_for_a4 <= 1204;
        o_index_for_a5 <= 2267; 
        o_index_for_a6 <= 2304; 
    end
    1116: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 17;
        o_index_for_a1 <= 570;
        o_index_for_a2 <= 691;
        o_index_for_a3 <= 1090;
        o_index_for_a4 <= 1205;
        o_index_for_a5 <= 2268; 
        o_index_for_a6 <= 2304; 
    end
    1117: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 18;
        o_index_for_a1 <= 571;
        o_index_for_a2 <= 692;
        o_index_for_a3 <= 1091;
        o_index_for_a4 <= 1206;
        o_index_for_a5 <= 2269; 
        o_index_for_a6 <= 2304; 
    end
    1118: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 19;
        o_index_for_a1 <= 572;
        o_index_for_a2 <= 693;
        o_index_for_a3 <= 1092;
        o_index_for_a4 <= 1207;
        o_index_for_a5 <= 2270; 
        o_index_for_a6 <= 2304; 
    end
    1119: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 20;
        o_index_for_a1 <= 573;
        o_index_for_a2 <= 694;
        o_index_for_a3 <= 1093;
        o_index_for_a4 <= 1208;
        o_index_for_a5 <= 2271; 
        o_index_for_a6 <= 2304; 
    end
    1120: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 21;
        o_index_for_a1 <= 574;
        o_index_for_a2 <= 695;
        o_index_for_a3 <= 1094;
        o_index_for_a4 <= 1209;
        o_index_for_a5 <= 2272; 
        o_index_for_a6 <= 2304; 
    end
    1121: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 22;
        o_index_for_a1 <= 575;
        o_index_for_a2 <= 696;
        o_index_for_a3 <= 1095;
        o_index_for_a4 <= 1210;
        o_index_for_a5 <= 2273; 
        o_index_for_a6 <= 2304; 
    end
    1122: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 23;
        o_index_for_a1 <= 480;
        o_index_for_a2 <= 697;
        o_index_for_a3 <= 1096;
        o_index_for_a4 <= 1211;
        o_index_for_a5 <= 2274; 
        o_index_for_a6 <= 2304; 
    end
    1123: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 24;
        o_index_for_a1 <= 481;
        o_index_for_a2 <= 698;
        o_index_for_a3 <= 1097;
        o_index_for_a4 <= 1212;
        o_index_for_a5 <= 2275; 
        o_index_for_a6 <= 2304; 
    end
    1124: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 25;
        o_index_for_a1 <= 482;
        o_index_for_a2 <= 699;
        o_index_for_a3 <= 1098;
        o_index_for_a4 <= 1213;
        o_index_for_a5 <= 2276; 
        o_index_for_a6 <= 2304; 
    end
    1125: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 26;
        o_index_for_a1 <= 483;
        o_index_for_a2 <= 700;
        o_index_for_a3 <= 1099;
        o_index_for_a4 <= 1214;
        o_index_for_a5 <= 2277; 
        o_index_for_a6 <= 2304; 
    end
    1126: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 27;
        o_index_for_a1 <= 484;
        o_index_for_a2 <= 701;
        o_index_for_a3 <= 1100;
        o_index_for_a4 <= 1215;
        o_index_for_a5 <= 2278; 
        o_index_for_a6 <= 2304; 
    end
    1127: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 28;
        o_index_for_a1 <= 485;
        o_index_for_a2 <= 702;
        o_index_for_a3 <= 1101;
        o_index_for_a4 <= 1216;
        o_index_for_a5 <= 2279; 
        o_index_for_a6 <= 2304; 
    end
    1128: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 29;
        o_index_for_a1 <= 486;
        o_index_for_a2 <= 703;
        o_index_for_a3 <= 1102;
        o_index_for_a4 <= 1217;
        o_index_for_a5 <= 2280; 
        o_index_for_a6 <= 2304; 
    end
    1129: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 30;
        o_index_for_a1 <= 487;
        o_index_for_a2 <= 704;
        o_index_for_a3 <= 1103;
        o_index_for_a4 <= 1218;
        o_index_for_a5 <= 2281; 
        o_index_for_a6 <= 2304; 
    end
    1130: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 31;
        o_index_for_a1 <= 488;
        o_index_for_a2 <= 705;
        o_index_for_a3 <= 1104;
        o_index_for_a4 <= 1219;
        o_index_for_a5 <= 2282; 
        o_index_for_a6 <= 2304; 
    end
    1131: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 32;
        o_index_for_a1 <= 489;
        o_index_for_a2 <= 706;
        o_index_for_a3 <= 1105;
        o_index_for_a4 <= 1220;
        o_index_for_a5 <= 2283; 
        o_index_for_a6 <= 2304; 
    end
    1132: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 33;
        o_index_for_a1 <= 490;
        o_index_for_a2 <= 707;
        o_index_for_a3 <= 1106;
        o_index_for_a4 <= 1221;
        o_index_for_a5 <= 2284; 
        o_index_for_a6 <= 2304; 
    end
    1133: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 34;
        o_index_for_a1 <= 491;
        o_index_for_a2 <= 708;
        o_index_for_a3 <= 1107;
        o_index_for_a4 <= 1222;
        o_index_for_a5 <= 2285; 
        o_index_for_a6 <= 2304; 
    end
    1134: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 35;
        o_index_for_a1 <= 492;
        o_index_for_a2 <= 709;
        o_index_for_a3 <= 1108;
        o_index_for_a4 <= 1223;
        o_index_for_a5 <= 2286; 
        o_index_for_a6 <= 2304; 
    end
    1135: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 36;
        o_index_for_a1 <= 493;
        o_index_for_a2 <= 710;
        o_index_for_a3 <= 1109;
        o_index_for_a4 <= 1224;
        o_index_for_a5 <= 2287; 
        o_index_for_a6 <= 2304; 
    end
    1136: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 37;
        o_index_for_a1 <= 494;
        o_index_for_a2 <= 711;
        o_index_for_a3 <= 1110;
        o_index_for_a4 <= 1225;
        o_index_for_a5 <= 2288; 
        o_index_for_a6 <= 2304; 
    end
    1137: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 38;
        o_index_for_a1 <= 495;
        o_index_for_a2 <= 712;
        o_index_for_a3 <= 1111;
        o_index_for_a4 <= 1226;
        o_index_for_a5 <= 2289; 
        o_index_for_a6 <= 2304; 
    end
    1138: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 39;
        o_index_for_a1 <= 496;
        o_index_for_a2 <= 713;
        o_index_for_a3 <= 1112;
        o_index_for_a4 <= 1227;
        o_index_for_a5 <= 2290; 
        o_index_for_a6 <= 2304; 
    end
    1139: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 40;
        o_index_for_a1 <= 497;
        o_index_for_a2 <= 714;
        o_index_for_a3 <= 1113;
        o_index_for_a4 <= 1228;
        o_index_for_a5 <= 2291; 
        o_index_for_a6 <= 2304; 
    end
    1140: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 41;
        o_index_for_a1 <= 498;
        o_index_for_a2 <= 715;
        o_index_for_a3 <= 1114;
        o_index_for_a4 <= 1229;
        o_index_for_a5 <= 2292; 
        o_index_for_a6 <= 2304; 
    end
    1141: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 42;
        o_index_for_a1 <= 499;
        o_index_for_a2 <= 716;
        o_index_for_a3 <= 1115;
        o_index_for_a4 <= 1230;
        o_index_for_a5 <= 2293; 
        o_index_for_a6 <= 2304; 
    end
    1142: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 43;
        o_index_for_a1 <= 500;
        o_index_for_a2 <= 717;
        o_index_for_a3 <= 1116;
        o_index_for_a4 <= 1231;
        o_index_for_a5 <= 2294; 
        o_index_for_a6 <= 2304; 
    end
    1143: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 44;
        o_index_for_a1 <= 501;
        o_index_for_a2 <= 718;
        o_index_for_a3 <= 1117;
        o_index_for_a4 <= 1232;
        o_index_for_a5 <= 2295; 
        o_index_for_a6 <= 2304; 
    end
    1144: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 45;
        o_index_for_a1 <= 502;
        o_index_for_a2 <= 719;
        o_index_for_a3 <= 1118;
        o_index_for_a4 <= 1233;
        o_index_for_a5 <= 2296; 
        o_index_for_a6 <= 2304; 
    end
    1145: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 46;
        o_index_for_a1 <= 503;
        o_index_for_a2 <= 720;
        o_index_for_a3 <= 1119;
        o_index_for_a4 <= 1234;
        o_index_for_a5 <= 2297; 
        o_index_for_a6 <= 2304; 
    end
    1146: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 47;
        o_index_for_a1 <= 504;
        o_index_for_a2 <= 721;
        o_index_for_a3 <= 1120;
        o_index_for_a4 <= 1235;
        o_index_for_a5 <= 2298; 
        o_index_for_a6 <= 2304; 
    end
    1147: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 48;
        o_index_for_a1 <= 505;
        o_index_for_a2 <= 722;
        o_index_for_a3 <= 1121;
        o_index_for_a4 <= 1236;
        o_index_for_a5 <= 2299; 
        o_index_for_a6 <= 2304; 
    end
    1148: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 49;
        o_index_for_a1 <= 506;
        o_index_for_a2 <= 723;
        o_index_for_a3 <= 1122;
        o_index_for_a4 <= 1237;
        o_index_for_a5 <= 2300; 
        o_index_for_a6 <= 2304; 
    end
    1149: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 50;
        o_index_for_a1 <= 507;
        o_index_for_a2 <= 724;
        o_index_for_a3 <= 1123;
        o_index_for_a4 <= 1238;
        o_index_for_a5 <= 2301; 
        o_index_for_a6 <= 2304; 
    end
    1150: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 51;
        o_index_for_a1 <= 508;
        o_index_for_a2 <= 725;
        o_index_for_a3 <= 1124;
        o_index_for_a4 <= 1239;
        o_index_for_a5 <= 2302; 
        o_index_for_a6 <= 2304; 
    end
    1151: begin
        o_branch_for_a0 <= 2;
        o_branch_for_a1 <= 5;
        o_branch_for_a2 <= 5;
        o_branch_for_a3 <= 5;
        o_branch_for_a4 <= 2;
        o_branch_for_a5 <= 1; 
        o_branch_for_a6 <= 7; 
        o_index_for_a0 <= 52;
        o_index_for_a1 <= 509;
        o_index_for_a2 <= 726;
        o_index_for_a3 <= 1125;
        o_index_for_a4 <= 1240;
        o_index_for_a5 <= 2303; 
        o_index_for_a6 <= 2304; 
    end
    default: begin // This case is for simulation purposes only.
        o_branch_for_a0 <= 'x;
        o_branch_for_a1 <= 'x;
        o_branch_for_a2 <= 'x;
        o_branch_for_a3 <= 'x;
        o_branch_for_a4 <= 'x;
        o_branch_for_a5 <= 'x; 
        o_branch_for_a6 <= 'x; 
        o_index_for_a0 <= 'x;
        o_index_for_a1 <= 'x;
        o_index_for_a2 <= 'x;
        o_index_for_a3 <= 'x;
        o_index_for_a4 <= 'x;
        o_index_for_a5 <= 'x; 
        o_index_for_a6 <= 'x; 
    end
    endcase
end

endmodule: ldpc_row_to_column_rom

`default_nettype wire
