
typedef struct {
    logic [15:0] magnitude;
    logic        sign;
} belief_t;
