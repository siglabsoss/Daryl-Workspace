// tb_ldpc_encoder.sv

`timescale 10ps / 10ps

`default_nettype none

module tb_ldpc_encoder;

localparam integer WIDTH = 8;

// Clock and Reset
logic                i_clock;
logic                i_reset;
// Upstream signaling
logic [WIDTH-1:0]    i_in_data;
logic                i_in_valid;
logic                o_in_ready;
// Downstream signaling
logic [WIDTH-1:0]    o_out_data;
logic                o_out_valid;
logic                i_out_ready;

localparam CLENGTH = 2304;
localparam SLENGTH = CLENGTH / 2;
localparam logic [0:CLENGTH-1] ldpc_codeword_0 = {
    32'b01000111100000001110001001110101,
    32'b10100000101010111101001000011000,
    32'b11010100110011111001001010001011,
    32'b10011011101111110110110010110000,
    32'b10001111000000011100010011101011,
    32'b01000001010101111010010000110001,
    32'b10101001100111110010010100010111,
    32'b00110111011111101101100101100001,
    32'b00011110000000111000100111010110,
    32'b10000010101011110100100001100011,
    32'b01010011001111100100101000101110,
    32'b01101110111111011011001011000010,
    32'b00111100000001110001001110101101,
    32'b00000101010111101001000011000110,
    32'b10100110011111001001010001011100,
    32'b11011101111110110110010110000100,
    32'b01111000000011100010011101011010,
    32'b00001010101111010010000110001101,
    32'b01001100111110010010100010111001,
    32'b10111011111101101100101100001000,
    32'b11110000000111000100111010110100,
    32'b00010101011110100100001100011010,
    32'b10011001111100100101000101110011,
    32'b01110111111011011001011000010001,
    32'b11100000001110001001110101101000,
    32'b00101010111101001000011000110101,
    32'b00110011111001001010001011100110,
    32'b11101111110110110010110000100011,
    32'b11000000011100010011101011010000,
    32'b01010101111010010000110001101010,
    32'b01100111110010010100010111001101,
    32'b11011111101101100101100001000111,
    32'b10000000111000100111010110100000,
    32'b10101011110100100001100011010100,
    32'b11001111100100101000101110011011,
    32'b10111111011011001011000010001111,
    32'b01011000111110110011101001110010,
    32'b00101011001100111010111111011100,
    32'b11011101010101000111001101010001,
    32'b11001011010111111110100110110011,
    32'b10000110110000011011001001001011,
    32'b00000111000001110111101000011100,
    32'b01000100001011100010111100011010,
    32'b10001010101010111101010110000010,
    32'b01000010110010100001011010101100,
    32'b11101001001010110111001010110011,
    32'b01101111001011111010110110001100,
    32'b01100101100100000101010010010000,
    32'b10111111010010111010100000011111,
    32'b10101110100110100010101001111011,
    32'b01011011001110000000111101011110,
    32'b01001010000010010111011001101101,
    32'b00011101100011101001010011010011,
    32'b00000000001110100100011111111011,
    32'b10101010100011010101000110010101,
    32'b01101001011110111001001101010100,
    32'b00010011001110010011110100001101,
    32'b10100111001000011100111001010010,
    32'b00001011111011000100001110101010,
    32'b00101000001011011000001110100101,
    32'b11001100000101111110011100101111,
    32'b01011011010110101100111100100010,
    32'b00111010010100011111010110001100,
    32'b11000100111010100011100000001000,
    32'b00000001010011101100111100011010,
    32'b10100111001110011100001101000111,
    32'b01101110111111001100101110011101,
    32'b10011001011110000111010100110110,
    32'b00101100101100011101000100101100,
    32'b10011101001111110011001101110001,
    32'b11001011100111010101011100110010,
    32'b11101001100111100111101100111010
};

// Example from Behrooze
// {
//     32'b01000111100000001110001001110101,
//     32'b10100000101010111101001000011000,
//     32'b11010100110011111001001010001011,
//     32'b10011011101111110110110010110000,
//     32'b10001111000000011100010011101011,
//     32'b01000001010101111010010000110001,
//     32'b10101001100111110010010100010111,
//     32'b00110111011111101101100101100001,
//     32'b00011110000000111000100111010110,
//     32'b10000010101011110100100001100011,
//     32'b01010011001111100100101000101110,
//     32'b01101110111111011011001011000010,
//     32'b00111100000001110001001110101101,
//     32'b00000101010111101001000011000110,
//     32'b10100110011111001001010001011100,
//     32'b11011101111110110110010110000100,
//     32'b01111000000011100010011101011010,
//     32'b00001010101111010010000110001101,
//     32'b01001100111110010010100010111001,
//     32'b10111011111101101100101100001000,
//     32'b11110000000111000100111010110100,
//     32'b00010101011110100100001100011010,
//     32'b10011001111100100101000101110011,
//     32'b01110111111011011001011000010001,
//     32'b11100000001110001001110101101000,
//     32'b00101010111101001000011000110101,
//     32'b00110011111001001010001011100110,
//     32'b11101111110110110010110000100011,
//     32'b11000000011100010011101011010000,
//     32'b01010101111010010000110001101010,
//     32'b01100111110010010100010111001101,
//     32'b11011111101101100101100001000111,
//     32'b10000000111000100111010110100000,
//     32'b10101011110100100001100011010100,
//     32'b11001111100100101000101110011011,
//     32'b10111111011011001011000010001111,
//     32'b11101011110101100100000100000001,
//     32'b10010101111011110110100100011001,
//     32'b00111100010100111101001111000010,
//     32'b11110011000100100111101000111101,
//     32'b11111000010100001100110000001101,
//     32'b01100110100110010001111101001110,
//     32'b11100100001001010010100000100101,
//     32'b00101100100111110101111010000110,
//     32'b11111100100100110011101001101011,
//     32'b10110111000110100100000000001111,
//     32'b11011000000110010110101110110100,
//     32'b11110010001100101011011100100111,
//     32'b11100001011110101001101011100111,
//     32'b00010100110110001100101111111101,
//     32'b01010100100110101110110011101001,
//     32'b10110101010100101110010100110110,
//     32'b10000101110110101000011111000101,
//     32'b00101011100001110110011010110110,
//     32'b11110100100100011101011110100010,
//     32'b10001000000000110110110000000000,
//     32'b00101000010110100111000001011011,
//     32'b00111001101011000001010001011010,
//     32'b01100100010001100100001110101010,
//     32'b00111110101010101111011110101010,
//     32'b01101011010101101011010101100011,
//     32'b00111101110001010110110000000000,
//     32'b00101000010110010110001110100010,
//     32'b10001101101111100110000110101100,
//     32'b10101111010010111010000010100010,
//     32'b11001110001001111011011100000000,
//     32'b00110101010100100011001111001111,
//     32'b00011001101010100101110011010100,
//     32'b11100111010110101110011110110111,
//     32'b00101000110110000110110010011010,
//     32'b01001001000111001101000001011011,
//     32'b00000100111010111010110001001000
// };

logic [0:CLENGTH-1] ldpc_encoded_codeword_0;

ldpc_encoder uut (.*);

always begin: clock_gen
    #5 i_clock = 1'b1;
    #5 i_clock = 1'b0;
end

// debug variable declarations
logic [31:0] glbl_err_count = 0;
logic [31:0] test_number = 1;
logic [31:0] run_count = 0;
logic [31:0] count = 0;

// Used by check process, declared here so it
// can be included in the final tall for the
// global error count.
logic [31:0] local_err_count = 0;

task reset_all;
    i_reset = 1'b1;
    i_in_data = 0;
    i_in_valid = 1'b0;
    i_out_ready = 1'b0;
    #1000;
    @(negedge i_clock) i_reset = 1'b0;
endtask: reset_all

initial begin: stimulus
    i_reset = 1'b1;
    #1000;
    reset_all();

    // Test 1: No data in = no data out.
    $display("Test 1 Started!");
    test_number = 1;
    reset_all();
    #1000;
    @(negedge i_clock) begin
        i_in_valid = 1'b0;
        #(10000);
    end
    i_in_valid = 1'b0;
    #1000;
    if (run_count > 0) begin
        $display("Error: Test 1 failed! No data input, but data output received.");
        glbl_err_count++;
    end
    #100;
    $display("Test 1 Done!");

    // Test 2: Produce codeword 0.
    $display("Test 2 Started!");
    test_number = 2;
    reset_all();
    #10000;
    i_out_ready = 1'b1;
    #1000;
    for (count = 0; count < SLENGTH/8; count++) begin
        @(negedge i_clock) begin
            i_in_valid = 1'b1;
            i_in_data = {
                ldpc_codeword_0[count*8 + 7],
                ldpc_codeword_0[count*8 + 6],
                ldpc_codeword_0[count*8 + 5],
                ldpc_codeword_0[count*8 + 4],
                ldpc_codeword_0[count*8 + 3],
                ldpc_codeword_0[count*8 + 2],
                ldpc_codeword_0[count*8 + 1],
                ldpc_codeword_0[count*8    ]
            };
            if (o_in_ready == 1'b1) begin
                #10;
            end else begin
                @(posedge o_in_ready) begin
                    #10;
                end
            end
        end
    end
    i_in_data = 0;
    i_in_valid = 1'b0;
    #(10*(4*CLENGTH));
    i_out_ready = 1'b0;
    #100;
    if (run_count != CLENGTH/8) begin
        $display("Error: Test 2 failed! Expected %d but received %d outputs.", CLENGTH/8, run_count);
        glbl_err_count++;
    end
    $display("Test 1 Done!");

    // Finished
    #10000;
    glbl_err_count = glbl_err_count + local_err_count;
    #10;
    $display("Simulation done!");
    if (glbl_err_count > 0) begin
        $display("Found %d errors!", glbl_err_count);
    end else begin
        $display("<< Success! >>");
    end

    $display("rx_cwd = [",);
    for (count = 0; count < CLENGTH; count++) begin
        $display("%b", ldpc_encoded_codeword_0[count]);
    end
    $display("];",);
    $finish();

end

// Tests the output sequence to make sure it matches the input
logic [7:0] expected_value;
always @(posedge i_clock) begin: seq_check
    if (i_reset == 1'b1) begin
        run_count <= 0;
    end else begin
        // Track number of outputs received
        if ((o_out_valid == 1'b1) && (i_out_ready == 1'b1)) begin
            if (test_number == 2) begin
                expected_value = {
                    ldpc_codeword_0[8 * run_count + 7],
                    ldpc_codeword_0[8 * run_count + 6],
                    ldpc_codeword_0[8 * run_count + 5],
                    ldpc_codeword_0[8 * run_count + 4],
                    ldpc_codeword_0[8 * run_count + 3],
                    ldpc_codeword_0[8 * run_count + 2],
                    ldpc_codeword_0[8 * run_count + 1],
                    ldpc_codeword_0[8 * run_count    ]
                };
                if (o_out_data != expected_value) begin
                    $display("Expected %b but received %b (run_count = %d)",
                        expected_value, o_out_data, run_count);
                    local_err_count++;
                end
                ldpc_encoded_codeword_0[8 * run_count + 7] <= o_out_data[7];
                ldpc_encoded_codeword_0[8 * run_count + 6] <= o_out_data[6];
                ldpc_encoded_codeword_0[8 * run_count + 5] <= o_out_data[5];
                ldpc_encoded_codeword_0[8 * run_count + 4] <= o_out_data[4];
                ldpc_encoded_codeword_0[8 * run_count + 3] <= o_out_data[3];
                ldpc_encoded_codeword_0[8 * run_count + 2] <= o_out_data[2];
                ldpc_encoded_codeword_0[8 * run_count + 1] <= o_out_data[1];
                ldpc_encoded_codeword_0[8 * run_count    ] <= o_out_data[0];
            end
            run_count <= run_count + 1;
        end
    end
end

endmodule: tb_ldpc_encoder

`default_nettype wire
