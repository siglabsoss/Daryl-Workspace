`timescale 10ps / 10ps

`default_nettype none

module ldpc_decode_stage (

);



endmodule: ldpc_decode_stage

`default_nettype wire